library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;


package cc_regn is

    procedure regn_check (constant program : in instructions);

end package;


package body cc_regn is

    procedure regn_check (constant program : in instructions) is
    begin

        assert program(0).src = 1 report "0 src Failed" severity FAILURE;
        assert program(0).dst = 2 report "0 dst Failed" severity FAILURE;
        assert program(1).src = 2 report "1 src Failed" severity FAILURE;
        assert program(1).dst = 1 report "1 dst Failed" severity FAILURE;
        assert program(2).src = 6 report "2 src Failed" severity FAILURE;
        assert program(2).dst = 6 report "2 dst Failed" severity FAILURE;
        assert program(3).src = 0 report "3 src Failed" severity FAILURE;
        assert program(3).dst = 1 report "3 dst Failed" severity FAILURE;
        assert program(4).src = 3 report "4 src Failed" severity FAILURE;
        assert program(4).dst = 6 report "4 dst Failed" severity FAILURE;
        assert program(5).dst = 7 report "5 dst Failed" severity FAILURE;
        assert program(6).src = 2 report "6 src Failed" severity FAILURE;
        assert program(6).dst = 3 report "6 dst Failed" severity FAILURE;
        assert program(7).src = 0 report "7 src Failed" severity FAILURE;
        assert program(7).dst = 0 report "7 dst Failed" severity FAILURE;
        assert program(8).src = 5 report "8 src Failed" severity FAILURE;
        assert program(8).dst = 1 report "8 dst Failed" severity FAILURE;
        assert program(9).dst = 7 report "9 dst Failed" severity FAILURE;
        assert program(10).src = 1 report "10 src Failed" severity FAILURE;
        assert program(10).dst = 0 report "10 dst Failed" severity FAILURE;
        assert program(11).src = 3 report "11 src Failed" severity FAILURE;
        assert program(11).dst = 3 report "11 dst Failed" severity FAILURE;
        assert program(12).src = 3 report "12 src Failed" severity FAILURE;
        assert program(12).dst = 1 report "12 dst Failed" severity FAILURE;
        assert program(13).src = 4 report "13 src Failed" severity FAILURE;
        assert program(13).dst = 4 report "13 dst Failed" severity FAILURE;
        assert program(14).dst = 6 report "14 dst Failed" severity FAILURE;
        assert program(15).src = 0 report "15 src Failed" severity FAILURE;
        assert program(15).dst = 1 report "15 dst Failed" severity FAILURE;
        assert program(16).src = 1 report "16 src Failed" severity FAILURE;
        assert program(16).dst = 2 report "16 dst Failed" severity FAILURE;
        assert program(17).src = 0 report "17 src Failed" severity FAILURE;
        assert program(17).dst = 4 report "17 dst Failed" severity FAILURE;
        assert program(18).src = 3 report "18 src Failed" severity FAILURE;
        assert program(18).dst = 6 report "18 dst Failed" severity FAILURE;
        assert program(19).dst = 5 report "19 dst Failed" severity FAILURE;
        assert program(20).src = 0 report "20 src Failed" severity FAILURE;
        assert program(20).dst = 2 report "20 dst Failed" severity FAILURE;
        assert program(21).src = 3 report "21 src Failed" severity FAILURE;
        assert program(21).dst = 0 report "21 dst Failed" severity FAILURE;
        assert program(22).src = 0 report "22 src Failed" severity FAILURE;
        assert program(22).dst = 5 report "22 dst Failed" severity FAILURE;
        assert program(23).src = 3 report "23 src Failed" severity FAILURE;
        assert program(23).dst = 0 report "23 dst Failed" severity FAILURE;
        assert program(24).src = 7 report "24 src Failed" severity FAILURE;
        assert program(24).dst = 0 report "24 dst Failed" severity FAILURE;
        assert program(25).src = 4 report "25 src Failed" severity FAILURE;
        assert program(25).dst = 2 report "25 dst Failed" severity FAILURE;
        assert program(26).src = 5 report "26 src Failed" severity FAILURE;
        assert program(26).dst = 2 report "26 dst Failed" severity FAILURE;
        assert program(27).src = 0 report "27 src Failed" severity FAILURE;
        assert program(27).dst = 3 report "27 dst Failed" severity FAILURE;
        assert program(28).dst = 2 report "28 dst Failed" severity FAILURE;
        assert program(29).src = 4 report "29 src Failed" severity FAILURE;
        assert program(29).dst = 5 report "29 dst Failed" severity FAILURE;
        assert program(30).src = 3 report "30 src Failed" severity FAILURE;
        assert program(30).dst = 2 report "30 dst Failed" severity FAILURE;
        assert program(31).src = 6 report "31 src Failed" severity FAILURE;
        assert program(31).dst = 1 report "31 dst Failed" severity FAILURE;
        assert program(32).src = 1 report "32 src Failed" severity FAILURE;
        assert program(32).dst = 1 report "32 dst Failed" severity FAILURE;
        assert program(33).src = 0 report "33 src Failed" severity FAILURE;
        assert program(33).dst = 3 report "33 dst Failed" severity FAILURE;
        assert program(34).src = -1 report "34 src Failed" severity FAILURE;
        assert program(34).dst = 0 report "34 dst Failed" severity FAILURE;
        assert program(35).dst = 9 report "35 dst Failed" severity FAILURE;
        assert program(36).src = 3 report "36 src Failed" severity FAILURE;
        assert program(36).dst = 5 report "36 dst Failed" severity FAILURE;
        assert program(37).dst = 7 report "37 dst Failed" severity FAILURE;
        assert program(38).dst = 1 report "38 dst Failed" severity FAILURE;
        assert program(39).src = -1 report "39 src Failed" severity FAILURE;
        assert program(39).dst = 5 report "39 dst Failed" severity FAILURE;
        assert program(40).src = 0 report "40 src Failed" severity FAILURE;
        assert program(40).dst = 5 report "40 dst Failed" severity FAILURE;
        assert program(41).src = 3 report "41 src Failed" severity FAILURE;
        assert program(41).dst = 0 report "41 dst Failed" severity FAILURE;
        assert program(42).src = 0 report "42 src Failed" severity FAILURE;
        assert program(42).dst = 6 report "42 dst Failed" severity FAILURE;
        assert program(43).dst = 2 report "43 dst Failed" severity FAILURE;
        assert program(44).src = 5 report "44 src Failed" severity FAILURE;
        assert program(44).dst = 3 report "44 dst Failed" severity FAILURE;
        assert program(45).src = 0 report "45 src Failed" severity FAILURE;
        assert program(45).dst = 4 report "45 dst Failed" severity FAILURE;
        assert program(46).src = 6 report "46 src Failed" severity FAILURE;
        assert program(46).dst = 7 report "46 dst Failed" severity FAILURE;
        assert program(47).src = 6 report "47 src Failed" severity FAILURE;
        assert program(47).dst = 0 report "47 dst Failed" severity FAILURE;
        assert program(48).src = 1 report "48 src Failed" severity FAILURE;
        assert program(48).dst = 1 report "48 dst Failed" severity FAILURE;
        assert program(49).src = 0 report "49 src Failed" severity FAILURE;
        assert program(49).dst = 2 report "49 dst Failed" severity FAILURE;
        assert program(50).src = 2 report "50 src Failed" severity FAILURE;
        assert program(50).dst = 0 report "50 dst Failed" severity FAILURE;
        assert program(51).src = 3 report "51 src Failed" severity FAILURE;
        assert program(51).dst = 2 report "51 dst Failed" severity FAILURE;
        assert program(52).src = -1 report "52 src Failed" severity FAILURE;
        assert program(52).dst = 7 report "52 dst Failed" severity FAILURE;
        assert program(53).src = 2 report "53 src Failed" severity FAILURE;
        assert program(53).dst = 0 report "53 dst Failed" severity FAILURE;
        assert program(54).src = 6 report "54 src Failed" severity FAILURE;
        assert program(54).dst = 3 report "54 dst Failed" severity FAILURE;
        assert program(55).dst = 1 report "55 dst Failed" severity FAILURE;
        assert program(57).src = 1 report "57 src Failed" severity FAILURE;
        assert program(57).dst = 0 report "57 dst Failed" severity FAILURE;
        assert program(58).src = -1 report "58 src Failed" severity FAILURE;
        assert program(58).dst = 1 report "58 dst Failed" severity FAILURE;
        assert program(59).dst = 7 report "59 dst Failed" severity FAILURE;
        assert program(60).src = 3 report "60 src Failed" severity FAILURE;
        assert program(60).dst = 6 report "60 dst Failed" severity FAILURE;
        assert program(61).src = 4 report "61 src Failed" severity FAILURE;
        assert program(61).dst = 3 report "61 dst Failed" severity FAILURE;
        assert program(62).src = 0 report "62 src Failed" severity FAILURE;
        assert program(62).dst = 3 report "62 dst Failed" severity FAILURE;
        assert program(63).src = 2 report "63 src Failed" severity FAILURE;
        assert program(63).dst = 3 report "63 dst Failed" severity FAILURE;
        assert program(64).src = 2 report "64 src Failed" severity FAILURE;
        assert program(64).dst = 6 report "64 dst Failed" severity FAILURE;
        assert program(65).src = 5 report "65 src Failed" severity FAILURE;
        assert program(65).dst = 0 report "65 dst Failed" severity FAILURE;
        assert program(66).src = 3 report "66 src Failed" severity FAILURE;
        assert program(66).dst = 1 report "66 dst Failed" severity FAILURE;
        assert program(67).src = 1 report "67 src Failed" severity FAILURE;
        assert program(67).dst = 7 report "67 dst Failed" severity FAILURE;
        assert program(68).src = 4 report "68 src Failed" severity FAILURE;
        assert program(68).dst = 7 report "68 dst Failed" severity FAILURE;
        assert program(69).src = 3 report "69 src Failed" severity FAILURE;
        assert program(69).dst = 2 report "69 dst Failed" severity FAILURE;
        assert program(70).src = 0 report "70 src Failed" severity FAILURE;
        assert program(70).dst = 2 report "70 dst Failed" severity FAILURE;
        assert program(71).dst = 6 report "71 dst Failed" severity FAILURE;
        assert program(72).dst = 3 report "72 dst Failed" severity FAILURE;
        assert program(73).src = 5 report "73 src Failed" severity FAILURE;
        assert program(73).dst = 0 report "73 dst Failed" severity FAILURE;
        assert program(74).src = 0 report "74 src Failed" severity FAILURE;
        assert program(74).dst = 1 report "74 dst Failed" severity FAILURE;
        assert program(75).src = 0 report "75 src Failed" severity FAILURE;
        assert program(75).dst = 1 report "75 dst Failed" severity FAILURE;
        assert program(76).src = 1 report "76 src Failed" severity FAILURE;
        assert program(76).dst = 2 report "76 dst Failed" severity FAILURE;
        assert program(77).src = 1 report "77 src Failed" severity FAILURE;
        assert program(77).dst = 0 report "77 dst Failed" severity FAILURE;
        assert program(78).dst = 1 report "78 dst Failed" severity FAILURE;
        assert program(79).src = 7 report "79 src Failed" severity FAILURE;
        assert program(79).dst = 0 report "79 dst Failed" severity FAILURE;
        assert program(80).src = 4 report "80 src Failed" severity FAILURE;
        assert program(80).dst = 3 report "80 dst Failed" severity FAILURE;
        assert program(81).src = 1 report "81 src Failed" severity FAILURE;
        assert program(81).dst = 4 report "81 dst Failed" severity FAILURE;
        assert program(82).src = 4 report "82 src Failed" severity FAILURE;
        assert program(82).dst = 0 report "82 dst Failed" severity FAILURE;
        assert program(83).src = 4 report "83 src Failed" severity FAILURE;
        assert program(83).dst = 1 report "83 dst Failed" severity FAILURE;
        assert program(84).src = 5 report "84 src Failed" severity FAILURE;
        assert program(84).dst = 3 report "84 dst Failed" severity FAILURE;
        assert program(85).src = 5 report "85 src Failed" severity FAILURE;
        assert program(85).dst = 3 report "85 dst Failed" severity FAILURE;
        assert program(86).src = 2 report "86 src Failed" severity FAILURE;
        assert program(86).dst = 3 report "86 dst Failed" severity FAILURE;
        assert program(87).dst = 1 report "87 dst Failed" severity FAILURE;
        assert program(88).src = 4 report "88 src Failed" severity FAILURE;
        assert program(88).dst = 3 report "88 dst Failed" severity FAILURE;
        assert program(89).src = 1 report "89 src Failed" severity FAILURE;
        assert program(89).dst = 2 report "89 dst Failed" severity FAILURE;
        assert program(90).src = 2 report "90 src Failed" severity FAILURE;
        assert program(90).dst = 7 report "90 dst Failed" severity FAILURE;
        assert program(91).src = 5 report "91 src Failed" severity FAILURE;
        assert program(91).dst = 3 report "91 dst Failed" severity FAILURE;
        assert program(92).src = 1 report "92 src Failed" severity FAILURE;
        assert program(92).dst = 2 report "92 dst Failed" severity FAILURE;
        assert program(93).dst = 2 report "93 dst Failed" severity FAILURE;
        assert program(94).src = 2 report "94 src Failed" severity FAILURE;
        assert program(94).dst = 0 report "94 dst Failed" severity FAILURE;
        assert program(95).src = 2 report "95 src Failed" severity FAILURE;
        assert program(95).dst = 0 report "95 dst Failed" severity FAILURE;
        assert program(96).src = 1 report "96 src Failed" severity FAILURE;
        assert program(96).dst = 0 report "96 dst Failed" severity FAILURE;
        assert program(97).src = 6 report "97 src Failed" severity FAILURE;
        assert program(97).dst = 4 report "97 dst Failed" severity FAILURE;
        assert program(98).src = 5 report "98 src Failed" severity FAILURE;
        assert program(98).dst = 3 report "98 dst Failed" severity FAILURE;
        assert program(99).src = 2 report "99 src Failed" severity FAILURE;
        assert program(99).dst = 0 report "99 dst Failed" severity FAILURE;
        assert program(100).src = 0 report "100 src Failed" severity FAILURE;
        assert program(100).dst = 5 report "100 dst Failed" severity FAILURE;
        assert program(101).src = 0 report "101 src Failed" severity FAILURE;
        assert program(101).dst = 2 report "101 dst Failed" severity FAILURE;
        assert program(102).src = 2 report "102 src Failed" severity FAILURE;
        assert program(102).dst = 6 report "102 dst Failed" severity FAILURE;
        assert program(103).src = 6 report "103 src Failed" severity FAILURE;
        assert program(103).dst = 4 report "103 dst Failed" severity FAILURE;
        assert program(104).src = 6 report "104 src Failed" severity FAILURE;
        assert program(104).dst = 0 report "104 dst Failed" severity FAILURE;
        assert program(105).src = 2 report "105 src Failed" severity FAILURE;
        assert program(105).dst = 4 report "105 dst Failed" severity FAILURE;
        assert program(106).src = -1 report "106 src Failed" severity FAILURE;
        assert program(106).dst = 0 report "106 dst Failed" severity FAILURE;
        assert program(107).src = 1 report "107 src Failed" severity FAILURE;
        assert program(107).dst = 2 report "107 dst Failed" severity FAILURE;
        assert program(108).src = 4 report "108 src Failed" severity FAILURE;
        assert program(108).dst = 0 report "108 dst Failed" severity FAILURE;
        assert program(109).src = 5 report "109 src Failed" severity FAILURE;
        assert program(109).dst = 3 report "109 dst Failed" severity FAILURE;
        assert program(110).src = 4 report "110 src Failed" severity FAILURE;
        assert program(110).dst = 3 report "110 dst Failed" severity FAILURE;
        assert program(111).src = 1 report "111 src Failed" severity FAILURE;
        assert program(111).dst = 0 report "111 dst Failed" severity FAILURE;
        assert program(112).src = 4 report "112 dst Failed" severity FAILURE;
        assert program(113).dst = 6 report "113 dst Failed" severity FAILURE;
        assert program(114).src = 6 report "114 src Failed" severity FAILURE;
        assert program(114).dst = 7 report "114 dst Failed" severity FAILURE;
        assert program(115).dst = 2 report "115 dst Failed" severity FAILURE;
        assert program(116).src = 2 report "116 src Failed" severity FAILURE;
        assert program(116).dst = 6 report "116 dst Failed" severity FAILURE;
        assert program(117).src = 1 report "117 src Failed" severity FAILURE;
        assert program(117).dst = 0 report "117 dst Failed" severity FAILURE;
        assert program(118).src = 0 report "118 src Failed" severity FAILURE;
        assert program(118).dst = 0 report "118 dst Failed" severity FAILURE;
        assert program(119).src = 0 report "119 src Failed" severity FAILURE;
        assert program(119).dst = 2 report "119 dst Failed" severity FAILURE;
        assert program(120).src = 3 report "120 src Failed" severity FAILURE;
        assert program(120).dst = 7 report "120 dst Failed" severity FAILURE;
        assert program(121).src = 7 report "121 src Failed" severity FAILURE;
        assert program(121).dst = 7 report "121 dst Failed" severity FAILURE;
        assert program(122).src = -1 report "122 src Failed" severity FAILURE;
        assert program(122).dst = 3 report "122 dst Failed" severity FAILURE;
        assert program(123).src = 7 report "123 src Failed" severity FAILURE;
        assert program(123).dst = 2 report "123 dst Failed" severity FAILURE;
        assert program(124).dst = 7 report "124 dst Failed" severity FAILURE;
        assert program(125).src = 2 report "125 src Failed" severity FAILURE;
        assert program(125).dst = 0 report "125 dst Failed" severity FAILURE;
        assert program(126).src = 2 report "126 src Failed" severity FAILURE;
        assert program(126).dst = 3 report "126 dst Failed" severity FAILURE;
        assert program(127).src = 4 report "127 src Failed" severity FAILURE;
        assert program(127).dst = 6 report "127 dst Failed" severity FAILURE;
        assert program(128).src = 4 report "128 src Failed" severity FAILURE;
        assert program(128).dst = 2 report "128 dst Failed" severity FAILURE;
        assert program(129).src = 0 report "129 src Failed" severity FAILURE;
        assert program(129).dst = 2 report "129 dst Failed" severity FAILURE;
        assert program(130).src = 6 report "130 src Failed" severity FAILURE;
        assert program(130).dst = 4 report "130 dst Failed" severity FAILURE;
        assert program(131).dst = 5 report "131 dst Failed" severity FAILURE;
        assert program(132).src = 1 report "132 src Failed" severity FAILURE;
        assert program(132).dst = 1 report "132 dst Failed" severity FAILURE;
        assert program(133).src = 6 report "133 src Failed" severity FAILURE;
        assert program(133).dst = 4 report "133 dst Failed" severity FAILURE;
        assert program(134).dst = 5 report "134 dst Failed" severity FAILURE;
        assert program(135).src = 4 report "135 src Failed" severity FAILURE;
        assert program(135).dst = 4 report "135 dst Failed" severity FAILURE;
        assert program(136).src = 2 report "136 src Failed" severity FAILURE;
        assert program(136).dst = 1 report "136 dst Failed" severity FAILURE;
        assert program(137).src = 2 report "137 src Failed" severity FAILURE;
        assert program(137).dst = 0 report "137 dst Failed" severity FAILURE;
        assert program(138).dst = 1 report "138 dst Failed" severity FAILURE;
        assert program(139).src = 7 report "139 src Failed" severity FAILURE;
        assert program(139).dst = 5 report "139 dst Failed" severity FAILURE;
        assert program(140).src = 2 report "140 src Failed" severity FAILURE;
        assert program(140).dst = 7 report "140 dst Failed" severity FAILURE;
        assert program(141).dst = 3 report "141 dst Failed" severity FAILURE;
        assert program(142).src = 3 report "142 src Failed" severity FAILURE;
        assert program(142).dst = 7 report "142 dst Failed" severity FAILURE;
        assert program(143).src = 2 report "143 src Failed" severity FAILURE;
        assert program(143).dst = 2 report "143 dst Failed" severity FAILURE;
        assert program(144).src = 1 report "144 src Failed" severity FAILURE;
        assert program(144).dst = 7 report "144 dst Failed" severity FAILURE;
        assert program(145).src = 0 report "145 src Failed" severity FAILURE;
        assert program(145).dst = 3 report "145 dst Failed" severity FAILURE;
        assert program(146).src = 5 report "146 src Failed" severity FAILURE;
        assert program(146).dst = 3 report "146 dst Failed" severity FAILURE;
        assert program(147).src = 0 report "147 src Failed" severity FAILURE;
        assert program(147).dst = 3 report "147 dst Failed" severity FAILURE;
        assert program(148).src = 5 report "148 src Failed" severity FAILURE;
        assert program(148).dst = 3 report "148 dst Failed" severity FAILURE;
        assert program(149).src = 2 report "149 src Failed" severity FAILURE;
        assert program(149).dst = 3 report "149 dst Failed" severity FAILURE;
        assert program(150).src = 3 report "150 src Failed" severity FAILURE;
        assert program(150).dst = 1 report "150 dst Failed" severity FAILURE;
        assert program(151).src = 5 report "151 src Failed" severity FAILURE;
        assert program(151).dst = 6 report "151 dst Failed" severity FAILURE;
        assert program(152).dst = 5 report "152 dst Failed" severity FAILURE;
        assert program(153).src = 0 report "153 src Failed" severity FAILURE;
        assert program(153).dst = 1 report "153 dst Failed" severity FAILURE;
        assert program(154).src = 2 report "154 src Failed" severity FAILURE;
        assert program(154).dst = 5 report "154 dst Failed" severity FAILURE;
        assert program(155).src = 2 report "155 src Failed" severity FAILURE;
        assert program(155).dst = 1 report "155 dst Failed" severity FAILURE;
        assert program(156).src = 2 report "156 src Failed" severity FAILURE;
        assert program(156).dst = 5 report "156 dst Failed" severity FAILURE;
        assert program(157).src = 0 report "157 src Failed" severity FAILURE;
        assert program(157).dst = 5 report "157 dst Failed" severity FAILURE;
        assert program(158).src = 2 report "158 src Failed" severity FAILURE;
        assert program(158).dst = 2 report "158 dst Failed" severity FAILURE;
        assert program(159).dst = 7 report "159 dst Failed" severity FAILURE;
        assert program(160).src = 2 report "160 src Failed" severity FAILURE;
        assert program(160).dst = 1 report "160 dst Failed" severity FAILURE;
        assert program(161).src = 2 report "161 src Failed" severity FAILURE;
        assert program(161).dst = 1 report "161 dst Failed" severity FAILURE;
        assert program(162).src = 1 report "162 src Failed" severity FAILURE;
        assert program(162).dst = 2 report "162 dst Failed" severity FAILURE;
        assert program(163).src = 3 report "163 src Failed" severity FAILURE;
        assert program(163).dst = 7 report "163 dst Failed" severity FAILURE;
        assert program(164).dst = 7 report "164 dst Failed" severity FAILURE;
        assert program(165).src = -1 report "165 src Failed" severity FAILURE;
        assert program(165).dst = 7 report "165 dst Failed" severity FAILURE;
        assert program(166).src = 1 report "166 src Failed" severity FAILURE;
        assert program(166).dst = 0 report "166 dst Failed" severity FAILURE;
        assert program(167).src = 2 report "167 src Failed" severity FAILURE;
        assert program(167).dst = 0 report "167 dst Failed" severity FAILURE;
        assert program(168).dst = 6 report "168 dst Failed" severity FAILURE;
        assert program(169).src = 3 report "169 src Failed" severity FAILURE;
        assert program(169).dst = 0 report "169 dst Failed" severity FAILURE;
        assert program(170).src = -1 report "170 src Failed" severity FAILURE;
        assert program(170).dst = 2 report "170 dst Failed" severity FAILURE;
        assert program(171).dst = 3 report "171 dst Failed" severity FAILURE;
        assert program(172).src = 3 report "172 src Failed" severity FAILURE;
        assert program(172).dst = 2 report "172 dst Failed" severity FAILURE;
        assert program(173).src = 2 report "173 src Failed" severity FAILURE;
        assert program(173).dst = 3 report "173 dst Failed" severity FAILURE;
        assert program(174).dst = 0 report "174 dst Failed" severity FAILURE;
        assert program(175).src = 1 report "175 src Failed" severity FAILURE;
        assert program(175).dst = 2 report "175 dst Failed" severity FAILURE;
        assert program(176).src = 2 report "176 src Failed" severity FAILURE;
        assert program(176).dst = 1 report "176 dst Failed" severity FAILURE;
        assert program(177).src = 0 report "177 src Failed" severity FAILURE;
        assert program(177).dst = 1 report "177 dst Failed" severity FAILURE;
        assert program(178).src = 1 report "178 src Failed" severity FAILURE;
        assert program(178).dst = 1 report "178 dst Failed" severity FAILURE;
        assert program(179).src = 6 report "179 src Failed" severity FAILURE;
        assert program(179).dst = 1 report "179 dst Failed" severity FAILURE;
        assert program(180).src = 6 report "180 src Failed" severity FAILURE;
        assert program(180).dst = 1 report "180 dst Failed" severity FAILURE;
        assert program(181).src = 6 report "181 src Failed" severity FAILURE;
        assert program(181).dst = 4 report "181 dst Failed" severity FAILURE;
        assert program(182).src = 6 report "182 src Failed" severity FAILURE;
        assert program(182).dst = 0 report "182 dst Failed" severity FAILURE;
        assert program(183).dst = 0 report "183 dst Failed" severity FAILURE;
        assert program(184).dst = 6 report "184 dst Failed" severity FAILURE;
        assert program(185).src = 6 report "185 src Failed" severity FAILURE;
        assert program(185).dst = 2 report "185 dst Failed" severity FAILURE;
        assert program(186).src = 1 report "186 src Failed" severity FAILURE;
        assert program(186).dst = 2 report "186 dst Failed" severity FAILURE;
        assert program(187).dst = 6 report "187 dst Failed" severity FAILURE;
        assert program(188).dst = 2 report "188 dst Failed" severity FAILURE;
        assert program(189).src = 2 report "189 src Failed" severity FAILURE;
        assert program(189).dst = 0 report "189 dst Failed" severity FAILURE;
        assert program(190).src = 6 report "190 src Failed" severity FAILURE;
        assert program(190).dst = 3 report "190 dst Failed" severity FAILURE;
        assert program(191).dst = 5 report "191 dst Failed" severity FAILURE;
        assert program(192).src = -1 report "192 src Failed" severity FAILURE;
        assert program(192).dst = 2 report "192 dst Failed" severity FAILURE;
        assert program(193).src = 6 report "193 src Failed" severity FAILURE;
        assert program(193).dst = 5 report "193 dst Failed" severity FAILURE;
        assert program(194).src = 4 report "194 src Failed" severity FAILURE;
        assert program(194).dst = 3 report "194 dst Failed" severity FAILURE;
        assert program(195).dst = 7 report "195 dst Failed" severity FAILURE;
        assert program(196).dst = 1 report "196 dst Failed" severity FAILURE;
        assert program(197).dst = 4 report "197 dst Failed" severity FAILURE;
        assert program(198).dst = 3 report "198 dst Failed" severity FAILURE;
        assert program(199).src = 0 report "199 src Failed" severity FAILURE;
        assert program(199).dst = 2 report "199 dst Failed" severity FAILURE;
        assert program(200).src = 3 report "200 src Failed" severity FAILURE;
        assert program(200).dst = 0 report "200 dst Failed" severity FAILURE;
        assert program(201).src = 1 report "201 src Failed" severity FAILURE;
        assert program(201).dst = 3 report "201 dst Failed" severity FAILURE;
        assert program(202).src = 2 report "202 src Failed" severity FAILURE;
        assert program(202).dst = 3 report "202 dst Failed" severity FAILURE;
        assert program(203).src = 2 report "203 src Failed" severity FAILURE;
        assert program(203).dst = 3 report "203 dst Failed" severity FAILURE;
        assert program(204).src = 2 report "204 src Failed" severity FAILURE;
        assert program(204).dst = 0 report "204 dst Failed" severity FAILURE;
        assert program(205).src = 3 report "205 src Failed" severity FAILURE;
        assert program(205).dst = 6 report "205 dst Failed" severity FAILURE;
        assert program(206).src = 3 report "206 src Failed" severity FAILURE;
        assert program(206).dst = 6 report "206 dst Failed" severity FAILURE;
        assert program(207).src = 5 report "207 src Failed" severity FAILURE;
        assert program(207).dst = 7 report "207 dst Failed" severity FAILURE;
        assert program(208).src = 3 report "208 src Failed" severity FAILURE;
        assert program(208).dst = 3 report "208 dst Failed" severity FAILURE;
        assert program(209).src = 0 report "209 src Failed" severity FAILURE;
        assert program(209).dst = 2 report "209 dst Failed" severity FAILURE;
        assert program(210).dst = 2 report "210 dst Failed" severity FAILURE;
        assert program(211).src = 0 report "211 src Failed" severity FAILURE;
        assert program(211).dst = 5 report "211 dst Failed" severity FAILURE;
        assert program(212).src = 5 report "212 src Failed" severity FAILURE;
        assert program(212).dst = 7 report "212 dst Failed" severity FAILURE;
        assert program(213).src = 5 report "213 src Failed" severity FAILURE;
        assert program(213).dst = 3 report "213 dst Failed" severity FAILURE;
        assert program(214).src = 2 report "214 src Failed" severity FAILURE;
        assert program(214).dst = 4 report "214 dst Failed" severity FAILURE;
        assert program(215).dst = 6 report "215 dst Failed" severity FAILURE;
        assert program(216).dst = 2 report "216 dst Failed" severity FAILURE;
        assert program(217).src = -1 report "217 src Failed" severity FAILURE;
        assert program(217).dst = 1 report "217 dst Failed" severity FAILURE;
        assert program(218).src = 1 report "218 src Failed" severity FAILURE;
        assert program(218).dst = 4 report "218 dst Failed" severity FAILURE;
        assert program(219).src = 6 report "219 src Failed" severity FAILURE;
        assert program(219).dst = 3 report "219 dst Failed" severity FAILURE;
        assert program(220).src = 5 report "220 src Failed" severity FAILURE;
        assert program(220).dst = 3 report "220 dst Failed" severity FAILURE;
        assert program(221).src = 2 report "221 src Failed" severity FAILURE;
        assert program(221).dst = 0 report "221 dst Failed" severity FAILURE;
        assert program(222).src = 0 report "222 src Failed" severity FAILURE;
        assert program(222).dst = 1 report "222 dst Failed" severity FAILURE;
        assert program(223).src = 0 report "223 src Failed" severity FAILURE;
        assert program(223).dst = 7 report "223 dst Failed" severity FAILURE;
        assert program(224).src = 3 report "224 src Failed" severity FAILURE;
        assert program(224).dst = 1 report "224 dst Failed" severity FAILURE;
        assert program(225).src = 1 report "225 src Failed" severity FAILURE;
        assert program(225).dst = 3 report "225 dst Failed" severity FAILURE;
        assert program(226).src = 3 report "226 src Failed" severity FAILURE;
        assert program(226).dst = 3 report "226 dst Failed" severity FAILURE;
        assert program(227).src = 3 report "227 src Failed" severity FAILURE;
        assert program(227).dst = 1 report "227 dst Failed" severity FAILURE;
        assert program(228).src = 0 report "228 src Failed" severity FAILURE;
        assert program(228).dst = 1 report "228 dst Failed" severity FAILURE;
        assert program(229).src = 3 report "229 src Failed" severity FAILURE;
        assert program(229).dst = 0 report "229 dst Failed" severity FAILURE;
        assert program(230).src = 1 report "230 src Failed" severity FAILURE;
        assert program(230).dst = 1 report "230 dst Failed" severity FAILURE;
        assert program(231).src = 2 report "231 src Failed" severity FAILURE;
        assert program(231).dst = 4 report "231 dst Failed" severity FAILURE;
        assert program(232).src = 1 report "232 src Failed" severity FAILURE;
        assert program(232).dst = 2 report "232 dst Failed" severity FAILURE;
        assert program(233).src = 2 report "233 src Failed" severity FAILURE;
        assert program(233).dst = 0 report "233 dst Failed" severity FAILURE;
        assert program(234).dst = 0 report "234 dst Failed" severity FAILURE;
        assert program(235).src = 1 report "235 src Failed" severity FAILURE;
        assert program(235).dst = 4 report "235 dst Failed" severity FAILURE;
        assert program(236).src = -1 report "236 src Failed" severity FAILURE;
        assert program(236).dst = 4 report "236 dst Failed" severity FAILURE;
        assert program(237).src = 3 report "237 src Failed" severity FAILURE;
        assert program(237).dst = 3 report "237 dst Failed" severity FAILURE;
        assert program(238).src = 5 report "238 src Failed" severity FAILURE;
        assert program(238).dst = 0 report "238 dst Failed" severity FAILURE;
        assert program(239).src = 7 report "239 src Failed" severity FAILURE;
        assert program(239).dst = 3 report "239 dst Failed" severity FAILURE;
        assert program(240).src = 3 report "240 src Failed" severity FAILURE;
        assert program(240).dst = 1 report "240 dst Failed" severity FAILURE;
        assert program(241).src = 1 report "241 src Failed" severity FAILURE;
        assert program(241).dst = 0 report "241 dst Failed" severity FAILURE;
        assert program(242).src = 0 report "242 src Failed" severity FAILURE;
        assert program(242).dst = 1 report "242 dst Failed" severity FAILURE;
        assert program(243).src = 0 report "243 src Failed" severity FAILURE;
        assert program(243).dst = 5 report "243 dst Failed" severity FAILURE;
        assert program(244).src = 3 report "244 src Failed" severity FAILURE;
        assert program(244).dst = 1 report "244 dst Failed" severity FAILURE;
        assert program(245).src = 7 report "245 src Failed" severity FAILURE;
        assert program(245).dst = 3 report "245 dst Failed" severity FAILURE;
        assert program(246).src = 7 report "246 src Failed" severity FAILURE;
        assert program(246).dst = 0 report "246 dst Failed" severity FAILURE;
        assert program(247).src = 2 report "247 src Failed" severity FAILURE;
        assert program(247).dst = 2 report "247 dst Failed" severity FAILURE;
        assert program(248).src = 1 report "248 src Failed" severity FAILURE;
        assert program(248).dst = 7 report "248 dst Failed" severity FAILURE;
        assert program(249).src = 3 report "249 src Failed" severity FAILURE;
        assert program(249).dst = 3 report "249 dst Failed" severity FAILURE;
        assert program(250).src = 7 report "250 src Failed" severity FAILURE;
        assert program(250).dst = 3 report "250 dst Failed" severity FAILURE;
        assert program(251).src = 1 report "251 src Failed" severity FAILURE;
        assert program(251).dst = 1 report "251 dst Failed" severity FAILURE;
        assert program(252).src = 0 report "252 src Failed" severity FAILURE;
        assert program(252).dst = 4 report "252 dst Failed" severity FAILURE;
        assert program(253).dst = 2 report "253 dst Failed" severity FAILURE;
        assert program(254).src = 1 report "254 src Failed" severity FAILURE;
        assert program(254).dst = 0 report "254 dst Failed" severity FAILURE;
        assert program(255).src = 0 report "255 src Failed" severity FAILURE;
        assert program(255).dst = 3 report "255 dst Failed" severity FAILURE;

    end;

end cc_regn;