library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;


package cc_opcode is

    procedure opcode_check (constant program : in instructions);

end package;


package body cc_opcode is

    procedure opcode_check (constant program : in instructions) is
    begin

        assert program(0).op = FSUB_M report "0 FSUB_M Failed" severity FAILURE;
        assert program(1).op = FSUB_R report "1 FSUB_R Failed" severity FAILURE;
        assert program(2).op = IADD_RS report "2 IADD_RS Failed" severity FAILURE;
        assert program(3).op = IMUL_M report "3 IMUL_M Failed" severity FAILURE;
        assert program(4).op = IMUL_R report "4 IMUL_R Failed" severity FAILURE;
        assert program(5).op = CBRANCH report "5 CBRANCH Failed" severity FAILURE;
        assert program(6).op = FADD_R report "6 FADD_R Failed" severity FAILURE;
        assert program(7).op = FSUB_R report "7 FSUB_R Failed" severity FAILURE;
        assert program(8).op = IXOR_R report "8 IXOR_R Failed" severity FAILURE;
        assert program(9).op = FSWAP_R report "9 FSWAP_R Failed" severity FAILURE;
        assert program(10).op = IADD_RS report "10 IADD_RS Failed" severity FAILURE;
        assert program(11).op = FMUL_R report "11 FMUL_R Failed" severity FAILURE;
        assert program(12).op = IMUL_R report "12 IMUL_R Failed" severity FAILURE;
        assert program(13).op = ISTORE report "13 ISTORE Failed" severity FAILURE;
        assert program(14).op = IMUL_RCP report "14 IMUL_RCP Failed" severity FAILURE;
        assert program(15).op = ISUB_M report "15 ISUB_M Failed" severity FAILURE;
        assert program(16).op = IMUL_M report "16 IMUL_M Failed" severity FAILURE;
        assert program(17).op = IADD_RS report "17 IADD_RS Failed" severity FAILURE;
        assert program(18).op = ISWAP_R report "18 ISWAP_R Failed" severity FAILURE;
        assert program(19).op = CBRANCH report "19 CBRANCH Failed" severity FAILURE;
        assert program(20).op = ISMULH_R report "20 ISMULH_R Failed" severity FAILURE;
        assert program(21).op = ISUB_R report "21 ISUB_R Failed" severity FAILURE;
        assert program(22).op = IADD_RS report "22 IADD_RS Failed" severity FAILURE;
        assert program(23).op = FSUB_R report "23 FSUB_R Failed" severity FAILURE;
        assert program(24).op = ISUB_R report "24 ISUB_R Failed" severity FAILURE;
        assert program(25).op = FSUB_M report "25 FSUB_M Failed" severity FAILURE;
        assert program(26).op = IADD_RS report "26 IADD_RS Failed" severity FAILURE;
        assert program(27).op = FSUB_R report "27 FSUB_R Failed" severity FAILURE;
        assert program(28).op = CBRANCH report "28 CBRANCH Failed" severity FAILURE;
        assert program(29).op = ISMULH_M report "29 ISMULH_M Failed" severity FAILURE;
        assert program(30).op = FSUB_R report "30 FSUB_R Failed" severity FAILURE;
        assert program(31).op = FSUB_M report "31 FSUB_M Failed" severity FAILURE;
        assert program(32).op = FADD_R report "32 FADD_R Failed" severity FAILURE;
        assert program(33).op = ISTORE report "33 ISTORE Failed" severity FAILURE;
        assert program(34).op = IMUL_R report "34 IMUL_R Failed" severity FAILURE;
        assert program(35).op = FSWAP_R report "35 FSWAP_R Failed" severity FAILURE;
        assert program(36).op = ISUB_R report "36 ISUB_R Failed" severity FAILURE;
        assert program(37).op = CBRANCH report "37 CBRANCH Failed" severity FAILURE;
        assert program(38).op = FSWAP_R report "38 FSWAP_R Failed" severity FAILURE;
        assert program(39).op = ISUB_R report "39 ISUB_R Failed" severity FAILURE;
        assert program(40).op = IXOR_M report "40 IXOR_M Failed" severity FAILURE;
        assert program(41).op = ISUB_R report "41 ISUB_R Failed" severity FAILURE;
        assert program(42).op = IADD_RS report "42 IADD_RS Failed" severity FAILURE;
        assert program(43).op = FSWAP_R report "43 FSWAP_R Failed" severity FAILURE;
        assert program(44).op = IROL_R report "44 IROL_R Failed" severity FAILURE;
        assert program(45).op = IADD_M report "45 IADD_M Failed" severity FAILURE;
        assert program(46).op = ISUB_R report "46 ISUB_R Failed" severity FAILURE;
        assert program(47).op = IADD_M report "47 IADD_M Failed" severity FAILURE;
        assert program(48).op = FMUL_R report "48 FMUL_R Failed" severity FAILURE;
        assert program(49).op = FMUL_R report "49 FMUL_R Failed" severity FAILURE;
        assert program(50).op = FMUL_R report "50 FMUL_R Failed" severity FAILURE;
        assert program(51).op = FSUB_R report "51 FSUB_R Failed" severity FAILURE;
        assert program(52).op = IXOR_R report "52 IXOR_R Failed" severity FAILURE;
        assert program(53).op = FSUB_R report "53 FSUB_R Failed" severity FAILURE;
        assert program(54).op = ISUB_M report "54 ISUB_M Failed" severity FAILURE;
        assert program(55).op = CBRANCH report "55 CBRANCH Failed" severity FAILURE;
        assert program(56).op = NOP report "56 NOP Failed" severity FAILURE;
        assert program(57).op = FMUL_R report "57 FMUL_R Failed" severity FAILURE;
        assert program(58).op = IADD_M report "58 IADD_M Failed" severity FAILURE;
        assert program(59).op = CBRANCH report "59 CBRANCH Failed" severity FAILURE;
        assert program(60).op = ISUB_R report "60 ISUB_R Failed" severity FAILURE;
        assert program(61).op = IMUL_R report "61 IMUL_R Failed" severity FAILURE;
        assert program(62).op = ISUB_R report "62 ISUB_R Failed" severity FAILURE;
        assert program(63).op = FADD_R report "63 FADD_R Failed" severity FAILURE;
        assert program(64).op = IXOR_R report "64 IXOR_R Failed" severity FAILURE;
        assert program(65).op = IMULH_R report "65 IMULH_R Failed" severity FAILURE;
        assert program(66).op = IMULH_M report "66 IMULH_M Failed" severity FAILURE;
        assert program(67).op = ISUB_R report "67 ISUB_R Failed" severity FAILURE;
        assert program(68).op = IMUL_R report "68 IMUL_R Failed" severity FAILURE;
        assert program(69).op = FSUB_R report "69 FSUB_R Failed" severity FAILURE;
        assert program(70).op = FADD_R report "70 FADD_R Failed" severity FAILURE;
        assert program(71).op = CBRANCH report "71 CBRANCH Failed" severity FAILURE;
        assert program(72).op = CBRANCH report "72 CBRANCH Failed" severity FAILURE;
        assert program(73).op = IROR_R report "73 IROR_R Failed" severity FAILURE;
        assert program(74).op = FMUL_R report "74 FMUL_R Failed" severity FAILURE;
        assert program(75).op = FMUL_R report "75 FMUL_R Failed" severity FAILURE;
        assert program(76).op = FSUB_R report "76 FSUB_R Failed" severity FAILURE;
        assert program(77).op = IADD_RS report "77 IADD_RS Failed" severity FAILURE;
        assert program(78).op = FSQRT_R report "78 FSQRT_R Failed" severity FAILURE;
        assert program(79).op = IADD_RS report "79 IADD_RS Failed" severity FAILURE;
        assert program(80).op = ISWAP_R report "80 ISWAP_R Failed" severity FAILURE;
        assert program(81).op = ISMULH_M report "81 ISMULH_M Failed" severity FAILURE;
        assert program(82).op = IMULH_R report "82 IMULH_R Failed" severity FAILURE;
        assert program(83).op = FADD_M report "83 FADD_M Failed" severity FAILURE;
        assert program(84).op = FSUB_M report "84 FSUB_M Failed" severity FAILURE;
        assert program(85).op = ISUB_R report "85 ISUB_R Failed" severity FAILURE;
        assert program(86).op = FMUL_R report "86 FMUL_R Failed" severity FAILURE;
        assert program(87).op = CBRANCH report "87 CBRANCH Failed" severity FAILURE;
        assert program(88).op = IADD_RS report "88 IADD_RS Failed" severity FAILURE;
        assert program(89).op = IMUL_R report "89 IMUL_R Failed" severity FAILURE;
        assert program(90).op = ISUB_M report "90 ISUB_M Failed" severity FAILURE;
        assert program(91).op = FSUB_M report "91 FSUB_M Failed" severity FAILURE;
        assert program(92).op = ISUB_M report "92 ISUB_M Failed" severity FAILURE;
        assert program(93).op = FSCAL_R report "93 FSCAL_R Failed" severity FAILURE;
        assert program(94).op = IROR_R report "94 IROR_R Failed" severity FAILURE;
        assert program(95).op = FDIV_M report "95 FDIV_M Failed" severity FAILURE;
        assert program(96).op = FSUB_R report "96 FSUB_R Failed" severity FAILURE;
        assert program(97).op = IMUL_R report "97 IMUL_R Failed" severity FAILURE;
        assert program(98).op = IMUL_R report "98 IMUL_R Failed" severity FAILURE;
        assert program(99).op = FMUL_R report "99 FMUL_R Failed" severity FAILURE;
        assert program(100).op = IXOR_R report "100 IXOR_R Failed" severity FAILURE;
        assert program(101).op = FSUB_R report "101 FSUB_R Failed" severity FAILURE;
        assert program(102).op = ISUB_M report "102 ISUB_M Failed" severity FAILURE;
        assert program(103).op = IXOR_R report "103 IXOR_R Failed" severity FAILURE;
        assert program(104).op = ISUB_R report "104 ISUB_R Failed" severity FAILURE;
        assert program(105).op = ISTORE report "105 ISTORE Failed" severity FAILURE;
        assert program(106).op = IADD_M report "106 IADD_M Failed" severity FAILURE;
        assert program(107).op = FMUL_R report "107 FMUL_R Failed" severity FAILURE;
        assert program(108).op = IXOR_R report "108 IXOR_R Failed" severity FAILURE;
        assert program(109).op = ISTORE report "109 ISTORE Failed" severity FAILURE;
        assert program(110).op = IXOR_R report "110 IXOR_R Failed" severity FAILURE;
        assert program(111).op = FSUB_R report "111 FSUB_R Failed" severity FAILURE;
        assert program(112).op = CFROUND report "112 CFROUND Failed" severity FAILURE;
        assert program(113).op = CBRANCH report "113 CBRANCH Failed" severity FAILURE;
        assert program(114).op = IXOR_R report "114 IXOR_R Failed" severity FAILURE;
        assert program(115).op = FSCAL_R report "115 FSCAL_R Failed" severity FAILURE;
        assert program(116).op = IXOR_R report "116 IXOR_R Failed" severity FAILURE;
        assert program(117).op = FSUB_R report "117 FSUB_R Failed" severity FAILURE;
        assert program(118).op = FADD_R report "118 FADD_R Failed" severity FAILURE;
        assert program(119).op = FADD_R report "119 FADD_R Failed" severity FAILURE;
        assert program(120).op = IADD_M report "120 IADD_M Failed" severity FAILURE;
        assert program(121).op = IADD_RS report "121 IADD_RS Failed" severity FAILURE;
        assert program(122).op = IMUL_R report "122 IMUL_R Failed" severity FAILURE;
        assert program(123).op = FSUB_M report "123 FSUB_M Failed" severity FAILURE;
        assert program(124).op = CBRANCH report "124 CBRANCH Failed" severity FAILURE;
        assert program(125).op = FMUL_R report "125 FMUL_R Failed" severity FAILURE;
        assert program(126).op = IMUL_R report "126 IMUL_R Failed" severity FAILURE;
        assert program(127).op = IMUL_R report "127 IMUL_R Failed" severity FAILURE;
        assert program(128).op = IADD_M report "128 IADD_M Failed" severity FAILURE;
        assert program(129).op = FMUL_R report "129 FMUL_R Failed" severity FAILURE;
        assert program(130).op = IADD_RS report "130 IADD_RS Failed" severity FAILURE;
        assert program(131).op = IMUL_RCP report "131 IMUL_RCP Failed" severity FAILURE;
        assert program(132).op = FSUB_R report "132 FSUB_R Failed" severity FAILURE;
        assert program(133).op = IMUL_M report "133 IMUL_M Failed" severity FAILURE;
        assert program(134).op = IMUL_RCP report "134 IMUL_RCP Failed" severity FAILURE;
        assert program(135).op = IADD_RS report "135 IADD_RS Failed" severity FAILURE;
        assert program(136).op = FMUL_R report "136 FMUL_R Failed" severity FAILURE;
        assert program(137).op = FADD_R report "137 FADD_R Failed" severity FAILURE;
        assert program(138).op = FSCAL_R report "138 FSCAL_R Failed" severity FAILURE;
        assert program(139).op = IMULH_M report "139 IMULH_M Failed" severity FAILURE;
        assert program(140).op = IMUL_R report "140 IMUL_R Failed" severity FAILURE;
        assert program(141).op = CBRANCH report "141 CBRANCH Failed" severity FAILURE;
        assert program(142).op = ISUB_R report "142 ISUB_R Failed" severity FAILURE;
        assert program(143).op = FMUL_R report "143 FMUL_R Failed" severity FAILURE;
        assert program(144).op = ISTORE report "144 ISTORE Failed" severity FAILURE;
        assert program(145).op = FADD_R report "145 FADD_R Failed" severity FAILURE;
        assert program(146).op = FDIV_M report "146 FDIV_M Failed" severity FAILURE;
        assert program(147).op = FADD_R report "147 FADD_R Failed" severity FAILURE;
        assert program(148).op = IMUL_M report "148 IMUL_M Failed" severity FAILURE;
        assert program(149).op = FSUB_R report "149 FSUB_R Failed" severity FAILURE;
        assert program(150).op = IXOR_R report "150 IXOR_R Failed" severity FAILURE;
        assert program(151).op = ISUB_R report "151 ISUB_R Failed" severity FAILURE;
        assert program(152).op = CBRANCH report "152 CBRANCH Failed" severity FAILURE;
        assert program(153).op = FMUL_R report "153 FMUL_R Failed" severity FAILURE;
        assert program(154).op = IXOR_R report "154 IXOR_R Failed" severity FAILURE;
        assert program(155).op = FADD_R report "155 FADD_R Failed" severity FAILURE;
        assert program(156).op = IROR_R report "156 IROR_R Failed" severity FAILURE;
        assert program(157).op = IADD_RS report "157 IADD_RS Failed" severity FAILURE;
        assert program(158).op = FADD_R report "158 FADD_R Failed" severity FAILURE;
        assert program(159).op = CBRANCH report "159 CBRANCH Failed" severity FAILURE;
        assert program(160).op = IXOR_R report "160 IXOR_R Failed" severity FAILURE;
        assert program(161).op = FADD_R report "161 FADD_R Failed" severity FAILURE;
        assert program(162).op = IMUL_R report "162 IMUL_R Failed" severity FAILURE;
        assert program(163).op = IMUL_R report "163 IMUL_R Failed" severity FAILURE;
        assert program(164).op = CBRANCH report "164 CBRANCH Failed" severity FAILURE;
        assert program(165).op = IXOR_R report "165 IXOR_R Failed" severity FAILURE;
        assert program(166).op = IROL_R report "166 IROL_R Failed" severity FAILURE;
        assert program(167).op = IROL_R report "167 IROL_R Failed" severity FAILURE;
        assert program(168).op = FSWAP_R report "168 FSWAP_R Failed" severity FAILURE;
        assert program(169).op = FADD_R report "169 FADD_R Failed" severity FAILURE;
        assert program(170).op = ISUB_R report "170 ISUB_R Failed" severity FAILURE;
        assert program(171).op = FSQRT_R report "171 FSQRT_R Failed" severity FAILURE;
        assert program(172).op = FMUL_R report "172 FMUL_R Failed" severity FAILURE;
        assert program(173).op = FMUL_R report "173 FMUL_R Failed" severity FAILURE;
        assert program(174).op = FSQRT_R report "174 FSQRT_R Failed" severity FAILURE;
        assert program(175).op = FSUB_M report "175 FSUB_M Failed" severity FAILURE;
        assert program(176).op = FADD_R report "176 FADD_R Failed" severity FAILURE;
        assert program(177).op = FMUL_R report "177 FMUL_R Failed" severity FAILURE;
        assert program(178).op = FADD_R report "178 FADD_R Failed" severity FAILURE;
        assert program(179).op = IMUL_R report "179 IMUL_R Failed" severity FAILURE;
        assert program(180).op = IMUL_M report "180 IMUL_M Failed" severity FAILURE;
        assert program(181).op = ISTORE report "181 ISTORE Failed" severity FAILURE;
        assert program(182).op = IMUL_R report "182 IMUL_R Failed" severity FAILURE;
        assert program(183).op = FSCAL_R report "183 FSCAL_R Failed" severity FAILURE;
        assert program(184).op = IMUL_RCP report "184 IMUL_RCP Failed" severity FAILURE;
        assert program(185).op = IADD_M report "185 IADD_M Failed" severity FAILURE;
        assert program(186).op = IADD_RS report "186 IADD_RS Failed" severity FAILURE;
        assert program(187).op = CBRANCH report "187 CBRANCH Failed" severity FAILURE;
        assert program(188).op = CBRANCH report "188 CBRANCH Failed" severity FAILURE;
        assert program(189).op = FADD_R report "189 FADD_R Failed" severity FAILURE;
        assert program(190).op = ISTORE report "190 ISTORE Failed" severity FAILURE;
        assert program(191).op = IMUL_RCP report "191 IMUL_RCP Failed" severity FAILURE;
        assert program(192).op = IROR_R report "192 IROR_R Failed" severity FAILURE;
        assert program(193).op = ISWAP_R report "193 ISWAP_R Failed" severity FAILURE;
        assert program(194).op = ISTORE report "194 ISTORE Failed" severity FAILURE;
        assert program(195).op = CBRANCH report "195 CBRANCH Failed" severity FAILURE;
        assert program(196).op = CBRANCH report "196 CBRANCH Failed" severity FAILURE;
        assert program(197).op = CBRANCH report "197 CBRANCH Failed" severity FAILURE;
        assert program(198).op = INEG_R report "198 INEG_R Failed" severity FAILURE;
        assert program(199).op = FMUL_R report "199 FMUL_R Failed" severity FAILURE;
        assert program(200).op = FMUL_R report "200 FMUL_R Failed" severity FAILURE;
        assert program(201).op = FMUL_R report "201 FMUL_R Failed" severity FAILURE;
        assert program(202).op = ISMULH_M report "202 ISMULH_M Failed" severity FAILURE;
        assert program(203).op = FSUB_R report "203 FSUB_R Failed" severity FAILURE;
        assert program(204).op = IADD_RS report "204 IADD_RS Failed" severity FAILURE;
        assert program(205).op = ISTORE report "205 ISTORE Failed" severity FAILURE;
        assert program(206).op = IMUL_M report "206 IMUL_M Failed" severity FAILURE;
        assert program(207).op = IXOR_R report "207 IXOR_R Failed" severity FAILURE;
        assert program(208).op = FMUL_R report "208 FMUL_R Failed" severity FAILURE;
        assert program(209).op = IMULH_R report "209 IMULH_R Failed" severity FAILURE;
        assert program(210).op = FSCAL_R report "210 FSCAL_R Failed" severity FAILURE;
        assert program(211).op = ISTORE report "211 ISTORE Failed" severity FAILURE;
        assert program(212).op = ISTORE report "212 ISTORE Failed" severity FAILURE;
        assert program(213).op = ISTORE report "213 ISTORE Failed" severity FAILURE;
        assert program(214).op = IXOR_R report "214 IXOR_R Failed" severity FAILURE;
        assert program(215).op = IMUL_RCP report "215 IMUL_RCP Failed" severity FAILURE;
        assert program(216).op = FSCAL_R report "216 FSCAL_R Failed" severity FAILURE;
        assert program(217).op = ISUB_M report "217 ISUB_M Failed" severity FAILURE;
        assert program(218).op = ISUB_R report "218 ISUB_R Failed" severity FAILURE;
        assert program(219).op = IROR_R report "219 IROR_R Failed" severity FAILURE;
        assert program(220).op = FSUB_M report "220 FSUB_M Failed" severity FAILURE;
        assert program(221).op = IADD_RS report "221 IADD_RS Failed" severity FAILURE;
        assert program(222).op = FMUL_R report "222 FMUL_R Failed" severity FAILURE;
        assert program(223).op = ISUB_R report "223 ISUB_R Failed" severity FAILURE;
        assert program(224).op = FSUB_R report "224 FSUB_R Failed" severity FAILURE;
        assert program(225).op = FMUL_R report "225 FMUL_R Failed" severity FAILURE;
        assert program(226).op = FMUL_R report "226 FMUL_R Failed" severity FAILURE;
        assert program(227).op = IADD_RS report "227 IADD_RS Failed" severity FAILURE;
        assert program(228).op = FMUL_R report "228 FMUL_R Failed" severity FAILURE;
        assert program(229).op = FSUB_R report "229 FSUB_R Failed" severity FAILURE;
        assert program(230).op = ISTORE report "230 ISTORE Failed" severity FAILURE;
        assert program(231).op = IXOR_M report "231 IXOR_M Failed" severity FAILURE;
        assert program(232).op = FSUB_M report "232 FSUB_M Failed" severity FAILURE;
        assert program(233).op = FSUB_R report "233 FSUB_R Failed" severity FAILURE;
        assert program(234).op = CBRANCH report "234 CBRANCH Failed" severity FAILURE;
        assert program(235).op = IROR_R report "235 IROR_R Failed" severity FAILURE;
        assert program(236).op = ISUB_R report "236 ISUB_R Failed" severity FAILURE;
        assert program(237).op = FSUB_R report "237 FSUB_R Failed" severity FAILURE;
        assert program(238).op = ISUB_R report "238 ISUB_R Failed" severity FAILURE;
        assert program(239).op = IROR_R report "239 IROR_R Failed" severity FAILURE;
        assert program(240).op = FMUL_R report "240 FMUL_R Failed" severity FAILURE;
        assert program(241).op = IXOR_R report "241 IXOR_R Failed" severity FAILURE;
        assert program(242).op = FSUB_R report "242 FSUB_R Failed" severity FAILURE;
        assert program(243).op = ISTORE report "243 ISTORE Failed" severity FAILURE;
        assert program(244).op = FADD_R report "244 FADD_R Failed" severity FAILURE;
        assert program(245).op = FADD_M report "245 FADD_M Failed" severity FAILURE;
        assert program(246).op = IXOR_M report "246 IXOR_M Failed" severity FAILURE;
        assert program(247).op = FMUL_R report "247 FMUL_R Failed" severity FAILURE;
        assert program(248).op = ISUB_M report "248 ISUB_M Failed" severity FAILURE;
        assert program(249).op = FMUL_R report "249 FMUL_R Failed" severity FAILURE;
        assert program(250).op = IMUL_R report "250 IMUL_R Failed" severity FAILURE;
        assert program(251).op = FMUL_R report "251 FMUL_R Failed" severity FAILURE;
        assert program(252).op = IMUL_R report "252 IMUL_R Failed" severity FAILURE;
        assert program(253).op = IMUL_RCP report "253 IMUL_RCP Failed" severity FAILURE;
        assert program(254).op = IMUL_R report "254 IMUL_R Failed" severity FAILURE;
        assert program(255).op = IADD_M report "255 IADD_M Failed" severity FAILURE;
       
    end;

end cc_opcode;