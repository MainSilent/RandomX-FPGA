library ieee;
library std;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_textio.all;
use work.common.all;


entity dataset is
    port(
        clk  : in std_logic := '0';

        addr : in integer;

        r0 : out unsigned(63 downto 0);
        r1 : out unsigned(63 downto 0);
        r2 : out unsigned(63 downto 0);
        r3 : out unsigned(63 downto 0);
        r4 : out unsigned(63 downto 0);
        r5 : out unsigned(63 downto 0);
        r6 : out unsigned(63 downto 0);
        r7 : out unsigned(63 downto 0)
    );
end dataset;


architecture behavioral of dataset is
    signal data : regt_r;
begin

    r0 <= data(0);
    r1 <= data(1);
    r2 <= data(2);
    r3 <= data(3);
    r4 <= data(4);
    r5 <= data(5);
    r6 <= data(6);
    r7 <= data(7);


    process(clk)
    begin

        case addr is
            when 0 => data <= (x"7ff858e02ad8f271", x"36980e8ed41f6eb9", x"ff7dd9fe87d212d1", x"db4d552b31374355", x"26f7a38c6ced78b7", x"2c0c58361479b4a8", x"91c9c13d90ff16f4", x"680588a85ae222db");
            when 22361929 => data <= (x"b6a6d108cf002ba8", x"ca9f89e54d196842", x"402b7589ac10fba2", x"429305c8e5bd1c08", x"86b92ef8bd934211", x"f36fb4bae218e7f4", x"aad593e123bf52b3", x"fe2f46e0a047079f");
            when 3353257 => data <= (x"11b22cec623c0141", x"ad4a6cd227876f54", x"a8a78312928f2f5f", x"56dff386da5f9c08", x"0d7675e2f5d0f3c4", x"d3f554499d519f2e", x"490ae5de2cbce2d5", x"f21ce51c0a853377");
            when 16361667 => data <= (x"cb84b6f3f46d3a7b", x"abcd3cccb9654ea8", x"f8defef02c5df182", x"c340b682d290386d", x"556f4ffe9c76300a", x"f9058a960452b07c", x"94e75ae043a03d1f", x"8c0c7e54c0f6f9af");
            when 25730860 => data <= (x"adf42bbd2e389759", x"257a8cf822a82483", x"755450416975767a", x"8a817e0c2c3f59eb", x"aae75f6fba14d72a", x"9d3568baa5f76953", x"3d0e018a59387c56", x"47ed1767f682bdb3");
            when 22260599 => data <= (x"b4c8536f6e5ee32a", x"ae68de24edb68eaa", x"5ae9ee381712569d", x"089369b0df61098c", x"4106c01807051809", x"d96f16b7c1e4d520", x"50b34df805a45a39", x"fe9b820c37878d7b");
            when 638748 => data <= (x"b422d6830566ee19", x"fe66e826cc7d203d", x"87adeaa43e2098b6", x"80d489b2b2b1ddfa", x"ae2204dedaa05d14", x"a2a83faaacfe2ee4", x"86ef0bdc9336bd5c", x"6146b171ec729034");
            when 10587689 => data <= (x"f6ccc956b58cb5d0", x"43c66f842449f2e0", x"23058513401510a6", x"59d3c05aee235468", x"32dd94f069f6176d", x"63020ed6022977fe", x"bd738fe7fabc13a4", x"eabe5aade85fcc97");
            when 27362850 => data <= (x"0b0e47df860f4acf", x"b928545c8b518e8b", x"212f31755016f478", x"bc9fd47fd6d84284", x"3238fd94bcb48f3b", x"282cf9a3b9a7083e", x"d0f5c8f611934a96", x"fe2c2f2b1ef51dca");
            when 13340705 => data <= (x"6509a8dd6bf16f75", x"a2ea5141aba31532", x"e334c918d800b3dd", x"ea32314fd2da1857", x"0ed75c7c826748c9", x"f3b7b10cfa84b21a", x"f428a833a28e528f", x"dd9fe7abd2f143c9");
            when 23083496 => data <= (x"dd218cd25ca06344", x"3be6da4c85d08e41", x"c7f10afe99e42372", x"a021d1663d51bb26", x"dc12e4861940260d", x"ade374d7e2754cff", x"323b85f4a72ea4eb", x"59e38bdaa0e10bee");
            when 29841990 => data <= (x"35f78b8ccd56b85e", x"de75ef3ff8de244d", x"cbd5e5428107dde2", x"f4f48d610799a3d6", x"0f3712dc6ad19d70", x"4a54d989e36a06c4", x"ee8d4f2bc6be7bfa", x"2da5000694275dbe");
            when 20764566 => data <= (x"21690dd0ae1c2dfb", x"832aef3f4c4dfdd8", x"bdd9aa937a7991ec", x"d811939b77c7638f", x"abd89c3c3b95a5b7", x"8f5de18f73cc2743", x"1382df672be863e1", x"59bfd0a2f9ce35fb");
            when 3906883 => data <= (x"84dd2535643d2bba", x"4ee7452a2d9abdfa", x"9c3ea14f0a29a330", x"93e4ca427fdfbb5f", x"ee62344f0d7e8274", x"5c8a46637627e9a0", x"383fd82a3dbc28af", x"4acf2ee5ac8f47b3");
            when 13010091 => data <= (x"8227633b46fa97f1", x"e3a435344eaf7ffb", x"64c5ed453dd3fd19", x"182d4aa99592d028", x"b95f6f7e32d2a847", x"05ab612297f4f58d", x"6b59ef4b6149df1a", x"7d8e8f8df70b1f52");
            when 2560923 => data <= (x"d235c7bbfba4ebf0", x"97d5f6eef50d5559", x"a1c4eb7a0edccc22", x"d99c2128c810a238", x"398ed9e878d529e3", x"b3fe271541f43193", x"53e5855658d83c61", x"325dd9c2c47e7453");
            when 10100537 => data <= (x"9974c1b553b4ab26", x"ce11f61e47021e85", x"83250c97f897f1c0", x"dbcd06391f0775ce", x"78a2de4d1ac2f1a9", x"71bfd53eb09252ad", x"da6455ca61d33aa2", x"1750f197b305683e");
            when 29464686 => data <= (x"e36e501361a04884", x"2389bb25e8d96c8d", x"a1183e10cd9b6fd0", x"e628fd93d865312f", x"519ae3d1078c454d", x"19c99ad8b16800a8", x"1922b1c4063d4894", x"95dc250bad51f7b8");
            when 21067388 => data <= (x"66585cbb163918d7", x"fd4b862702a526d3", x"80deaf37f1b34db5", x"c8558074ffe0eda6", x"23424d3e2b62aa66", x"9ca5a52c8c376b5e", x"9fca76356b2f4a2f", x"3b0de88d1b25eb85");
            when 26083543 => data <= (x"4f81cdf745988874", x"ce1fadd9cf0aad5a", x"b9fddb582a42e4a0", x"61116284d92c392d", x"3f9a2065a540fe87", x"4bfb644f05377f66", x"55eb7aef815728a9", x"6b7853e4d4112302");
            when 29223637 => data <= (x"94f6fede7fd4ecb1", x"88630e234ab28b81", x"d60ab4c8f220c954", x"acede0cd2b938cff", x"6715b286b3c06e03", x"1fc286f7a748be19", x"b0c9a29e222071b8", x"c3477c69096452fd");
            when 30438012 => data <= (x"c8b2e2519a6121d7", x"994ff65009b6c58a", x"b3ed9b32572d610c", x"ca0d9f25bbef5b29", x"8154890d09cf5d38", x"19b9dae960ecf4bd", x"39dc7203d79889f2", x"535fa35a32ac16b8");
            when 1954482 => data <= (x"6a632dbbfc0cd531", x"f8f13354ab731c27", x"bdad3b3e4311c4f4", x"b5efbb3d63e1504a", x"b1c8525fea64d1cd", x"6641d37d8b2581ac", x"f3cc2fba6369937a", x"9d90ad0cf08297a7");
            when 28589478 => data <= (x"f8011c494c71436f", x"d8a08ee7d0e03e18", x"ebba1f6589390107", x"b8ee796683b13cf8", x"a417cd3ba943ccb6", x"74172644b7f1b4b4", x"560ff40b79cd2f90", x"98e052868227f838");
            when 7147741 => data <= (x"8f409e49edad24d1", x"d7ab305e4af03f60", x"8eae74b62ca05615", x"a169d5aae7cb8506", x"4ff9394a9800d20e", x"a1d7740d67e3675d", x"ee4cc224d211d2a3", x"0561468809ea533c");
            when 8541261 => data <= (x"616c5770831289b2", x"016ef8dc6ec37852", x"fe825c2f82a616c8", x"c96f6758791737fa", x"d40c5d0deeba0ed1", x"7be65bdec61faecf", x"b7f2cfd84b8d964d", x"264e9b89dc11456d");
            when 12524790 => data <= (x"ea43bb07981f3fe4", x"cab9fb2be1f5847e", x"277dc0dd9e5e08dd", x"a4455fadab6962ca", x"0eb9d9724cd0e082", x"fca6ebffa0ab67d9", x"fa7734529e81a793", x"30d6c33533e28e5b");
            when 29630525 => data <= (x"be7c5a7b32e7a39b", x"7912cdd3098c3557", x"5da0917a4887ba8a", x"51cabb87745983c0", x"19d8f6489fffb22e", x"63ec666a143900fd", x"9de9a2f2978d90c1", x"ae7e2351b06f1be0");
            when 10828145 => data <= (x"04ec6676953825f7", x"1eb064bac3d405a0", x"63ea789a75a6e7c5", x"6150b4382aaa16ca", x"a58546da971a242b", x"120d30876c61655f", x"9915aa37b97777d1", x"3fc05a35b4c4199d");
            when 4836230 => data <= (x"adfd1cbd0e841257", x"443ba044ffd352dc", x"88838f873b931237", x"1d30000894539c8e", x"223c32e75bd183c9", x"996576cad074dcf5", x"96ec255a19df0fde", x"1b5c1b4afd977a20");
            when 20934055 => data <= (x"1aa9ffb92bcf3df5", x"9cfd9f3c56efb110", x"0f9315f191b0fd95", x"48d7d009053c6875", x"655ed422067529fa", x"24f9037c0b13b9c5", x"4567e75dc57d435f", x"21024d55ded9ac0a");
            when 20246876 => data <= (x"cde823ea2e3bcffe", x"99847808f850f93f", x"908bd9b42d43f7b7", x"4a5223b70cc4c340", x"e83a846788bd04bc", x"efc5c9354ffd6d40", x"6bad5d1f5037858b", x"361ebadcf4361c3d");
            when 9969635 => data <= (x"12894ddda7294c2b", x"075d62dd5eb2d37e", x"3288df65216e20be", x"bff3d7a848d18855", x"db986febfdd49d64", x"0b8616620614acb7", x"34f478fbf31686f5", x"8ada3ea7b09f8ac9");
            when 13479743 => data <= (x"295c481a33721fa8", x"99070c83332e3655", x"fb6c82f0f134ba2d", x"dec958f9971c0da0", x"8cb41bc115d1c882", x"072511932ee1a0e8", x"0883ed6d69e45832", x"d6178eb428d1a774");
            when 29633621 => data <= (x"dc87e5733953d9fe", x"59e55ecd6df799cd", x"4f90844c24c74652", x"d4b0649f729bb29e", x"0e8b7182d50ed8a9", x"2c0b6ea1b2145f47", x"429e14ac71203653", x"5c3a753a30a4061c");
            when 8759488 => data <= (x"b36882fddd73fdcf", x"3ae293fecf1f6a5f", x"2cdf642f4adfc4cb", x"ac9c12be6533b81e", x"8d5d95035c1993b9", x"8d8ddaa9307311f3", x"a6e9b691b41f92d1", x"19f96c009326325a");
            when 1371113 => data <= (x"b9e2992e2c008674", x"73c3abaebd72ad74", x"3a12af24f6d409b1", x"1503098a5b63e207", x"e751e4a6ee273f0b", x"2732abc05e527681", x"202a3cc2c8d581e2", x"35c174b4017430ed");
            when 13584192 => data <= (x"1d64c256ae611790", x"7870e77da5f2b732", x"5855364bab494d88", x"da7f9e1707ca327a", x"4297d7a2b72b87ec", x"33d16bb554d2627d", x"3ac9a3c37d9f2a4b", x"61eddc50bff3f495");
            when 29162742 => data <= (x"a8c69cf13de3cdcb", x"24fde7155135a619", x"1b8cb219dde61ea6", x"2b2fa13a65675cee", x"198f339906d6b06a", x"c25f02b96242310c", x"01a54793772d7eea", x"787e432756534b0a");
            when 18250615 => data <= (x"1d6cb328934e64f5", x"67614ac5f48d0eea", x"0db525cb4225ddd6", x"bcefbc865b3051ce", x"a68813af3ec91c02", x"cf05846336815244", x"f337e8ea1e4e3e77", x"daa069678a5ab2ba");
            when 20022964 => data <= (x"09a50dc6dc0e2d11", x"608fdf847b6bee6e", x"32a48ce0935fae84", x"7a0ccf6b8a8459c2", x"93613c5a2467f450", x"58539137250b9cd9", x"8af4d446f4b75439", x"35cacb9418ae2989");
            when 19050661 => data <= (x"2e1e2d05f1b16373", x"74b51d6e37542dfa", x"52c90d9485ce32ce", x"c8a774918d2e3bb9", x"f32a9ff133bb64e6", x"1188d32779fe209e", x"05fee2695da556ce", x"d403a0e06c0d3e69");
            when 1055486 => data <= (x"821742c31833f942", x"6bf1a69fd0df74f6", x"141dc31a67e04a2f", x"7bf6d32c7e45497a", x"4839ea0d0fef388c", x"80521de703cbb895", x"bd0e5914b384ffcc", x"45714a1cefa25bfc");
            when 21226371 => data <= (x"56bd43884d582d0a", x"aebe0eb28c985dac", x"11a4260738638b6d", x"d5508a27208f9cfa", x"2ecb9e41c1a4705a", x"4ffc51a64d93ee01", x"56dc725aa0721402", x"b71904b5e10a313d");
            when 21516961 => data <= (x"527110300110d669", x"1bd87d907677198f", x"a682d2d2171e610a", x"0c4d40290e97925c", x"d90bad10f494fe7c", x"1d22051110ec1c7c", x"b6a70cf8ddcde80d", x"8456ad9a7ee42b62");
            when 2261468 => data <= (x"78d558bbb07f5a50", x"9da6f37afcadc07d", x"e655d46da329b2b4", x"38c22a5b893b0b2c", x"0d7cee0925d2c426", x"b75ce04d95fea0a8", x"1dac01f2900b1912", x"d98ec7f6cc246f49");
            when 2687377 => data <= (x"b2be1df741ef7d67", x"4fac3437d85216d2", x"896c04a214aec829", x"1c85f2f5cab41e89", x"8e7d771d7c89d451", x"7e826308a6fa1bdf", x"6b221d38ba37beb9", x"3949ec8d212303e3");
            when 17664291 => data <= (x"72640fbd88134c95", x"881d2608a650bf6f", x"5538f3fd7d0d95ee", x"e423551aa87ce633", x"90418c00bde8144a", x"add5a8027f865bb6", x"85716422a64184b7", x"93a0c5b8ec7e012b");
            when 10419439 => data <= (x"af27b8ae2128d69c", x"3d15d9c3a2c73aaf", x"c4d9bf7406390cc3", x"06471d31f2ab7398", x"9b0f4a9ee460e993", x"d99c6de68f2fe840", x"42559b9b78141687", x"d0ab538536b0439f");
            when 17362084 => data <= (x"f70feb75a35a79e5", x"13ba5518cbbc59b2", x"abf456d3c84d1fc1", x"26122e1252718c12", x"3b82cb2145b21001", x"73241958f3efc840", x"271674024cc762d4", x"77084e31746e8213");
            when 632961 => data <= (x"15ca0b55f4e59ed2", x"97c68f2fb576ce41", x"85696bf8c191d9b8", x"802c7b9b2ffae6b4", x"d81ec56d54a08f85", x"bf8e4b2f1831cb8e", x"4953a5e0c484d444", x"3efd91ec1ccda000");
            when 9880244 => data <= (x"85f920548f6131ee", x"fdfa9863ae229e56", x"74bc968a5a7ae6e8", x"6e756a2c70158183", x"0a024cf5f56a09f6", x"43f348f88f16cd36", x"b938f47f462b113b", x"5bb33f80033907b0");
            when 15328100 => data <= (x"23e4a469a82cc894", x"6c9450336c1d0c91", x"053593e3e8e70a16", x"42074c8cccc04ddd", x"2f50cbc0e1fd7f59", x"efafaa6398eb196c", x"db5286ed14b0be6c", x"c4ec782acf057aad");
            when 20646470 => data <= (x"180a0a7c3fa79058", x"c07951daf8208d9b", x"f07b8535b1dd2dad", x"263c32b6e0c19838", x"f5b2f7560eb81a1d", x"7587cf27b4d14d1b", x"7c7756b9388e480a", x"5e9079f951a0f829");
            when 27181809 => data <= (x"c0f50d5d5f0da916", x"f8d13a548df1a3a8", x"436a8df35ca6a29e", x"618aae5ee4439c62", x"688b2ce5238cfd4e", x"8b07f9d16b426e16", x"b377f4298ea8a53b", x"16c4666948511e41");
            when 28646097 => data <= (x"289eea493add8531", x"7b1c51d4c613a68e", x"f5eca9e45f452328", x"f36fd6b634ce1ea3", x"95890fb292f650e0", x"70e2c3be5742f0f7", x"7d86bbb3326454e8", x"4c6b00211d665b8e");
            when 28050641 => data <= (x"3157665f915ead36", x"92ec3794197acd9a", x"bf9cdcff7a24ea39", x"999817fc7aa87d4a", x"366f77b08c29110c", x"e1175ce97d02d4d2", x"3c60d9b0b0926c3d", x"49fb1fb1b39fde14");
            when 5040648 => data <= (x"b476d06755dc954e", x"2709386ee4765eaf", x"537f76611ecb7795", x"c27cbef7a1eea02e", x"1f377e1f11da7c27", x"41c0aa59959a5c4b", x"556bf93ee1388c8f", x"2a722badec5c9f1a");
            when 2048226 => data <= (x"e86ecc929af51da8", x"368e6fb31a34e9f4", x"8fb6b97bbb4a493b", x"507c580afe127d6c", x"e0d56adf55e010fd", x"3753ecd263a3a520", x"f62f0c0bcd0a2eda", x"e4c044eb58f75ee1");
            when 5733990 => data <= (x"7017a46c2b134d26", x"81d4784a261babc4", x"4334e39702ac7a0c", x"809c3923b9c4c3a3", x"cad334ebf51b4922", x"21e12e4f9a549870", x"de9472061eb9d2ad", x"2e83a0e91b1532fa");
            when 4771645 => data <= (x"f2798a889f8c7b53", x"b32ca93d9d91b7d2", x"499280d771228f41", x"fafbbc23473081e6", x"f19e2c2599bf62b5", x"b395ece8541a1f4a", x"c5f467d36a4d1d4c", x"16582220e4d9b9d8");
            when 8577776 => data <= (x"9a5721770c82a17d", x"d8d7259e0e2fd2fc", x"893dc81d8677c0c2", x"3ec3e507f38c3baa", x"b7d01d3f0b68f784", x"d328ab2c21b8da2f", x"4fcc619f014a71a3", x"8c8c143610edf9d7");
            when 15232546 => data <= (x"ccc2af9416eb9be1", x"002c829f290f84ff", x"5576e754292bd7a9", x"b7340e1b66f74c3e", x"9e2a6497dd199dba", x"f557f3addf556727", x"44ace8ad41f49898", x"25bdc4f231e1539c");
            when 7253742 => data <= (x"f220354958779614", x"86e433aa40a17f4a", x"bd32211c63b6a9fc", x"f1e6ffebc5a16a05", x"056f86b67d4270e5", x"e455f2b3000251a2", x"f466dec762c8298b", x"1fe7a73d222e6242");
            when 1380700 => data <= (x"8ac54f4982930997", x"c5ad3642ac57b8ea", x"a3b1133e2abb8451", x"d34cf5b1a5c24922", x"6c2b5d664f368a9c", x"8fd411c6e32b35bd", x"2010ce8f514ae4a1", x"d47d481aa542bbad");
            when 23251781 => data <= (x"7616d706f04f344f", x"88bc9d0ab9cdfce4", x"015dce65665692df", x"3cbb425bc4f00a93", x"3ff0942b335037c2", x"cf5b6d08b6d0b1c5", x"f44e248284253ff4", x"f0056c7997e44943");
            when 12014830 => data <= (x"db66a9febbd7e8fd", x"9ea3f5f99b44e35c", x"035069e9f909be04", x"08b601b368bb6f44", x"cab30d4483ea386f", x"410a6a8f3c4f24e5", x"3addef6baafd72c3", x"539378cd81abd2db");
            when 23343042 => data <= (x"4f49113029aa8352", x"02512a40ca54214c", x"66a7e0a7b23a981f", x"d2051fa19bd19d71", x"40c78c18ffeb9049", x"bc10f5358d50be68", x"3d79c5d6032ecab8", x"e55d61da1637b869");
            when 21922192 => data <= (x"4cc854b152471602", x"360714f1e17ef8aa", x"3b07832f95208075", x"ea997f4a7d193d2b", x"0258347eef205032", x"bff759662b935107", x"b55d60b8c9d70934", x"1d7b604ca86094ac");
            when 21189794 => data <= (x"b498ffe5d3b871b9", x"b5f37e53ea304fa0", x"e13d6448ecc3b25e", x"f897dce526ad277b", x"245ab8deb0691d54", x"57311bff2a53d5db", x"13eca56973d11f58", x"f21a6b40c365a456");
            when 12772675 => data <= (x"0f4cadd7d6c6d261", x"4b29be3e1e2bcaa3", x"474f21c1b3131e19", x"ad959f8ed4dee503", x"eebb9663fa02459f", x"2775d96a6211b811", x"ce7f5b4cd55e95db", x"73172e565fcd4f56");
            when 29364624 => data <= (x"8f3f66e1264d41f0", x"0a0c9438e60a2c5d", x"4d6ac045a4202956", x"551301d7b94785f3", x"270e4893ed96bbc7", x"cef160579d2ccd07", x"2fe20e6793b6e10f", x"3f646e0f21318c97");
            when 23770903 => data <= (x"ae40d013b7d2f7d1", x"6e2bce364f776124", x"389b7df4642bac78", x"9602328a23404813", x"6523c806e295600b", x"ab5e3c8b34849ef4", x"f701b2e95441f425", x"d93760491d03b755");
            when 23480835 => data <= (x"3206f47421f124b8", x"c8af482f6b0aaba8", x"4618936c6109734d", x"eea0a0023c4f70a1", x"7f91603e8ac54cb7", x"6f025f9ff11561b0", x"365ccdd6dd0f497c", x"e6bd738b5ec36f1a");
            when 23760574 => data <= (x"974ff8a9bcdfe368", x"ee8fbfd0442b4131", x"75e4b8fd4c43e8d5", x"5fb23fd37abd7df8", x"20220cdd6c3f0dd1", x"fd8a98081b7e2289", x"36eb479e315cabf2", x"c4724b24e6e520d6");
            when 24078763 => data <= (x"c5f69144b8261c3f", x"92323f25d94184ad", x"09bf442739263d94", x"d7e7a7ae89327a03", x"5cc2295583c4eb7f", x"c895860070482aa7", x"1cfc559c31e42d7a", x"0b2a6b35d864ba38");
            when 31313356 => data <= (x"2802870fcf5a0c6b", x"300a195763a6d652", x"53c8f2a80a147bb4", x"5a1b2700dffc44e7", x"f2a967ae7f09c0a0", x"57732a3d85a04971", x"063137de925627b4", x"4308fd3692581c2c");
            when 10135013 => data <= (x"de1ee100fa36b2d9", x"69c0652e62ac2512", x"4b264cc1b495561e", x"caad69388f781054", x"e8de96442a19424c", x"32c6a19f44098d47", x"a5eedde51d17d4d8", x"783e50c38c666139");
            when 21823870 => data <= (x"26a9cb2b652f6a26", x"7605a529bcd5479b", x"c967a6de2274f0d6", x"741c384a8dd9a316", x"cda9a8a14cd30e04", x"1705c43814268043", x"ef79aab38f769486", x"60976c53fb0250e3");
            when 17471869 => data <= (x"18960923764f756c", x"0320b326d81e3634", x"78057d812355eaba", x"b53f018087221aff", x"5786679cfad10c1a", x"2f7e8f7d14912da5", x"b98c63fede23e52f", x"3833f8466cba5c2c");
            when 32183550 => data <= (x"324ecf8b05c7a21f", x"d33c2855b541300d", x"bcf535e3eee0b00f", x"eea3531e23558de9", x"e6b59aecc94c0f1f", x"8d7a4b43fdfe1962", x"a0e7928e0530896c", x"3d504c540d04d14e");
            when 3643263 => data <= (x"275c0a9e2600c72c", x"d88a1d2fa9ad4a06", x"7191f5d7997634fe", x"5d9b20741b47de3b", x"19eb13a75a6a99d7", x"ad21c98e1494485b", x"a7b22db19e2cef85", x"9419c4ffdb792430");
            when 17778486 => data <= (x"731d43e022e72637", x"f9a9917b96bf451a", x"a4895583f7391ff6", x"44e47072b05c7bd7", x"0f11e7161237b86b", x"53a1a589f2b07843", x"b678de3fc036b5dc", x"e2b4bc542190fdb1");
            when 27105305 => data <= (x"f50d42d32a85eab7", x"d6611435ae288b35", x"d5bfe3ee7367c113", x"3d01d5abef1a7f92", x"5a4ff22af4e179a8", x"420ed72c3e5baeac", x"76d3ca4ad100e32f", x"28fd3ffd2f766435");
            when 29456092 => data <= (x"7d6d58789184a49d", x"5391360faedea7d6", x"c5da2d38c61bebe4", x"59af3184854ef7f9", x"d63dbc9c0390f431", x"0bb3b9512d3292e2", x"c77cc0834ca16439", x"d91d72b258c4394d");
            when 26538772 => data <= (x"34cb748b25398d01", x"913b5e39af24707a", x"a5ea334cdb27c9e1", x"b16a494dd18828d1", x"84b62096dec8d7af", x"662ac7402b18ef69", x"08e29a3cda5b85bb", x"e4ccb9ada80cd5e6");
            when 32070135 => data <= (x"48bad3892e5b1e89", x"8d56ed64c464d907", x"93e3a46d6351b2cc", x"b976b3ceb257b013", x"bf0afb83310bf822", x"cb9b7c1cb5ef5317", x"98d070424ab7d3c5", x"125e5845ac35d137");
            when 19183100 => data <= (x"660c2d1275da0e0a", x"cd968d11ee342ecc", x"45120c193bbdbcd9", x"88b3faaef0fc8447", x"ea52f01e4499e3c1", x"421d5dd0dc8716f1", x"0bcc1c7a809f2871", x"679f4908f69ca3e8");
            when 10813942 => data <= (x"9eadd1fac7f8cd1d", x"c03d3a8bc442ebdd", x"c98187b2fb69676c", x"8aa1f27ed5d208a0", x"01b385622952ecfd", x"224ef944b07868bb", x"f42ada9f42d2c22c", x"06d18ed22c885398");
            when 15068647 => data <= (x"0967c4aff648d251", x"9a3fcae014b6e097", x"4bc9d53a16135a1a", x"1ac13a53b8e3b555", x"4a5a87d25499e455", x"e69bf881e5d66be1", x"683e58c28c1cc202", x"83c469c8c7d8f475");
            when 6640067 => data <= (x"344c084bc1ba5fa9", x"2209a3ab27d8602a", x"6eb2ab5dda93af71", x"22b3bc1531f1febd", x"6b17dd6997424745", x"04edb94ca3d95bb9", x"0fb612ec86a2548a", x"9bb5337958270622");
            when 31592091 => data <= (x"954520424ea2f835", x"85433b4b4a8c5d76", x"3142f061509166d1", x"2e4b573f74fc976d", x"fd10628fa1fe6625", x"f6efc56890215e1d", x"0ae79bd9d925c78b", x"ea1600e0cc558b45");
            when 33039919 => data <= (x"1c560d94fa8db109", x"a05118b3de932f68", x"02ca9cf4c54c8125", x"1c2966b964dcd9ff", x"c43018beeddd7b94", x"0165c31d15ff94fb", x"8fdade627ce44907", x"50b89925dd2ca5d0");
            when 10472748 => data <= (x"28d6ffbd6822dc60", x"40135a71b3073ff6", x"bf24a1fd908a6723", x"27192ab669809484", x"cb51dcc4ff94af69", x"8559dc9473e2587e", x"0d4e3d4bb47ed5b8", x"dc308907021b791a");
            when 3450861 => data <= (x"e084319077f5132d", x"f5470e489aa8a03a", x"adf95338b8d5930f", x"1ed34660ca963ccf", x"afbe5d5792e4c9dc", x"58b3f9d3cd2968fa", x"70a83556e255e4f3", x"6d156f9624893157");
            when 3450863 => data <= (x"35eb38e0d7daa09d", x"d68420b8e22dd26f", x"dcaff5ec3da15e37", x"1ca23b0fa10f8909", x"d3d5f8aa8f7b2c6a", x"93ae497cd4496d1d", x"6b04a2b1f76d39a0", x"9fe00301b1f104d0");
            when 32102189 => data <= (x"0349dcae39f6b0e3", x"1d8450841d9550d9", x"7b52866b14250307", x"2bed85be2a4575a6", x"36848cff0496d97c", x"8288e141d2aa4084", x"84c5f05e6823ba23", x"fd7fb92e90fbe680");
            when 28863704 => data <= (x"6bc1a112b7933eae", x"ad761040e330768d", x"7ba763d3c79ad3b0", x"53e8217c587adca2", x"2552eb2226460630", x"6b58fbf568808fe4", x"39accb13a552d587", x"26c2cdf5d7069baa");
            when 4932723 => data <= (x"209d2a652c0fbaa6", x"97affecd31dca327", x"e9efa7d557ca587b", x"ce18fcd119573d1a", x"fd425b5e847682c2", x"4c3691e84d959365", x"88f0a0fe7d0656e5", x"6620c734eea8a62b");
            when 4156571 => data <= (x"1bde3161a3fba685", x"a47fdb74b531ffd6", x"ee5777ee112e20a6", x"bd7892627fb9845a", x"e3d2a2bcdf567e84", x"048789922c85d732", x"9c84441c4fecee04", x"ab71579a995b9f2a");
            when 5415288 => data <= (x"2e8d08453635ded4", x"20c465a5ba81d2e6", x"04d3f246d81d5d6a", x"3d2705f3663c86c7", x"8a5f9fef8392ce7c", x"e9e3181c4520413f", x"85f018a17b5991cc", x"da34d7a5137582e8");
            when 33329163 => data <= (x"5f8946b35b5e112f", x"0c96f121c3c40aa3", x"17ec9488b93a79ab", x"65d8e715fe460720", x"cb92256d443e7aa3", x"52d92124bb97a436", x"5d1bca410c42eeb0", x"387b76d64d600fe7");
            when 7483845 => data <= (x"76ad44c01cf248c3", x"c18b4e25a730e881", x"3b5cec4f9f393a66", x"3fabfc77b05ba527", x"eef8d3cfe0a78ef2", x"26afdd9dbcf245f4", x"21f652918a305ad1", x"4d804dea13951f08");
            when 18429247 => data <= (x"bbdf5db48230ac1d", x"d080389455e2a645", x"fc338b422b893fbf", x"4cc9c53999dfff38", x"24cc0fe55f027856", x"1a304761baa28025", x"c4f279e005441084", x"25318e1baa797e31");
            when 7672120 => data <= (x"e5acf35bedbd956a", x"7f3bbefd88a89f4b", x"02b75fca916a83e8", x"0ce97a2662b1626c", x"c6bc5d9d2115a35a", x"5d19df6dbb64646c", x"0935e1aefa372ad9", x"951e50311d9c6256");
            when 33905733 => data <= (x"b8e59fe0951ef190", x"632ab19a58a08558", x"2a86706c368006c9", x"c76212ddd37105b5", x"8e7954ba94d574ab", x"05d81bafbbe0a07c", x"4d003035b16270e7", x"5adc8ab654bbc792");
            when 26038976 => data <= (x"a1b47da7edb9942d", x"500874a8b77c6cbf", x"b031c3626b38fed6", x"8575986312a6c7f5", x"2ab78afa564c9260", x"2495e1273e3ff98e", x"3ce4eb14db0757a5", x"28384824bd726a89");
            when 4668363 => data <= (x"b1dd3bbb809c69e7", x"7531dd17b91d0e5e", x"7b842698292b2627", x"6df719920ae6af06", x"8648578ef7068707", x"ae7d0fa1f338956a", x"b79d838e1b4b0882", x"3fd2591335cfb098");
            when 840749 => data <= (x"d2613c67f22e0844", x"1d5a245095fd5640", x"85720c7c0069b9d6", x"3ccdcb09b9e3a59c", x"3c01a216280af49e", x"4720aa5b264ee6cf", x"4a7f7d4d9d422796", x"4731a6d3213d48f3");
            when 22959671 => data <= (x"4be0ed56d1970efa", x"17d94c1ae2322c32", x"f7dbfe63019f96b6", x"900ffa18331f810a", x"36bce9f8f8f21c0e", x"339be7da379d9390", x"7383af9d527f7008", x"149c96fbb666b437");
            when 29368471 => data <= (x"ecdb2924eb8124a0", x"8eecc36f08cf0156", x"c148d38897c142df", x"13514c24eeadc3c0", x"65b805b609b1c960", x"c7e72d9569af830f", x"c238787048cd8f10", x"9b5ad1a075d49abc");
            when 15883060 => data <= (x"1c74e352a9cfc3d4", x"982417eccf924182", x"beb07b676081a6c5", x"01c436630b1f104f", x"400cb9bdb68fa25a", x"7d129e70aa427af4", x"f19f885df6995a24", x"7ac22b9f41f80dc5");
            when 14402863 => data <= (x"f586120f0c967e05", x"a87868e4cc7e9297", x"74062c0acc285820", x"9c01d2985fba04ec", x"8c3b17c83c3c4550", x"b4f7e09978881bbc", x"e94a42180a71a860", x"18d051c63a00bf7b");
            when 33647126 => data <= (x"18e471d277b9a2b8", x"a5f3820a85ed11a3", x"0eac4b8e413f90a1", x"1273da542639c494", x"9a0fb4c9c335047a", x"6e57738f9efa710e", x"e491161a644cc4a6", x"b19b9679d7da941b");
            when 17689900 => data <= (x"f4436afc1c6231cb", x"0bb2b8a84448573e", x"063ce3df67b9fbf8", x"a373564f1f39431b", x"4ba6158ef2c26d9d", x"baf67d9022b421e3", x"5e72f56ef5179e26", x"dd382bbd955d3cf7");
            when 24894715 => data <= (x"805262f536b97b1a", x"113a5e59fbcae13f", x"3b87cb5401e8d3dc", x"2cdee23e605cd4f1", x"f28bd87e3f1f76f4", x"e2bef80511ab9389", x"5a57165d2472b96d", x"ad734528c2beef7a");
            when 13380252 => data <= (x"36968be33a67903c", x"9edff0646e78120a", x"9b70ff3ecae80125", x"d496932fa72c97f9", x"885d1e8aef62f020", x"0bb24c3e2a815881", x"d131aaa0ff5e9396", x"474196ccc86e1bbd");
            when 10875030 => data <= (x"6817633723f8779e", x"0f47e99130fdcbbb", x"3bf1735c6fb2bfb0", x"febe69ec0ef92c48", x"59ee2a72a88170b0", x"61abe16c188efdfd", x"2117e7c41cdff581", x"6ccec1cd1e6dcd8f");
            when 20394843 => data <= (x"513a390f07374d5c", x"edc2aee7dbbe5f07", x"4a49fbb514f7304e", x"1f8a884a3bbe9e2c", x"de529daba3203351", x"7c62166ded1e5271", x"3273aa345c3c66b5", x"0e01b5707f2a498e");
            when 29320555 => data <= (x"64d1280f270daae5", x"5f8c7adffdf28211", x"ccbffac0cfa467d6", x"c5040e11da7f5104", x"00b15b07cdfd5921", x"daf9d79a075ee2c0", x"80079618ef92b842", x"941799c5f03edd33");
            when 5071188 => data <= (x"057055c5aae27a47", x"cb5e5be2ff3ae1c9", x"6e9726dd3888d5f7", x"134beaa46b34a75e", x"38615c6560af1b42", x"37b32ddfd3ee9337", x"77352bf3ec8800e8", x"79ad6a0c88be97fc");
            when 4093822 => data <= (x"aa2513b70259ae9b", x"e5b47e231f7a8f96", x"35e71017fe34a691", x"bd7c02c6693c6f4e", x"8817a7076374290c", x"a10f86dffd3cd2d1", x"9bfa804d632b1d65", x"d5ecaaf96ab1674e");
            when 29471501 => data <= (x"fd3f1c40fd45584f", x"c46db0871ce7e403", x"b879864a8d0420b2", x"34f332e017aef048", x"319f8f9e195ecfe9", x"f197e5ed2bd5539f", x"40a96295c03e83c0", x"67cce25af377c8ec");
            when 4897473 => data <= (x"2108212ef04b6c9d", x"e6619314160d0a19", x"f6d3a9ba7fd9c702", x"0f43731c43fb95b6", x"9837b58020216bdc", x"f54ad11223d13c74", x"694960b77021785f", x"1cd3d4dff6b83a3e");
            when 18479866 => data <= (x"99f726e06bb80f44", x"7e93f03b60e4d178", x"e1684c60e9064807", x"9407161773da5256", x"1156107f62dc5fa0", x"f73c88215ff4a694", x"de2efd9e02c62c32", x"c6676b9f9c643788");
            when 16427314 => data <= (x"ec6a913033b2260e", x"bc2ed3daf62f159d", x"5542641f1af73fd2", x"49872947bcb1e946", x"ea15cc104802148a", x"600c7d295edcc991", x"2b93d351da626547", x"40a6445ac07daa77");
            when 32144114 => data <= (x"84463aab89313c5a", x"a61e4f0032f09fc4", x"ab1d20dd6d43b903", x"9acea9c0ed135ae3", x"ebe4832d311b6bc6", x"3f3e6efd15a2be7a", x"5235b08345c7648f", x"945109468075fc69");
            when 2038120 => data <= (x"e8dc7cbe972f9ede", x"0814999bd91fd472", x"7c99877d94772152", x"8d22ef5d8ab8da5f", x"619f630de6981196", x"da2ed54c68d2e683", x"608e51917d004fc7", x"e8b353a96483449d");
            when 17943524 => data <= (x"9315a3fdf56698c0", x"438528dcba2b7b58", x"d7e884af73e11095", x"0310c3e63ca3b333", x"946ac3d3832d5b07", x"ef0eed8ba99f312a", x"a86e2d029e9ecc2b", x"bde405561ac2fd4d");
            when 20519296 => data <= (x"4a5714dd2be23f12", x"58a9342a62e7deec", x"65e0eaa9b8f9335f", x"f3965d9afe244b6d", x"18b0600141f035f1", x"cbe0e80c76372d71", x"1ef62e65919f7a6a", x"7a1141e434f8caea");
            when 18380423 => data <= (x"d44bdcd3fbd3f1cf", x"5872fb793b3195c8", x"def111b2428f2abf", x"6a9c091ab0904713", x"ba6d0c8c2a356851", x"828650d0f9a5d210", x"982de5711aa027e1", x"4ef98e610d07e921");
            when 19262840 => data <= (x"12d6c119d2f7b79e", x"bf0460bfe93b4b09", x"8602f99fc5e0973e", x"a649157263e51b53", x"749a4eb8b67788d4", x"71da1d61a712ed03", x"62f4139a6a936ed9", x"2fe82fc8f41bcc6b");
            when 6019019 => data <= (x"d7bd6438b393bd3f", x"9d1374a8b6bc4be8", x"b1f354864f86ea24", x"1d8e1e3a0031331e", x"49cbbc718b395098", x"5e24d330fb7fa4cf", x"f02a2009c763eae8", x"92ddb58150b915c1");
            when 33191885 => data <= (x"5eec077d88544432", x"705207a21d067346", x"d2fd6d2ee6f776d3", x"c608d466ee3063da", x"74b4e11e788ecaf1", x"ff3e910a82f3853f", x"65ec2cd20e91accf", x"885a0aa6b16508e7");
            when 7230809 => data <= (x"64916fd930068fbc", x"7f3f239be20d48a4", x"5cf013147e93d3c0", x"699dadc6cbbf5340", x"018723913e660f0c", x"d408ba2a17e51a86", x"4956b5f0715da21f", x"dca952f9a10be00c");
            when 8151360 => data <= (x"9a5c18975a5b6cef", x"5bca677b7c1578eb", x"0f7e1417e90aa120", x"fabe6f530b4957a6", x"cbff3e15fc7396e7", x"6bd78768583199b2", x"0693c3ea0935e919", x"d8bc3b23c02f5250");
            when 30062161 => data <= (x"6b433195915210a0", x"35512eb35a0adbb8", x"61b93b2279627cb2", x"efbac1a7ad82aecc", x"d34eecddabc0dc23", x"c3069d310f56f2ec", x"f155cf85345d6815", x"0b130f8f58ee9dd7");
            when 6287027 => data <= (x"f2fd40fc65b7cbbb", x"f2c44bc1902cd24e", x"82141aebe218b495", x"28c0e9232bbd026e", x"795359a07e329361", x"7419ddaacc189881", x"88ff64a6ccf7946e", x"c5b5ba1825948aa6");
            when 29162511 => data <= (x"79df279712a1b249", x"6941e232315838d3", x"3692427df3e8565f", x"13410803d60178ba", x"42ec1068cc391418", x"7195b325ec60b4d7", x"c491cb5440a6fe66", x"6d1da80308725644");
            when 32269559 => data <= (x"9d9249fa9c5dbe32", x"de7f47aee382cc65", x"427fa5502eaafe59", x"c8a9af4186caee4e", x"5779cb43ff85e26d", x"198bd48a277cfbfe", x"d3cee6679f1d7fcc", x"a4fe50efe83bf5ba");
            when 29993620 => data <= (x"f410612af0bb9c89", x"28489af589f0cbb2", x"f85b7a2cce3ead80", x"80f471397e208dd4", x"9b3c22564232ab56", x"00484aeff7e1cffd", x"9198af0bd1879f28", x"51f17567e58ea0d3");
            when 33659458 => data <= (x"7f0e69f34f569f60", x"3d79209779b5b5d7", x"bec591527408086e", x"2421ad015c5ef32e", x"859e1dcf4ebcbd3b", x"3629321f97c563b7", x"606fdd8c6f84084a", x"9fc9794a31ea1476");
            when 921916 => data <= (x"67b4df40551ca129", x"ed1f48ea1a14a520", x"46bd8fb670775037", x"35961c1fe83dd11b", x"ce213a9a5e1d21fc", x"a6f059ae1144fbcb", x"1608b29efb81c2a4", x"1bf78ff88074bcc1");
            when 17556619 => data <= (x"1c594588fb93b4ff", x"cf96cd1c206bc093", x"a89bc6be3b2d2e5d", x"f08fabbf9661b837", x"6edf7b5e1a490059", x"1e6aad167edbf67f", x"fa95f730bb6f9b33", x"5c0d98842e430feb");
            when 26393367 => data <= (x"a736c27a50ffa446", x"452502d408de6fec", x"c873afd4e3ad41eb", x"da37269542729884", x"ad3b915732b22d01", x"9712b72c96acc134", x"064eef426603bfdf", x"418734771002f5d9");
            when 17603915 => data <= (x"3b053c6a7d97f424", x"27ae66fbfdcf4064", x"e5e6f140e33684d3", x"77994313696a428b", x"2ea0cec99334858b", x"70f3767302bd1074", x"e42fad5db18f21d2", x"ec1c26f455cbaed3");
            when 3499689 => data <= (x"28244ac2f02e3ce8", x"a844d2d3f585ac6d", x"a17ad7085db58244", x"d10ae1b9054da451", x"8c419e5e72531625", x"4d50d35406ccf9f2", x"5157e068062d590c", x"6447aafa8f41d101");
            when 14245342 => data <= (x"f54fc3ead8ef0981", x"e98f8001775c934a", x"30b91e8f4958e236", x"b139a38d8d2bc564", x"ee51c312299ff8c6", x"dd147704ae99547e", x"25cfb6d52f43649c", x"59997f46331b1349");
            when 9234649 => data <= (x"2426552246ee0800", x"ad14c7b23b29fa25", x"6db03095c2621db8", x"2361dbad92c35192", x"ba90494355a1b17b", x"d4d97942fd016c8b", x"ae253d632baa1b00", x"f0078104d30f2157");
            when 27842156 => data <= (x"7775184ec470b371", x"a95711804e3c7692", x"b73b137c4c52a885", x"e077515d88c6f908", x"e718ad6b6c9554ed", x"7ae4eafb9131032b", x"6ddf88214c863af1", x"e0ca59d23fedfaaf");
            when 10103854 => data <= (x"bc04fc670118601b", x"67a2f154f9f2737f", x"ae92ded6e0d44220", x"a66faf5eb5f41293", x"0bf35a1b8c0189e7", x"f5214cdb22142b9e", x"2c2110be67bae87e", x"5b91131747a92e67");
            when 28278640 => data <= (x"113ce3f13952d42e", x"b7588eb9323cb934", x"50ba543064491fc0", x"b9e95eaa29d3547a", x"bd685448b9dcb713", x"4fdd8a958c1ea2e3", x"d87e5210f6bd9f3e", x"60e7e62833786b35");
            when 20573034 => data <= (x"62b69221315879e8", x"96e3dc2f5678891f", x"4d21ca87201f2e2d", x"2fbd2f841eb10ef5", x"04ffadec0c75f8a4", x"c48b742a6b34b111", x"3e4e11d51f2adbf2", x"33dcdbf35cb17c00");
            when 19986903 => data <= (x"bbcbefc61a754efd", x"0148839e6f5bf341", x"4e05bf1fa37d3e80", x"f05d73dd344dad7d", x"7b3461d6762375b9", x"23d26181c8bc3ea2", x"f1e52ae2a674bf00", x"308ea7a4a3b8c124");
            when 1441313 => data <= (x"b66c4dbb2067f232", x"52d00861d43a0edc", x"30f64be5a7c72a45", x"7bc5c0d1d94d87d4", x"3afd47d284763743", x"10ea25b57318057d", x"1cf894a72083ca09", x"c7739f90fdb64eea");
            when 25046919 => data <= (x"cb7f4dca106258ae", x"527591ebe3bd859a", x"8eb5346187edd1f2", x"c79504af8a28178b", x"01c08ae6a3b8ecfb", x"113861b1ed6fe97a", x"cd8938ccfb79d9bf", x"85552daf048aa833");
            when 21209330 => data <= (x"d40026492047b44f", x"e282ec6fb88e3450", x"1bd02d5b8149c4f0", x"cb0072d4a8a9c31e", x"66e4ab9b3fe73d09", x"f7e6aba691104c0f", x"76a1e533dc17d8fe", x"275371bb3be4e93b");
            when 8328084 => data <= (x"850a1397c0d078ff", x"e3e1e52cf2c8f785", x"8827d7c01fd58b4a", x"79158a9619f4cac2", x"335d7d88472d70ee", x"0cfc820d1ab0aeb1", x"70ec8444f0afabb4", x"042133cbb77ede9d");
            when 26774301 => data <= (x"15166c7b5578bced", x"6ba837e3d225f443", x"8fb46434f00be72f", x"8525afef5aa220d4", x"c714ab0696669286", x"4d2dbeb911ad4c55", x"914c4046139d42ef", x"17a3d3d4d1a326e1");
            when 31473590 => data <= (x"7ba3f07e17ce93af", x"dd52d288a3883530", x"4089570a5c4a8359", x"e1e8bfe19788e0a9", x"059326d6b1628189", x"0eea140e4938c784", x"aec16fdf844b014b", x"910bf506ae0869a2");
            when 8079399 => data <= (x"4ff5ca416117f203", x"cdfd1b76ae4472c5", x"f6c0cd2a8cef7493", x"c9a7e8b38d7179ba", x"e9c63923549a9922", x"926866de3000543c", x"7587332a49b388f9", x"f3b3c45f6a7189ca");
            when 2703112 => data <= (x"3a2fd5291014d45f", x"006a4c3a3d03870c", x"9a8221dde26b2a5d", x"35061b357ae2b6fe", x"2e986130a25d09e9", x"7bf867a513b8b03b", x"781cb35055c6a68b", x"8e0a6788e6c78fec");
            when 22540406 => data <= (x"9abb52b87145a2ff", x"c006c88ae1f040a5", x"e51901f18cd6b86c", x"4a9ccf5f2b47c709", x"fd40bee0b12a92a9", x"60cf7231a2d0d215", x"53e4ea5645df4cb1", x"b5cf2c5ffea8e3c3");
            when 31573804 => data <= (x"8161d59cb883a05c", x"8d6ef90e03d94157", x"9423f0dae5061ea1", x"1a8e8b8ed945f782", x"9786ea6271707589", x"6b7774f2dc0c77be", x"78bc2420eecd144c", x"727830e51196c1d1");
            when 28143926 => data <= (x"b0d054e3edb39071", x"0edb6ecd79bbcd67", x"2253dcb99769e480", x"0478e86a21da8869", x"1b6dadfe644a5530", x"572516dc9ea454ef", x"64cec0dab9a579a4", x"c99ad99e91cac2cd");
            when 24716447 => data <= (x"12d882caa6f16180", x"5ae3681f48abfd5f", x"69907874f98c16c3", x"6dac5f3b01cfc26b", x"8a3d596bb4aa6685", x"55b33627114fa646", x"1262993908c34566", x"c36db7a1e0eb4c24");
            when 33872887 => data <= (x"dc79da19ff6e5e8d", x"74d46bd23ad63d60", x"ba268b06be71733b", x"29f859dbe1cacfbf", x"6b9ad1ba1863b074", x"6b6ec1476bc3dc9b", x"177916aa61372eb2", x"2dbcd216f7b1b720");
            when 32792207 => data <= (x"df0b51f6a264520a", x"bc71417b867153e6", x"59a6b9b7dd1f2017", x"a69466d6fdb9a73a", x"3359b9fe26fa5985", x"61a536e0c6a947ec", x"c34e356b6528ae0a", x"5c8c79eb580f4ccc");
            when 17656642 => data <= (x"f8aa347ced98ac78", x"ea1df3bfbf9dff67", x"7bd118c8a54ee2ff", x"2e254f32c64f4487", x"cbbee1c2b8a0744a", x"26e74e8b7b812282", x"a2b97bd0de9cec19", x"469711897d1a8fa2");
            when 8413107 => data <= (x"c9f5d515d5f9bf11", x"dbc8fa4cb8afcdb4", x"07920e984bc3ddbb", x"65bde174d58221fe", x"0a4a22700b80241b", x"468c8f56f341c102", x"0bcfdac26288352d", x"d5f06b5bb8217903");
            when 1087460 => data <= (x"991d9747a0c1373f", x"fd47a041808cade5", x"de8d1ab807640cc6", x"dca26ce8042791d0", x"035ba32b20475a52", x"db958430fa05e896", x"014354f4b09a8959", x"10e4cfbd3284c72e");
            when 3114369 => data <= (x"6488142494b7aee7", x"c0d3b637179cd1e7", x"6cb6057a16a9e04c", x"9646f2d181c765ab", x"34781400746b2fd5", x"8735198268f921bb", x"2bb4f43bf945e6ca", x"b7dc1342995589ac");
            when 6596120 => data <= (x"e8ebbd23773dd1cd", x"fff18a80fa66adf3", x"b6f7557c915ed4a4", x"746bdb0de36d5bd9", x"149eb08cdebe0b03", x"aa6939231666a60c", x"f94f232031b72099", x"90cdde88ed14fa7d");
            when 23919230 => data <= (x"b95a021a78ffcc5b", x"8ff4f2409710ad7d", x"c1e84a257bab8308", x"ca5f4283359306b2", x"f9dc505f90773476", x"6ec777b8e52828e9", x"ae40a316a9f87c61", x"5b1cac3f8e0ce2d7");
            when 9965628 => data <= (x"a4ac248a6149e1af", x"404dc8639094aa7c", x"3049006b2d9828d2", x"6d383549f3f4fd99", x"7cbe85127edc1ba5", x"97e4a09413d5eb1c", x"60efa3630004b8d5", x"0cb53a2deacbabe7");
            when 9865151 => data <= (x"73593849feb0ce2f", x"452b9c6646bc0126", x"9949f7330111a2c9", x"310c87f1ace3f0b2", x"85b61a7d60123ca0", x"72e340eb29d1490f", x"411d1242f91f5a20", x"dd592b3c6c3db70a");
            when 22970091 => data <= (x"e9f69084933783c4", x"1ec5cc8f026f7114", x"7658c68ebd224a78", x"bff059c96187500f", x"a38df0ac5674c5fb", x"c813fce64d33802a", x"1b10f3341457c156", x"7b57c4f0c074c555");
            when 17403716 => data <= (x"1b9e990258a5e2e6", x"27ed21080cef202b", x"0105a2b362f36cc7", x"dbbc6696643161fa", x"8769c9847e096df6", x"c9b281b9a210e700", x"1f77ba3772920397", x"ab4f073832aabc76");
            when 22215139 => data <= (x"c71a73c0345ea5f4", x"7797d9d1621493e6", x"1c21d4adddc9610c", x"0d3834f54cc4f314", x"7f97e8a35e2ef6ec", x"671fe3a7048ae684", x"8275420135fea5ee", x"e2d2c69c1b4ba21a");
            when 13667950 => data <= (x"f20ea9bf1f77fbb7", x"0a338baf4d2374a6", x"750b6cb967c3a02d", x"a60d01be6dfc6063", x"9ac28f38e044a257", x"c1160baf1b9bba4d", x"923c9b6355008660", x"48d4c7d802b7fb8f");
            when 17121476 => data <= (x"28740cce3aba5180", x"74a843bb68e6b685", x"6b0af20319de7b26", x"c70ff940852175cf", x"5e5cfa6a5883ff2a", x"93fe052fb517fbd7", x"02f4949773cb1947", x"83f5f97d2dc8d88c");
            when 23965237 => data <= (x"6ccdcbf0bc631c7d", x"a756bb42d80785a8", x"dce5a675ff1db224", x"6f5ba5a63a9db73b", x"e306505c17ba6c62", x"93f8281f6bfe9504", x"d7d32387f0a7e3df", x"2105042ccbd1067b");
            when 1778691 => data <= (x"1c282f9c62376676", x"396ccf181e3ee051", x"e0ccdba853be81a6", x"282dd38c585d61a8", x"cc98d8b3a426d13d", x"1bff5e4db7eecc66", x"b6e37660f8911841", x"b5292bed0dbc49f3");
            when 22862409 => data <= (x"4879523a869411e1", x"a6a134b98ba1fd6a", x"563e040d86bfe315", x"30b0fc66a73f379f", x"229d6bf0fa1fbf75", x"a359f15a9567163a", x"550bf8f6bb032763", x"0a32e027ce1cf896");
            when 22370155 => data <= (x"02742e4bb6412b05", x"8dcec853b4d97dd8", x"90cd1fa13b3d527b", x"03a61fedb95399e7", x"b609b0804c024d0c", x"d3abe3463034107d", x"d7fc3c6385cecf5e", x"4f39c94504907dfe");
            when 30577545 => data <= (x"22927fc7ec0610e0", x"5aa8b7b28bed32b1", x"584385ea99b4874e", x"13ff18c54edf17d7", x"7a32f84d1fd2f8a4", x"665416a93aaf7e54", x"bb516b5945b079ed", x"f7bcc74f3e19d43c");
            when 9233335 => data <= (x"dd7c1a6ff518bd7b", x"f04b593020ec5a41", x"a71d1b319f140f5f", x"096e410d078696a6", x"98f44f215bd114c1", x"79e413b36115c90d", x"6794cf39e23d80f0", x"2d101e5f9684641c");
            when 21311820 => data <= (x"09734c9d7ef455f5", x"32a1c4f4df79b738", x"e33685a5b232593c", x"883cd39ba46048dc", x"f3cdbf83445ac2a9", x"e43d955e6ab7aa3e", x"4052380e282c0b67", x"904ed26e67a35e78");
            when 14802218 => data <= (x"d188c17630b08708", x"38850a4e0b0a2c7b", x"a28de2f149d571f5", x"cd9a712ea3ff7f4a", x"1a0c255975656df5", x"d65a2672bda181e5", x"7dcdc1aeaf85ca4c", x"62cd8cf432ab61bc");
            when 16967564 => data <= (x"4d0659abd9ece754", x"4cc6e5aaa8928533", x"34e52a5ff7264853", x"c4143374fe96d9cf", x"e0abed33e7f5a1cc", x"b75b47ecb863bdbf", x"8e1f19112de78ab9", x"bed6d304e445a99c");
            when 14570070 => data <= (x"681108df1bddcedf", x"dce40af98b41485c", x"e11651554ca2a0ad", x"d9c92224b09f4bc7", x"300737438f6b968f", x"58711b82caac3b09", x"87e49c0372c6ff4f", x"d6a3073764964aa7");
            when 20398263 => data <= (x"2370d00a0417c70e", x"6428b9596b167097", x"73960b5f1cbd5243", x"3d5035e4fb4e4a8e", x"dcf6089753543fdb", x"8a47008cd5dd2614", x"e7a903b6298d0efd", x"33f80faedc30f39b");
            when 1053268 => data <= (x"0e0015726429c6f5", x"5314cdb674678917", x"2bc2250b529ded6e", x"e8b4d566b1b7b394", x"66d658515f2b0d9a", x"c85dbbe7b054b5f2", x"9329b9bc353e7f7c", x"3c8f11df34e0a625");
            when 22422796 => data <= (x"84212da33cbea524", x"4804a1ad663bc6de", x"0e8e0d60f7f3a5a5", x"b671760a56e1ddc0", x"4cafd1637340bbe9", x"7d15388b89e787c2", x"f2b1aa0c17f65364", x"c08974ef131af448");
            when 32113332 => data <= (x"9b0544381b454d33", x"c0035e38eb2b6aa4", x"512e00d5901f90d1", x"7ac8185ebf327cb5", x"29146b27a00d3d9e", x"e476ff29e9af5087", x"c1e5c0109720c8c5", x"22c32d8b01506941");
            when 23019458 => data <= (x"240725103ac16efe", x"55f7c06234cc5fb3", x"800f09360bb91f69", x"78831d2668d2f417", x"824b5a63906b2d7a", x"369f4984aead235e", x"7420e3e65ce4a718", x"8df74e1f34758af8");
            when 26696900 => data <= (x"60fb91448eb6fb0c", x"62d99f936389b9e9", x"26bb169a42416719", x"b7040578dec415b1", x"e15018d42356d77e", x"95837e3b8df94c4d", x"40d29d6d00083f33", x"8b92bd01417a933b");
            when 10497163 => data <= (x"794cdeba52f5c4f2", x"05edd5a941d5c836", x"5b8f9efa1b1ecfe2", x"8a15d2cb08eafbc2", x"45b6f74d8bc0ffd0", x"00886d1960c93a2b", x"29f46aa8a738ab9d", x"bfd10afde747e093");
            when 451296 => data <= (x"d6e77507f573609c", x"38179fa4c2ec102d", x"196312bb7530e2c1", x"afa5d2862a330444", x"20633c407cb96265", x"4d0ca54bf46617ca", x"684777dbd250da4e", x"e740521029be8997");
            when 28054670 => data <= (x"e88c20d83c2c146e", x"b09c6de03ee802df", x"35fd396e8eded876", x"a4489a16d9984fd2", x"711cac21b1a805ab", x"ca108751a28fc618", x"b32008b1bb220986", x"078afd4b906ee95d");
            when 20376750 => data <= (x"f893c4e6c9dbdc2e", x"2bff144532f32d56", x"5bf1ebf224665959", x"cf439b5a7d73574a", x"8f90d6bf8e116fb8", x"1922755ebe18224d", x"58936b49520e3847", x"aa79c1c61db410de");
            when 26481720 => data <= (x"b59bfd13edf3c1e1", x"1989b2d9b6810dab", x"ee80906725ae7581", x"317532424dbba12d", x"93a67d77b7883799", x"1b2005c5a907ee64", x"ee62415635b1a930", x"fceed680c5a6bee1");
            when 30383288 => data <= (x"cf6317978e07996f", x"1858724b8de45e71", x"bacd14ed46ea5904", x"6634d90a720439a8", x"a6bf1a113a880b4a", x"afe6a9b23d6d08ef", x"3e5459987948bf11", x"c61a2bfd078226e5");
            when 19641814 => data <= (x"c196bcd41327f671", x"f9149b24a387068e", x"5d05bdac6b42f581", x"9e87720b4803bf78", x"a1ba00ab92f17b5d", x"e9c53203bbbf7553", x"331a4383098fe959", x"7fb4554f6bc929be");
            when 14054139 => data <= (x"de2970e80cc4520c", x"08c3588c7a4e0773", x"db74f7451073487b", x"4e670ef8ab6b0590", x"f8ca5a691d4242bc", x"a34fec343fdb144d", x"6e28ea485cb96921", x"971301774535d919");
            when 19926300 => data <= (x"b34f59b94fdbf79a", x"88f2b0128d5f3884", x"3a5b511690130db9", x"85972552d79568ea", x"baa97133e3f5a525", x"894bcbda7fb64a33", x"cccf3066a905bd46", x"0b3b44bcf9bf73af");
            when 26009366 => data <= (x"299e6e43026e8de6", x"2da028d10cb37628", x"212db6572be3f9b6", x"d676138f2c2147d0", x"bb724166d291a542", x"26d3895962846853", x"ca0c3b52ca2dd0bc", x"2f0d0607a47fbd7b");
            when 12615906 => data <= (x"3d8f420e2908c7b8", x"0c2efd852f66f367", x"c3977fea748442d9", x"46c57e68e5f9ca7e", x"215560bdc02c6cd3", x"095755188acad215", x"0433ea845c2e39fe", x"3b5af17f7e0295c3");
            when 27894284 => data <= (x"00a3e93eb710e357", x"8a35c23c13e8f130", x"82f0e342eab9ab79", x"b46afae80aa1c1ab", x"586a24fe61cdeeeb", x"f8bbd3473ad05419", x"a49ab897ff3c8b28", x"1f256810fa91a524");
            when 29424588 => data <= (x"c521f0c28fb8d9a9", x"744453b70527249e", x"b9b83b22bde6810c", x"02ca49d995dea3b2", x"ec0e66d044caf634", x"d093765bc737fb60", x"b2a49de7aa3f278b", x"3123e7899b629482");
            when 13940274 => data <= (x"70ba8a9a82b73fbd", x"d3f30d499ab69172", x"0be16376b9108666", x"76b3079f98b016ca", x"66460a1a8b16b5fb", x"edd058c426ef7f99", x"bafbdb20789c81cb", x"999527f8f9f099a5");
            when 24172763 => data <= (x"4dc659c1d6fb90f3", x"39be522a0ec183a4", x"7c678fefda3b3fe4", x"99ac67cee7471737", x"82f9f76ae5a278e7", x"0a88c78ce2d86fc4", x"d43a4f0cc05199ca", x"c5889793807f66f7");
            when 3336498 => data <= (x"c64ae4de63efc473", x"587ce9038f8d8700", x"8f2a201f3a20c8de", x"a1efb13a528280c9", x"31962f900d537926", x"65eb6741b975b6ef", x"0b497cd9850e2733", x"ca119e219f95b0c6");
            when 8983648 => data <= (x"ff54bc26fabc6e7e", x"51192889b4b01cb9", x"99d0fdbb25a4fe58", x"c9f44625448a099f", x"a8b99e46d0000c55", x"d28acca52ae77230", x"6780b27e2117dd78", x"e1d2581d07a0c083");
            when 29780487 => data <= (x"474907bd47b01c0d", x"a9532db3cc3a82c3", x"3ca9f482b86f3ddd", x"ae285c750dcbeea8", x"77d960729701007a", x"d6c6311990f01228", x"42e75661f040c225", x"539eb650c5b1e03b");
            when 23769849 => data <= (x"465f3f64ba1c8570", x"dfd76e878cc0b906", x"4dfac84dc3234fbf", x"fc91ed3441015508", x"aa2e98307e645ba8", x"a0205a4802710776", x"c57e0b67a2793f57", x"c2978ae7d1be5569");
            when 1910567 => data <= (x"0ad5408f5e7e9a91", x"3b6dadaa3bc116b3", x"a30cfa8756392a76", x"9decd50e95e8105e", x"5a1abb4e462d00dc", x"b2b519883df665cb", x"04ce06b62e77ef5c", x"8d6d5d2050e4ab62");
            when 3450217 => data <= (x"99c952ad590861d0", x"356d4115fee544d5", x"3b216275b3cf5129", x"a1a31e239fa19cbf", x"4c21d6fe565bdc89", x"054a1d8f3d41f052", x"e450d50cdfe3df4d", x"6564055f459a8fbf");
            when 7037448 => data <= (x"f3342fe0f7bc66e0", x"4a9dccd2d1097c17", x"320b4c1d1a867526", x"065bf7f9f7fd5f9e", x"a365bd1c4b5a20d5", x"cd19a0ad37f5ac69", x"0613827936cb9bc7", x"cf99300f60a2c8e5");
            when 22444529 => data <= (x"d9f0ada54b3c06bc", x"9e9f38b84374a291", x"aac04c7f0f61099e", x"493824c6d46d4c9a", x"3397a4df1ba09e4f", x"6c4549259db41fcf", x"c1713b71c692f770", x"2cfac5e34276e8f2");
            when 18772286 => data <= (x"b6ee1268db91218c", x"8f55d4cc9c50f767", x"95067e855571a3b1", x"be774323c9443068", x"e9834303b692faf0", x"5f89d0d603e73c6d", x"3d33c76fab82d83a", x"e887abe3ff5bbe85");
            when 15887325 => data <= (x"cd6f186849389f0d", x"e94b6744eca8155c", x"b167d4a992aae1c7", x"93dd96ffab3b1bc6", x"ddc5ed8bbc841a43", x"295c4e3f8c89a7d8", x"e3321cc050c9cbf8", x"f735c4ce35da5fe2");
            when 23273676 => data <= (x"b2be218af61da87b", x"7b5f3ccfd063f910", x"9b0ece95f2854752", x"08237537ada4530a", x"a22be591ebb9dd23", x"f463023b54b4346b", x"5b4b058d5a4187b9", x"e92832dbb38f2125");
            when 16141951 => data <= (x"285449b0dcaf98f2", x"838464713e762ef0", x"366a777690f1c574", x"1819005ff6dac1bb", x"b8eb4af2ecfc074a", x"37cc50ff54cfb024", x"f5df9298f277624b", x"dbce0c98f8bdf9f1");
            when 28999832 => data <= (x"dad7a52f27c89d2d", x"f61c3b8359f2dbcc", x"68b08ef5733b55a7", x"f09cc237cea45a0c", x"55b6e2a3d5440549", x"116dcdc41f4846b1", x"775957407ad631ae", x"7b51f2bbb38f6bd6");
            when 12235628 => data <= (x"ae542a66026632a5", x"fc447575fd22edd8", x"ca573210e26bbcf6", x"d05ce4a699ac1add", x"9d80cca66a391755", x"36b7e9fe600c60c8", x"21eb3e4d376dc409", x"b8109800d363db0c");
            when 2115023 => data <= (x"73057e1cd7fec972", x"b3ea365351645462", x"06b35278642f821b", x"3f5c87c88f0da2c6", x"eb32f68b286ee878", x"30351bb478271069", x"f819270ebea734da", x"f340ed79f226c2f4");
            when 23274169 => data <= (x"3ecd4e7b56b6ab3a", x"c44d9c7847ea7d38", x"f0c604a73999cd1e", x"1fe2fac9a4f1d803", x"e3c9d0ba2b1bb014", x"bce95c1d5ee8a6f9", x"64a7b8625c73c934", x"891eff676bf41d60");
            when 27126540 => data <= (x"e9a56d361b934aa0", x"491b66c5874a428c", x"b23552ad202acd29", x"5c25b5133065190e", x"c90daf3d8ff613dc", x"d0de88fb546b9154", x"02fa044f4d2c4d61", x"9be537021ed0105f");
            when 30096050 => data <= (x"258a0240211e51fb", x"cc3dc3eca7cb0557", x"772ad1b9d3c90201", x"4869125a79a365ec", x"48d23fd1de4035b7", x"ffd2295045cde5f6", x"e9ecb86716507543", x"0c6c97fe5e474e2e");
            when 11639918 => data <= (x"84b61efcaa690a37", x"206663d1fc12dba6", x"bf0da81fa8c45ea9", x"4fa13c718517dc48", x"77c81d0a54796d7e", x"e9e0fbd2f9b0e661", x"59cb7ce16d6ad79a", x"176dd403a6db8bd2");
            when 25474762 => data <= (x"3d16031ee09dc303", x"94796407b09609b6", x"0ab8c8bacc6e06b5", x"71d2952f77fe04f7", x"f67aceba899fc578", x"d556d282c6798934", x"19e7d7786cb0c4cf", x"7aca40052f3097c6");
            when 22530936 => data <= (x"fb1113189b5c3af2", x"20d22f45dbdcaca9", x"59b68686790418ef", x"6c68d6110b2425f2", x"de58c11ede592c7a", x"e18b82fcece6cf0d", x"ec6465659403d3ed", x"309ad20b6bc8d4f9");
            when 24996707 => data <= (x"d7b1d0d9495cb5a1", x"46a0a3291a8edd72", x"51a6af980dd2d906", x"06f74a2fa6eb16a8", x"94b6c45489d70100", x"352b0cc65e212f39", x"61f5f55dcad7b55f", x"46bb571bcea866f3");
            when 20693218 => data <= (x"327223689f895b52", x"c51b282e883ff77a", x"fad22d64518bfd88", x"ff50b55ff547e763", x"679a8139a21215ee", x"71428de4bf4eae65", x"abc56785fe5aabc8", x"ee20cce206bd2ae1");
            when 13107094 => data <= (x"fc389bc81999ad9f", x"e189253767be01f9", x"becad4d69222f153", x"cecdb9e92102d9dc", x"b709b0fd8d5e0a2a", x"a6549d7bc3b580ba", x"e30a5500e54ead49", x"53576bbaf482bb9e");
            when 24140522 => data <= (x"8edfdcd364218eb3", x"f67e9c6aef161527", x"895d9d84c5666475", x"7d7d14cbe0d16a8f", x"a82fd139fcc7345a", x"ab52842dae1df2ae", x"c2eb250fb6b41fa6", x"a9c56cbda8fa9c0c");
            when 28372358 => data <= (x"c8c7fb52eecd4119", x"7ed4d53f86922ac2", x"09c39b958cce5275", x"1649677ec7422ab0", x"e6f84e9d1bc8eddc", x"d842414957ad2739", x"2a68a33418c62e0f", x"1314a1d001e485f6");
            when 10537678 => data <= (x"bd12a235eb74435d", x"5c969edab04022e2", x"3c1c85af398030d6", x"ed63a2a07a6eb9c6", x"5c04cd3159d8b7e6", x"1969b9dac0f61986", x"22bf198472976093", x"0fb2d56c04d8ea3a");
            when 28990677 => data <= (x"5c362efc18ea5d3d", x"419a87978730afde", x"ef4cdd0e3b992f83", x"f93679aa967e7735", x"52cfc497438f3697", x"6c0c28646a5ef87c", x"678db62aa7307b5a", x"68889ee3eef8f642");
            when 12270960 => data <= (x"96cf2908d5aabe33", x"947ee95fe4f028b7", x"f20657e83af61978", x"a83976fd00a1630e", x"06a655cbda1ff35a", x"95bb6c8af98e00a3", x"e72ffb9eeef8e415", x"eba583c8ae5c0d0f");
            when 19002324 => data <= (x"433fa8b6ae570145", x"1512928cb8f995aa", x"a7d570edd8d5b0a2", x"61881cd64ac1e41a", x"b76f742bf6204bb8", x"aec7836d068f6058", x"3600a38203c5dd81", x"21b3f5266a4e44ef");
            when 18267766 => data <= (x"7366f6a338f53fd5", x"86d9c1c566550bed", x"8ee1de62b6026981", x"2a04fce627483849", x"d26cd98df3a0d43e", x"32ce5c21b0b91aad", x"55f54c1cc7f45b2a", x"f7fe5cfb5ecaa4ac");
            when 28932782 => data <= (x"143f2d83260aa5fb", x"2cfc5aa44dbe116e", x"4a8d235c77f3b8c5", x"cbab693af69037cc", x"73c876e1b76d4bef", x"0149736901bd137e", x"8b970cca2b0819f1", x"001255a070addd85");
            when 22047612 => data <= (x"6c15b284476e2f0b", x"2399b9d0da719297", x"06b61d9e97a97c5c", x"bb59d0897674a75b", x"12b21caee2136a48", x"b6fb1144f415105d", x"ed4e98dc9794e854", x"86473480c57c7639");
            when 22412494 => data <= (x"b0c947afbd513d09", x"7dbae08788f6fbc5", x"e0df47b2cb9db6ae", x"ac06c9a55ed5bd7a", x"77facfd46b98ecde", x"2b4837b04eaf8e5f", x"cf8fd45c2d626884", x"4d58843561ca0d58");
            when 6326992 => data <= (x"c6a1dd203140339d", x"835d73da1b42c1ec", x"cdc1b2e10cc3c19b", x"40b6b4eac93c9cae", x"a60442b6cf9fd01d", x"35d3a63f2aee3668", x"5fcf55ba7acccc00", x"4ccf70e99135cb7a");
            when 7499585 => data <= (x"dab11e23e9257bb2", x"88f895c721d544e8", x"eec6409b79504d47", x"e385cd826b2b73ac", x"401d5a49a0b2a04a", x"81e45ee48a9b3c6e", x"7437c616a0ea604c", x"5c66dc14fe37cbbc");
            when 13772006 => data <= (x"50a6bf0b0b7a7d00", x"9d1ece804c13fd82", x"aa0175c38712024c", x"82a2bf932224eb90", x"2ef4dd196229994a", x"15c1a3f7d0e3c930", x"670d8d3533a0d81b", x"6e7397565ef5304d");
            when 10701234 => data <= (x"92f50692043a8342", x"04e74d8381b25d4f", x"d04c2cb582a7b157", x"5b85cd71f74f5d92", x"caa681f6ea890edb", x"1da7a8b16cf6ea36", x"8e43d4ad9e13a547", x"3a0168f02728e7c2");
            when 467605 => data <= (x"7779856933e42124", x"f2e5ce9930b0b59c", x"f0f1441c29b2aec2", x"eebeb672f4dfcdfc", x"7dc6cff9f8372e11", x"c342cc226ffc31f2", x"9681e0c3bf72ba4c", x"975add5f1d907dc8");
            when 3652438 => data <= (x"f16cf876f490a762", x"4b8ead708229215c", x"b0fdd4acd22eacca", x"134199502714f953", x"3fb68aa7d8feebe6", x"4c83f3331dbe246e", x"c75f35225dfb977e", x"bac8ffb9ff24027f");
            when 3721956 => data <= (x"763b1b9e7e25e18d", x"53c39136bcf3826c", x"bc65f60ca169e7bd", x"0e87e4f849889df9", x"004bc7b09ace13de", x"473ac69f1ec01f9b", x"0bff05481c75e518", x"f6f5fe33b536c594");
            when 8986308 => data <= (x"37402866ba3f8a7d", x"01ed7430b24d5114", x"998df50308e69f50", x"2a53db7a8453c0f8", x"5b6c1e29a4a5bed8", x"916251803b9de66d", x"0d407f6b91337441", x"94aeddb97dfd5d89");
            when 1633793 => data <= (x"f1496d97253db65b", x"7d384322d5aef042", x"91f2b5d94cc20eaf", x"1ebf39e895cf936a", x"04d1735a47d4121f", x"551371c590d1c256", x"7233ec03da9e4ea8", x"d7bf10ff795990cc");
            when 21078227 => data <= (x"42fe4a346db139b2", x"acc7a77f36cfe74e", x"d0acbcf3a2cb5a0f", x"039462c68262ef96", x"31e7815ff1e4a576", x"b58ce81792eeac85", x"9704253ed367dae5", x"5d12aaa937bd547f");
            when 29354883 => data <= (x"b36a5ae57f1e5e08", x"9c27289ccdfe599c", x"51a7f8a882c118eb", x"65344a087779df65", x"64a25e265238848b", x"20f0bc61f59055a8", x"9355707f01454584", x"a22a3487e5ad207a");
            when 20742321 => data <= (x"157c94939010599c", x"4fb53162f8046ecd", x"23ce9c46eaa0a7a8", x"e6a7b2f7f54a76c6", x"238fec6f5e3db858", x"7eb417e95c38a3b9", x"4ec8ba6ff0494b63", x"2c22ffdd2d8e48ed");
            when 24608154 => data <= (x"1d970b7db25b112d", x"a25b51a2d66af863", x"1c00b1413d9bf365", x"0ea6df7b2fe32ca4", x"542801c9cbe6c461", x"0c4b80c1de88ddab", x"e83bfaa9efcc8aba", x"c76442facd788657");
            when 6686733 => data <= (x"b2564958d0754f13", x"18e876e9bf66416e", x"c9194b7aac37996b", x"4ad1a41eb2651c8e", x"ff7293da1ac39bd4", x"3b6d3e52cb4a6e0b", x"ac55b45d85d33367", x"05d210464b203c8b");
            when 5178520 => data <= (x"7ce18e02453c9432", x"fa22a0497f200390", x"9becbbf9aaf5ab92", x"98dcabb0c69db12f", x"ef503f328e65ea1e", x"a6717027ece9690c", x"b867e6027f8e76aa", x"30b2f8b11c672499");
            when 16740621 => data <= (x"13deca74b8a4ecbe", x"1a6710cbcb5247ff", x"0fb08790fa6d2105", x"0131e9f68b8a9177", x"5553591afd364e79", x"d1ec8c84bef62c85", x"e47a4cc9f83459de", x"5aad0b4d573f8d84");
            when 9285875 => data <= (x"ec5f5901c1f9ce18", x"249dca91051a7f32", x"ec6516b73b71c46d", x"54632960d21c54f1", x"1c8a4b4fb34268bd", x"f0c41285891b4f4d", x"b6d31b39dddec15d", x"6d6b8245af47002a");
            when 33918767 => data <= (x"fc779449348a8835", x"6c5702413aeb58f4", x"bc7743f69b9b9b84", x"11d2e35492fce4d3", x"558c27d03dcff561", x"b7192502679e7479", x"9aa629caf9661f8c", x"6f8fbce149da8c34");
            when 20750443 => data <= (x"a32ac19595deee39", x"fa6d828c7a5b0805", x"dacb6f269da4fb03", x"f38f8ec5a937dfef", x"0055f330a2d5b3bb", x"9369df6b8286167f", x"7533a1189acd196a", x"0292c9eb294433bb");
            when 5226143 => data <= (x"e52a7e19f43dfe6c", x"d21f383dac8bf360", x"8493701f00650334", x"672ad749849c1baf", x"eb457e75107ab859", x"0c2885a359ab550c", x"470235d936801791", x"39e816b7e9ca1613");
            when 30885798 => data <= (x"b9ba101bfdb6ecb5", x"e8f4435a04855b44", x"4341f084f20d4c06", x"d826d5c1396fb681", x"f7e3acb94ac04612", x"aef48f5a9fd8b3d4", x"e684914a9426861f", x"fec5519bc28ccf91");
            when 6506026 => data <= (x"1cee002caeb7a1fe", x"19f6d86a9629c52a", x"edf5a62932ee098c", x"3b1e36b3cbcfb5a8", x"b6e112de9a236c52", x"4f5368595d67c228", x"78dd5e26d793ae92", x"3465c5973f8a5439");
            when 8243701 => data <= (x"07753a8ba3546baf", x"970149fc9704abc0", x"6ce78ac12711eeca", x"713e0dfec931b723", x"cc0cfaf86f7bb698", x"94bf7346eb23a92e", x"39b3c1fff71a71b5", x"55993e566460c4b7");
            when 22182781 => data <= (x"b992d247424f0bf1", x"582007a6a4460d99", x"2e6fcdb4fdaac8ca", x"c508fb01ed5a719d", x"23a7b5fc96bc93a4", x"4b4c56ab3e02ea83", x"7f9534f571c6ad45", x"5e3fc39b52a31267");
            when 23321267 => data <= (x"6e19a00f60d8474e", x"e0818a403120db60", x"637e53b5a218b84a", x"9317b36bf80b7a22", x"d36190ef46cc5883", x"59249fd09b615cba", x"3a641e8d348c314e", x"a0565e931bb9a24e");
            when 29764568 => data <= (x"cb1db8d920553800", x"4917ff6d7ec336ef", x"2fb4cf9aba9682e8", x"57eb388dcedbb3d5", x"6c0560988170f2b6", x"7d51d410d44b8250", x"b6582a7d90174208", x"7507da1154db4a3b");
            when 12970822 => data <= (x"d9d919fcf70712fb", x"1950c5ded67d769d", x"fd173f2d0a03dc2a", x"efee7c913980180d", x"a97a1f37443717f9", x"32cc8d995c350a9b", x"69d25a7e95e58971", x"ac507c13dc7f8d47");
            when 20771445 => data <= (x"61c76ad2cb65b519", x"572b09aac62ef59f", x"01302485bcad043c", x"9eb0992c53e7605b", x"20e9cb6736a43cbb", x"b33c826b922f06e0", x"a16a0db0c67769af", x"3fda1616db2e2f63");
            when 17561376 => data <= (x"f51522468f4c7a10", x"e90f27faec7f8168", x"c0bc0c44f4ffdaac", x"14629d93c8cccc8a", x"dcb8b384c290f111", x"58e998bcc76d0744", x"d537fce0c7c5814f", x"210a7cbb917576a7");
            when 24656685 => data <= (x"592211b7ee87a05d", x"b768bded1b02c082", x"2131e9298b79ae54", x"3d75ed93372067e1", x"c210fe80f1cb253f", x"e4e10efdacdd5ccb", x"5a5dd8f76afbaf7f", x"f97cf3855b1dfba0");
            when 7215102 => data <= (x"3e8926a9925702dc", x"259f77626f96678f", x"31e6777d101d5fed", x"0044a9e3c2374f7a", x"ca4a5f8f79138759", x"ef9913d43a8c544a", x"8a6a2d7dddc64f0b", x"8dd4cc5545f18e85");
            when 32036870 => data <= (x"7cccb638c08be259", x"eebb4f31b03d99cf", x"07644996ead4542e", x"7db73df72d2194b0", x"1b54c4201924cce0", x"8370f9c289f399f7", x"00e547559a1fc501", x"0af9b28fa29e23cb");
            when 30727640 => data <= (x"569fb42450280bcc", x"85fae5c783b9fd38", x"9f5bb5370217e524", x"fdb84ded65c4b025", x"c9cd775e2b2432de", x"3464ccedfb5af297", x"4282acb80ab5c10b", x"0342fd5126d14fe3");
            when 5839051 => data <= (x"188f78ae00d8efa7", x"ef612429136cf5e3", x"326d89eb83eb1442", x"391448fbdfbf2419", x"aa69fac175e3bedb", x"bd6ba6c3bccf83e0", x"bc2fc681068de1ad", x"6f41cc4122d17a48");
            when 23944715 => data <= (x"62bbf28e57af07be", x"409b71414b0989d4", x"02773f8ba5e4773e", x"67e678b8f01cd21b", x"a881f489465bf7fe", x"77ab730c54fbd87c", x"ed79f0c53f572325", x"394ddfd0f66d562b");
            when 26242448 => data <= (x"f9afd3157e3336d4", x"5f091138f9412165", x"b7e4096293b08bcb", x"90893802b3ec989b", x"fb84a29b06ea1782", x"248d2f943a8417c7", x"ce60b0dad960257d", x"76d8bd758830278c");
            when 28282502 => data <= (x"63d6f3069396e037", x"cde2d7390220cb69", x"1b94815b83f30919", x"a342f2680055dd3c", x"fb26a0d6c2ed897d", x"b816deeb34af42a9", x"9b9c6f1b700a114e", x"87323e111848f368");
            when 28625415 => data <= (x"36b49334424c70b9", x"d50d99934c6ff69c", x"3c63ea716c86a6e2", x"03a9c3f325cbbfcb", x"47b541c4e9a26163", x"cfdbc5d44ffbc683", x"6946ecfcbb3af91d", x"2dc898bb54f2fe5d");
            when 29550439 => data <= (x"c0ba4b599497d06f", x"54b5abdfae96369d", x"6d7442eff0db3d76", x"4d7699ca4f36ffcc", x"7e111c013bc81552", x"78093c3c61ce4902", x"2200024615a398f0", x"26ccc8f649dee04a");
            when 33786172 => data <= (x"105e373d594f672e", x"50298d7bcfa484c5", x"45da1839cbf5dce4", x"99a3b5ec0066d09d", x"53162b3b37189a68", x"f051daff08b03718", x"0fd99d5eb9b77615", x"a0960e585dfc9434");
            when 33340458 => data <= (x"9776583d9d6dc4a6", x"bd3e257481ff00f0", x"a48604a2d5ddf981", x"1fc6311a5b21b2ef", x"c90a3be376b0d10f", x"90fe747920b90c48", x"ced897a7018b8eb4", x"c58d62405bb10728");
            when 1152577 => data <= (x"a95f65882a6dd663", x"8f614e98b5eec466", x"a0f6293f9fdd6954", x"e6ebb396dc269638", x"a34ad751a2a625d2", x"b048d2eee5768a62", x"7d2a300f433ae08d", x"a2ac6b3f3956dfe9");
            when 1414953 => data <= (x"60e3ce2bf1879756", x"b4110577686eaee5", x"e5fa18a9de345100", x"0d47f6186fbc8637", x"84476d8e31cbe316", x"8f4be3ca08eb22c7", x"f82a7fbb80330291", x"dee2bb163b51c4d8");
            when 12751504 => data <= (x"06cfcc2d677562ea", x"065a3d8ab126f802", x"408b81bf4024daab", x"ecdc40726f058ec6", x"bb3adfae3686123a", x"1929e34bfc9d2572", x"e22c5c81133cc3cb", x"ff7b6671f4439ab3");
            when 10412312 => data <= (x"9d69b77acf1e11f8", x"c101626fbd48009b", x"0a22934eeb1c738c", x"7a2ca35efbde6ca3", x"e778780d4c8380b4", x"55749d405565b3e5", x"b2369fe7afda813a", x"29bdbd4bd120eaf1");
            when 9116600 => data <= (x"bff12d950cae38ac", x"551c43409a9e709f", x"3c26196a69ce7381", x"c823d4484374d4fb", x"16a0b8c53688c686", x"46288aa28679d5a4", x"11d2f1b0a67b1848", x"77497f07047531ac");
            when 20759552 => data <= (x"a018d773b666d6c4", x"554d16afaedfd295", x"8599d44ea09c98ed", x"32e2f6994362973e", x"a5cafeb2689983dd", x"a5ac6fa296a4dc55", x"8a776e909d4df78a", x"9902caa9c4c4707d");
            when 730618 => data <= (x"7a98e9f25ad0811a", x"11a8959b554e3a48", x"620b399ad019f9da", x"c187929c40ea0617", x"ae1d0e64bc3b8536", x"67df6827b94d7906", x"0153d1ee2005eb33", x"171d47448b3e65b7");
            when 12199450 => data <= (x"e781822a3da25e2c", x"f0fae68c49ec5c6b", x"8ce677c55661fce7", x"7ef62f37dfd198df", x"a231f3465ba48b1a", x"214d27a7baf0d20f", x"fbdd842f4cd692da", x"258a3465ee95a0f3");
            when 28549695 => data <= (x"0f214e789c4d83ef", x"2f84c9f8b9720652", x"8f712809e6489fe2", x"29f9f3c525d96566", x"9b672956e8d7da9c", x"1a7b29f92fbf20a2", x"843dd691c86eaf74", x"08c16f7d844efb42");
            when 30503980 => data <= (x"00cbffb012250fa0", x"6743d846ae9a6dd8", x"a0530381f0e0e6cd", x"7685ef4719401262", x"3cbd4bae9c72a65c", x"daa78456ccf61ab7", x"754e6b1296ac2c68", x"1d9d27e07ff8caf2");
            when 9316166 => data <= (x"01f180f35e247436", x"e066cd08f3d1d7d0", x"38f72e3e1f72fe9b", x"6d7fa29072e6091a", x"2fb4c4b56ecc8f41", x"998329e19a80e34e", x"0a16a1cae84cb574", x"ab49e51fb0b592df");
            when 24959304 => data <= (x"c40ff24ea5cffa39", x"63f18423ef95fc40", x"3b6fc2e54e44c113", x"0a11a3b5691c4e26", x"d5b9e1da6e367338", x"0c7b5c8bc71763d7", x"522048ddb943f4d8", x"aeef75dc3da0d6d9");
            when 2099797 => data <= (x"23b619f2883bb8bb", x"21c73df1d17cafba", x"2c30ac0f8655ea6f", x"262237e147c3bc07", x"3850fb4b08b8ecb0", x"56e0ea9b9e20a46e", x"b86c59137bc04e73", x"9b5bdf30ab8d9a8a");
            when 16892590 => data <= (x"39e92e638e60cd42", x"51d749d41f6d21e2", x"6a63153a25858b11", x"a58600de8630ab39", x"5764a93acb46ca20", x"9babd1e5d5880e67", x"06e4ae663e773c5c", x"287f543503bac94e");
            when 16518632 => data <= (x"cfcd641ff18a068f", x"4c94d19c9bce8a71", x"f37737347a259cc7", x"21e8878cced4ec14", x"5298e03039a9b1cd", x"040eeab3ade96790", x"5d214fbcf1920bbe", x"bfe81661f19af98c");
            when 25452195 => data <= (x"1143e384ca8052eb", x"e25d784de0f9b8c3", x"234e0bcc7a6a45a5", x"2dc4359dbfa4df97", x"a045b20bee1b5b48", x"2b63e81d67dfccde", x"27d2a063621b9a2e", x"da59f16a8bbf805f");
            when 15064032 => data <= (x"b3a2f13d6a43beeb", x"51896e379ffee96f", x"637812db07f866eb", x"c3da9b02416e69d7", x"aec6a362b2629cfd", x"c688dbcda5f97b5b", x"205c8dc0d92a20cc", x"89763547202b920a");
            when 6991240 => data <= (x"59b51dc83870d051", x"40ff4857f52b4e04", x"5bcc53eadbba5b48", x"7bc2fc42eb32cafc", x"c28cde8ef4dc98ea", x"6d798979990b26e7", x"2cf1a32fab3566ff", x"dbd9d705a9dff0a4");
            when 32595530 => data <= (x"6f32ed3f0e7b5b9d", x"10d11f29c7f8bc5a", x"db3b1ddaff164fdf", x"4ad1ddafbecaeaaf", x"b54f1976be554605", x"af27619482cdbfc4", x"fcaa3131bdc9a572", x"a75d88c9a9b9d0f3");
            when 7961868 => data <= (x"fb63f4dfa71723fb", x"cf669c3068f2d158", x"acc2627442ad930e", x"98f801c399be7341", x"27c00e2a8309487f", x"06c928871d431022", x"8ad5143870a963c1", x"3cdfc35be09e9bfe");
            when 16709748 => data <= (x"fc39dcba2a59ed30", x"14be462554f8273e", x"03fd5c7cd31cf579", x"20480cef75dd2834", x"bf3ef1854b6d89c4", x"aea2ef4545dce3bc", x"6fd3d78ea0755980", x"248339d347c88894");
            when 12333586 => data <= (x"61ce37e4a9c1a13d", x"df0f5335896438b6", x"62ae32d8569c1362", x"5cccaf31b2429154", x"82bdf70f39aec368", x"4a3b0c9041871c4d", x"6a016e0fc355fc44", x"a2c88f4dea73cdbc");
            when 15967746 => data <= (x"f14c4a66bb85133b", x"9ff57066b4f46d4a", x"18bae03c76031c93", x"fbf02515878d4873", x"718a4eedc86e3e37", x"c8ecb936a3d4fef9", x"ab38554f24725148", x"3fc856fd902aadda");
            when 28019849 => data <= (x"711b039c986acdf5", x"01b183696f0c9d86", x"e48ed9455b06c5c8", x"e69da4cee5743c72", x"64b40e90095ddc71", x"63ad8eb394113f9a", x"f838f8870631d957", x"a4a06d0113b3aed9");
            when 25319287 => data <= (x"8453f13faf722f4a", x"60329b5f82177aed", x"b3eac56e0c16669d", x"19a4f8014305ffef", x"95c49a95f917f31a", x"deb47b30e4671d8f", x"a3bb1ca1063f2c39", x"927f79302be2d1c9");
            when 26102616 => data <= (x"204a75c029c65128", x"7f3d6a6fe7a86159", x"3031ecd65a6758a8", x"1bd76f0e5b013d71", x"434d8ec163c43f7f", x"7d01e3033264e715", x"cf55e87b5661667b", x"2f2e24120292a433");
            when 21048275 => data <= (x"a956338f829d9f9b", x"6161df6eeef440c7", x"d15f1f51b0d3eb08", x"94ff5c5bf81fcf89", x"cec5624b2799dd00", x"2bc51b04e868bdd3", x"d38e90638fd91343", x"60d99a0bd20c4ac3");
            when 17275886 => data <= (x"ade21b64ee883668", x"c6d8d8e5b072381c", x"64697050cd5ec495", x"a90670d7f2c52875", x"17506e92d4fd4b65", x"d2ecab96e289ca81", x"195e073564a66a75", x"f51b3613b7626bbc");
            when 19598661 => data <= (x"9546876ed9fd8f0c", x"d21883d2675f59f0", x"3e54c9c646a0a7b7", x"1d349d1f3cdd8e9a", x"62ae67a8d3a214b8", x"6c3a511f7a2af1f9", x"b65ecd3ef71241ba", x"0fd160e49179e7fe");
            when 9189485 => data <= (x"3b66fef7260e7773", x"1e5e6431791ec5ef", x"95a99c245fd11d33", x"50b308cc58d14395", x"0cbe8fb2529892d9", x"dbce8a7a3458bc66", x"e004608b1cf4bc4c", x"58381d33a7104c19");
            when 21822581 => data <= (x"93a792a14442b3f1", x"baa22b15fa97f2b0", x"e432b8b75e520a07", x"2bebf18bf0200365", x"6d220fb84ec3fb9e", x"491ceddcca0d2e18", x"d28a549e6a7d33de", x"1d0928ac98209a4d");
            when 8021326 => data <= (x"1c65fc5070a49026", x"92418f3f082d37bd", x"6071818e331fcbfb", x"acbd8d4b3cb7d80d", x"3a0a882a72510ecb", x"714a66485ebc37d4", x"65a1cced89c51bc5", x"be26eef2a884255b");
            when 4859223 => data <= (x"a80062c889f9c012", x"fc674748012ec4eb", x"bc53a1293be77bfd", x"bd8011b76858d5fb", x"879328144b9467e6", x"8d6f9b9a7d1e62bd", x"180f894dc9a3f990", x"d9497d4ad9485d75");
            when 20416360 => data <= (x"30bbbd3eab87b345", x"c43bab500d0b44a5", x"3edd9975a3afad22", x"46521f2db67f06ed", x"23d64fdb76bf5cb8", x"c153c9cdb49dcdc6", x"d11156fab7d9f550", x"a0fab9fa581952c2");
            when 1023327 => data <= (x"992d415f8db98970", x"b2b5891d2ebdc9f3", x"e354dc93bb12f9f3", x"96b9982b587f5a9a", x"14ea776a7fe30a68", x"3028c3e2fdf578a9", x"a81dace2da7f68c6", x"89999a1d1795dfb3");
            when 6879909 => data <= (x"723afc29935cab19", x"e7c401a370a793b2", x"fb458adb4b67f013", x"1751d879107c1123", x"c416ddb516ead8ae", x"af4326ff85935c5d", x"b00137b1330fa506", x"133718980f5e1ac9");
            when 1248700 => data <= (x"d555caaf4f590f1d", x"05235f4aada753c2", x"13db2de0be1e432b", x"80a1fdfbf87a3563", x"785b5d370d0e2f62", x"4c3dd8b2583d3e48", x"54bf51e9e5207bb7", x"4b2b7f7fb6f16ca6");
            when 8411212 => data <= (x"777a3c5dcf7db924", x"938314b06e82f091", x"700b93a7def9081b", x"3f20e45332a52bfa", x"80e6f2332b807679", x"9fcbc3cb284af027", x"76c37ee2058d99bf", x"692b65fef641e1fd");
            when 11419185 => data <= (x"1ae5b0ae868349d8", x"db1a12f115f38b07", x"b15d7167782e3e60", x"fef8aa1cbaa94213", x"2505f4e92ccc93b0", x"74146ca9c35d14e8", x"b28c09e2f0e5b28b", x"18eb3a2416d6b2f4");
            when 18300951 => data <= (x"e718ddf9818631a2", x"c743a7ff08cd768d", x"768bb6d7fcb48908", x"1132b36539206745", x"7cb567fa27f2f904", x"d2c621119005bd42", x"6c7651d5a9d77854", x"973806b336926bfd");
            when 16320375 => data <= (x"f2161a43fa48e94a", x"e6f78b7317ba5348", x"35b307557452c747", x"f5c1a202475d09c6", x"6c4730104a859320", x"c4ec7face6ed8541", x"f17e8671990109ff", x"a42e8caa21b1b870");
            when 32178189 => data <= (x"c10cbfd1befea856", x"702191b0d7834d8d", x"d929e80a0be477cf", x"854358def8d7afcd", x"13bc8d7b5899715b", x"8bf345573c073323", x"c21749de3354e79c", x"ef71171c80aa12b7");
            when 11346066 => data <= (x"cec259d4e4876964", x"9302088cf131c3a3", x"4c97505960d84f11", x"7bc491e1af7bd46a", x"e476159026104a55", x"e5a38617b74109c0", x"a5957b8b1cc1d700", x"fcf9b9d832a02f97");
            when 20366733 => data <= (x"593d026ca54d1135", x"e0dcea6d091316f6", x"bb3e901c4d393f98", x"29c42de9122ed0d5", x"ab7a583a20fc422f", x"74ca99cf72efede2", x"449f0491eb05a827", x"cf85be9ecd6a292b");
            when 7701267 => data <= (x"2e435be5f0dcc9af", x"c1871f092d46b377", x"154578e15c960e72", x"f14fb4411f47be76", x"9b97e518cd46692b", x"65ce0e0df2011673", x"636f0c5cf07acad7", x"d170a0cdb2f759dc");
            when 3262955 => data <= (x"3429df8dad6d8ac3", x"4366a207ef2c614d", x"f1d205625d4124f0", x"24b2761284578b4f", x"b943d872bba4f437", x"4e87f563b2de7eb5", x"55ffc83c2376e778", x"f8bab64ca7769e5e");
            when 22398151 => data <= (x"c0a751d8bf824af0", x"9645df3cd8efc63a", x"9af4e10df8c1ea7a", x"4a10546b4661f473", x"2ab770d58a986d2a", x"949b2e5be5ee9bd4", x"473f6db97a62d242", x"6cb0a578541bed90");
            when 26700051 => data <= (x"3602eece4440b11d", x"99f61200d08a177b", x"a104906f62adbfc2", x"f6b72d8b14647e6d", x"69ef43ba6532f365", x"1fa58759ac30ca13", x"f03f3f5752fd0d73", x"23fa9b7a9cb5f2b3");
            when 25217972 => data <= (x"e672a80cf8e263a0", x"25e949a0e141e1d0", x"9e0580d18af2dd5f", x"58e6248051cd87eb", x"ab805e752085c4d6", x"b12489ff1c8006bd", x"1e37e2880b0669ff", x"194aad9cbcf448cc");
            when 19359838 => data <= (x"1b22623b74a1cc7f", x"509a30ee2118eeb4", x"24a7012b16d3d13f", x"b848d4f6f38147fe", x"9a80116ccc9b5124", x"bd80d5d956dc9fce", x"ace27d26c4133fdd", x"67edaaeb7f9f0864");
            when 21179406 => data <= (x"cb0d31320c9677a0", x"2287a262ff21c1a8", x"7e3613d5c91211e0", x"b52cc011be58405f", x"59504a32f292c22c", x"afa14d427eb32159", x"0826e8e76681766c", x"d8f4b9cf0bad2e47");
            when 29613180 => data <= (x"5dd9fb225637a981", x"0f30ffac6451b659", x"25ca8c0e524f9a6b", x"2d4113479789f4e9", x"c60602267e7c5b65", x"9fd552112dc94446", x"4765c5d2bf0c381c", x"6d7520834102425e");
            when 21781235 => data <= (x"15be0cf9da02addc", x"e12545f026c17a9e", x"5c73a4904245d5c2", x"9bb990e9d15f9812", x"c44934e3ca7434f4", x"639a4ae0a2a845ad", x"888ab926f9a9db46", x"0cf67afe02c70a15");
            when 939900 => data <= (x"2860aeb59cb00c0d", x"bb4b5dc6f2e4d15b", x"bf4b37e67c158958", x"cd9f481e14e77589", x"fe461182369645e5", x"2810711d2f6ca450", x"f876cb226913c5ea", x"ba0c7762d3da33ae");
            when 14939958 => data <= (x"59c7017032d69ee9", x"6df5804837025fc9", x"b36202d436b8c31a", x"c6e2425137932200", x"b39e4be637e37364", x"3bad53bfd76af9e8", x"353bfc0aa76c4430", x"2362f0cd489f2fd8");
            when 28276861 => data <= (x"5a27dfd863428bd2", x"0b735c6596170211", x"f7efed5f95f10ac9", x"77cad8d389e48600", x"b718cc8bf26b54ba", x"02c1972d3bf54739", x"5178af21565d7d57", x"cc79b7cafc1e8629");
            when 27508015 => data <= (x"40ec5953b7ac80de", x"8b3c5bedc9ccecdd", x"225f6e43810c6f08", x"d2c7a4456737e946", x"5791d99f00b22417", x"dc9fab8170ba1308", x"bf1b8076f11f810a", x"e275d0f8e1853e09");
            when 31640519 => data <= (x"0ca61ed109376e94", x"7c1e718e2c44fac9", x"583cf391722e045d", x"5b2518eb49351240", x"109c8f967dbae8f1", x"e3eeb018d6f78f4e", x"c1886180f68ef02d", x"c35df89ef113e14a");
            when 22460451 => data <= (x"54b3a7c5477f07c8", x"6c1c3a630fb0890d", x"171ecb2970d6cb70", x"bb02654401cd1cb0", x"9fc35379200f5278", x"7806bfcdedd8feff", x"6a4a5e04b00d26b8", x"672e8af9c23ab555");
            when 13629944 => data <= (x"66d09f05dc836938", x"1df20080c76461e4", x"351fc091e5f5eb8f", x"a03ef63f6b95c75e", x"6830b9f46b1198f2", x"088fd0b39aa825b5", x"08fce0112d181641", x"63a141983c54f674");
            when 14293756 => data <= (x"695e50a93ff8e46c", x"eb4d6b1a149ab021", x"b0ad516ee54121e5", x"9cc3a0939fc5f989", x"8edcb581ce7a3aeb", x"de522b177273eb3e", x"e082a813229be457", x"64e24d3210162a3f");
            when 7737181 => data <= (x"ed0777c1d0fef199", x"b90f4837cbafea15", x"7afcceb4a563adb7", x"da35efe651bbfbcf", x"d3ea08c4c9082979", x"39438e13d984c349", x"2b7f6bd105e01e6b", x"48b6645c1ee14406");
            when 31730150 => data <= (x"1c15fb0779a58e47", x"45b68d22d3e756cb", x"d3ddbde120d068b1", x"f8b27fdafb365184", x"004fcc1259626a8a", x"d94937e64f239894", x"e35b693572374448", x"1bc7b3d8a17411b0");
            when 31741081 => data <= (x"e496864c9d22d153", x"00402aacc5e33991", x"1bd3097c015daee9", x"d47a6532b657d6e4", x"ba74a8486d7b7fd9", x"c31fbd1d1f253511", x"a7b252d885f46165", x"76278c69e3dff583");
            when 19716423 => data <= (x"d6b17dd1fa1dfde9", x"77aba69f7585174b", x"54a0fb2eaa852b58", x"a52b36dda71259da", x"5601b497b7faa5fb", x"bb6e9555774bb04b", x"a18f3efea21292a1", x"ae58e014a170362f");
            when 18382816 => data <= (x"c4838d70b18117ba", x"12cb414d7bf33ebd", x"837741d5cf546540", x"0c0a90e771d9323b", x"250acd8e0b1bf00d", x"4322c0f9058e56fe", x"51552b90bd880665", x"d2acf5877a0e5506");
            when 21780876 => data <= (x"428f33d7280dece0", x"4f4eb9da763b9b8f", x"7f466f6aaab3c9ec", x"bdb662cb14dae56c", x"7f3d69c0a20ff0f4", x"93c2fa4aacd8615c", x"be99a1deb17c82de", x"eb25b7f97972be6c");
            when 26433021 => data <= (x"2ba3a00bbc7c28ea", x"6570776d527ddeed", x"4fd04e55c2888126", x"c2c7661ead725e43", x"c0442ceae2cd2b69", x"e2e9066379e61969", x"a3c30b50fea94ccc", x"3e260d419bd765da");
            when 4181065 => data <= (x"9c9faf60ad325866", x"fc1549703124af9c", x"e6d0627bbd30c3e7", x"1ae8796bb9843d57", x"8c98be3b473e44f5", x"440c1e5db827a878", x"9150072b19abb8e7", x"c0bb15ce829ece41");
            when 9622337 => data <= (x"68afc5a8a795e125", x"8cda67ef33fe44c1", x"ff49bde0c0c611d7", x"5a4b0684d024bfde", x"eccd1d3997ab9dfe", x"7af3d56b67b90d67", x"b72c6f043752c54e", x"ea417d7180dfd213");
            when 27947345 => data <= (x"34c6ce2008b802b8", x"58b5ca769a3661cb", x"cd6f26df03bbd386", x"593d290b59ff4a0b", x"01f0a2fd9f194c30", x"37b77767f00e790c", x"4176328e136e398f", x"27571938d3267842");
            when 5565886 => data <= (x"cc5167edf99d846e", x"ebee18f47ab5ecba", x"3a731a443861035c", x"1553e3e30de51e30", x"1a94af8e186d5b77", x"fec83c932a326edf", x"4517bf15d6db9448", x"7f9c700a1ae3ca23");
            when 30065981 => data <= (x"7b1ed96835e35d75", x"a8f51df0cf76c3cc", x"8dc47ad6f9e89b16", x"128b68381ed3cd0c", x"93f68d92f9b7a8b1", x"f49fb0fef37c2fa6", x"18745cdefe6c4aa4", x"745750ce5182ab96");
            when 31307092 => data <= (x"b8b0cd384b8f7d55", x"a8b181137610860c", x"c9fac50253310780", x"18cb41a6a7bbc877", x"333eb5b2824a7345", x"998e7c3e8a3b0985", x"efdb004609e2e632", x"739c604e43d22d79");
            when 22986982 => data <= (x"4463fe902c7541e5", x"683e10654eb79f5a", x"cc5e7a30e0aaca44", x"eafa991d82012b30", x"6c6520598d7de368", x"fcd2359e31637118", x"0c7574cce2a23c8b", x"65c77812243e6998");
            when 27892257 => data <= (x"497dfb2174d8ab5c", x"189a4928ecd2c81d", x"625fadb6cdbb7b7b", x"c066ce5a80f1ccfb", x"3f412841744daa5a", x"29ff7a9768cb787b", x"f8b54095e87b0339", x"f19873e38510f881");
            when 21135651 => data <= (x"ed36e6d58895e073", x"7101f57519f6ecae", x"dd215c0b9e594e9b", x"c8a6e8f6978da459", x"88eec112f1938164", x"6f208b166f2f9ca4", x"82b49d0e5c6dde7d", x"c8acd5e5adfd00e8");
            when 26289482 => data <= (x"1fdb8063f0688832", x"ac9d6c9fed5f925c", x"431d1389c2741a47", x"47793dca75aa5f90", x"9ff592ee0b58a367", x"2c8f9741368fc639", x"4cfeb2e6cc011c9f", x"417d6119ab83ae60");
            when 9718581 => data <= (x"d56dcd5cbec82709", x"36f95f695b7f6c6f", x"508bebaedab8fabd", x"395d9e7543009c6d", x"b63a619fda79d34e", x"04ab82dfa6be44f9", x"11a9485348a6878b", x"a7b8e84372f9f59a");
            when 13326563 => data <= (x"750b978e555741e2", x"2ba4b3ae79e1cf96", x"0b4387d9a5ade7a7", x"5e4c96299c839254", x"1d5b67517f916a4c", x"9678b738255365a5", x"23bb6c78a4a28bba", x"b45028c1a26e864a");
            when 18134080 => data <= (x"c47552cb0940d797", x"68b51fe8077432d9", x"f39507ec42eed8f6", x"278001aeee175891", x"0200618b97e993be", x"510758eaab9deb37", x"87032170f967aaac", x"a7d9c885516848e7");
            when 17948530 => data <= (x"d993e5d4d0d9f200", x"a15c0e48265a6ebe", x"290c62080b25e7ff", x"7d5151d27d66f295", x"4b521e0b59bf0a57", x"412a1a3ad9bb00da", x"883a223d3e6edce2", x"c793c8bf46805fff");
            when 9745695 => data <= (x"b3a2f32bb43e1523", x"2a0a20e0f369983e", x"5c3a2a39e28e1c9a", x"1db06f7769a59cb7", x"7e5f684ba87f7558", x"6f5d1c0775ba255d", x"7ba746613daccc52", x"13c95a77d5ab47a5");
            when 25135940 => data <= (x"396fe660f71a3b64", x"19f6148ee2e118e0", x"121ba98ed73e1d87", x"3bc775da108c238c", x"98314bb4607a085e", x"e3a03f59e8dd1794", x"d60aec15911fd933", x"502dd7ca373abdfa");
            when 31963334 => data <= (x"4a49f7206f3b2001", x"07e850238a208646", x"4174b457d8b31a82", x"fb5fbc9e6a1d9a6a", x"46e0fc16b48d0772", x"36e1357bcce87478", x"d198fa79eec851d1", x"69c01e5430f5d7a6");
            when 32458044 => data <= (x"997b44fd309d0494", x"5d732926d5a0efe7", x"5e3d08bb285e2b8d", x"be9b29367bb53b06", x"8d2c256d68a27d04", x"5ca5894df8809dcd", x"d7f6f20a1bc72804", x"710e040fbf921b76");
            when 22223214 => data <= (x"08cd5886a23f0890", x"7a0906273d281a72", x"e33d578bfbbb6be6", x"d7ceb4c0b092a602", x"85a02e57d7d1901c", x"50856e7e6413f6e9", x"f147f9962580ecf1", x"de88259831b73c45");
            when 27636428 => data <= (x"84aed8a4dd6943f2", x"0a908dbdff465e62", x"ffe115bb51b6b378", x"a00d6a59796b9108", x"db52189b1ef49bcc", x"8634388e0b94e547", x"6f48282792f84a77", x"ca428d9adbcfc85b");
            when 6198051 => data <= (x"7accf2fc7bfdaddc", x"3abecd12db360e07", x"d18b3dbd975e57e6", x"12e373ea26f5d43f", x"b4690117223d65cf", x"d74463aa4ce14790", x"f6688bb0208e0421", x"6b608329985a5284");
            when 2018377 => data <= (x"4b0c1cefa59e2cd3", x"b3e8970e1f82243c", x"df0f7909767bccfd", x"e5360f9a6e11177a", x"16c8fca8bfe42c08", x"a9c4710e70eb5bea", x"32275d512a642e68", x"2268dfc58e667973");
            when 12789331 => data <= (x"d268ca557213a4ea", x"45968ca653f849db", x"99dcfe8934fb4955", x"d4bf457cdf97267f", x"129c1b7159949585", x"076b043487bc4341", x"531edb867f9ed2ba", x"63041d58aa2e16fe");
            when 29923364 => data <= (x"8f0e5b40b2a0e882", x"bc73956e13f8102e", x"9f070bf7a748c0f7", x"c9036341870fc410", x"cacee47d944b6d30", x"5399135171dc21fa", x"555e4e1372568c59", x"dddee47fec37478b");
            when 7951141 => data <= (x"b438805c56b24105", x"f897f4e1d7aafda6", x"615800d2ca109578", x"817910587ad7a5f1", x"51e6f2dc83cd9eae", x"18208363317be7b9", x"f8c44fdf4c535c89", x"d44211e9bcaa4d0e");
            when 4304613 => data <= (x"d762b188eb0769ab", x"a9b201dc34af1dfc", x"bd0b85e29ef240b5", x"136827f2f21b7c6d", x"175a7f8d5032de90", x"49f8c752b8c3ea13", x"974dae092584d82f", x"18a203878e401932");
            when 12399144 => data <= (x"87368d9e8251dda3", x"3dc2f46290af3247", x"64310c86fb42fc48", x"b09fa67552798ec6", x"93529bcbcf255d41", x"94ac45efa8927dea", x"8b595af92a44aa68", x"f5729ed5fa072310");
            when 22073596 => data <= (x"ed441efc6d51cc41", x"8adef905f864fecc", x"08249cdaa0192f49", x"6920d59094e9acf4", x"9551fb65dc3e2673", x"82732cf50b6cdb98", x"4680bd5b48063666", x"674b7b4ca4679ef9");
            when 4783835 => data <= (x"fb3b0fa5658c3252", x"ed167025a02e0631", x"6a8d9bb9bba86d2e", x"656030c15843ffd3", x"1e386917a5cec67b", x"4d110b68eeff7862", x"162bf17d29becd28", x"afe8c2edf8d45b65");
            when 6359987 => data <= (x"b941fbf9adc25efc", x"0ade28a95dcbab11", x"1a8176c021e9249d", x"67a839ec5008e0fc", x"d3f853964d60b729", x"ceb31746a4607a68", x"89b0bc13aaeb6cdb", x"2672203562df5db7");
            when 13349114 => data <= (x"360a5eec9e7ad71d", x"2abec379c30833e0", x"8800cc902e523445", x"8348b88da9d08429", x"6cfde8675f2d68c3", x"a8dd050430b97088", x"cad5ccd615d57dc0", x"f0c9956c9f0e76ca");
            when 14784313 => data <= (x"04df8d93d9baaf11", x"b891a9b6750f56ce", x"46fcc5ddd9aa6f11", x"0e5938c530046828", x"54f4926d37cb68d1", x"0202c515cb3b615a", x"8a203012fa479fde", x"870253375ac15995");
            when 29329940 => data <= (x"ee9cac3a302782dc", x"0c44f5e9598635b8", x"6c41f6812623919b", x"c9e844e39405f4ac", x"fcec2a6bd7919c7b", x"68eabe393cfa9068", x"b7d2319918cb135b", x"9788b6b5ad6261b4");
            when 28065771 => data <= (x"dfd19db8d0b2b92f", x"87c04ffd712a7094", x"8aef900f5711698f", x"2d3591ea4542a31e", x"8ad3e38a4fec2d54", x"24c7ddabcdfbdb52", x"c94e68f60719ca2d", x"5e8bd0ae8a4abe46");
            when 3063450 => data <= (x"658446070b84b281", x"a516315e81aef27f", x"ead31c8d2ac8d6f5", x"0d1021c50865c7d6", x"344a366ec23b096b", x"36fd08be9affd1ee", x"a0d87d6fba461be6", x"2ea1a3bb00a71eda");
            when 20594133 => data <= (x"11371de334f3cc1b", x"ee252b62c495f7a6", x"4bcd1a834852756e", x"6f711ac0cf9536bc", x"f13e51fdf9cd39e8", x"0bd8b0b245a7c207", x"dfbc5d6a40ac4b89", x"49a6e19462de68a8");
            when 19515455 => data <= (x"5c0bec7f705bc77c", x"7e0f024f71500f81", x"6f6e256c6becc233", x"4094e1ec0c975d08", x"661db04352d7d5c7", x"918c7502db830101", x"956e0f7bdd96d8ed", x"ed2fc4310a75ffd7");
            when 1566757 => data <= (x"c39d9bf7af1c93d9", x"8084b9c5204e4a83", x"7fed34da7b23c9ed", x"076fbd6fcab24b0d", x"69cf1bbddabdf1bd", x"1d38f3cc0dd53db0", x"84f6c2d5cbb16ac6", x"52b50ddb3d1b3975");
            when 22143660 => data <= (x"f61111ecd3164206", x"611fc9baa4667f37", x"086801f5a3f315fe", x"f617b6cd7b137e2f", x"f28815fe57f0670c", x"96f49ca12b5ea286", x"bca437a8ae002ece", x"0ba3570dcb309947");
            when 5246147 => data <= (x"5be448080ce0d350", x"587580938dce4e26", x"51970b9bbc071507", x"47c0d72de24b8512", x"2942a1e872bb1dec", x"2b106899e2b128de", x"a80d666db8c3fd34", x"a4f0d3bac5cec4b7");
            when 5718451 => data <= (x"240e4b32daa796d8", x"640fd78cc1b00df2", x"5f5365d6472adb7a", x"9affd385b428a70c", x"5cbecd959fd410b3", x"af14d45947e41e0c", x"9194cf5b4e729212", x"fb6e3d27699165fd");
            when 4493210 => data <= (x"ad6c277a93ad7a86", x"4b06d8326e9ceb6e", x"5e6a35ac9b6a4968", x"5d06be78321cf391", x"2f5171c526ae8064", x"c3feb885d6237e3f", x"f549e611f09b7618", x"7b92e56229b54144");
            when 14917728 => data <= (x"a490baf78d9e2861", x"198fed8cba0bb14d", x"a2edf2578445a80b", x"e3bbbdc7ef7d15a6", x"b92314e5b1ff76e4", x"37e87214fd1ccb3a", x"759c6cc133bcd870", x"b0aff4a373cff968");
            when 33337656 => data <= (x"fc992fd1629a0c51", x"c7b182e4c6901677", x"89074b3ce9b32f53", x"dff7d3b74b68e5bf", x"672220207c6966bb", x"0bf222c7c8aad7d2", x"a75c9714c0b9cc74", x"d593daa99e5bba14");
            when 18064852 => data <= (x"a583d896fb3bf4ca", x"98e87d44c825d7ab", x"24e6ab2e188d4422", x"86fab178adcfd9bf", x"7532253b28c48c32", x"20cdce26607a3d94", x"689d5420b98d3717", x"f544571085bbba1e");
            when 13473817 => data <= (x"01289b6e6c2c2761", x"2c5ba44074c16ea1", x"c9fab058a4fb3b88", x"757504d4db433db9", x"b50775bdc0cfcd0b", x"69b3d1619959e446", x"11d8f7fc442ca0d7", x"6d1091f51f6a979d");
            when 22591625 => data <= (x"f52bb402fd651e5d", x"d0458e2371c8196f", x"b0916ea13969591c", x"85e7776b7af87198", x"bad27edca90ff6b2", x"4681d90644ccd80c", x"ad26c52943cac50a", x"a58515e3f5ea0dab");
            when 26522244 => data <= (x"3c8077ef09281008", x"3b282715b556cfda", x"efe4663574921563", x"c9a1ffacf550b702", x"bc9a7095d9236d5f", x"f3929233a6a4002d", x"73060e109c0ea6b8", x"46f9d5946e68275a");
            when 23009875 => data <= (x"6efcd1acf7fb3a7a", x"4fe6fade98539ebd", x"d9c067942b4b571e", x"e12304ad9d45fe14", x"07b6175694f29212", x"9babfa91ee20c188", x"89246f4ea788fbb0", x"637fcc1532a31332");
            when 28122372 => data <= (x"a32d0724356751a5", x"7d6eb4e1a38c67c9", x"a0a6578bd863b043", x"0bb201ceac0a321a", x"6758c859442c1260", x"40eee6a74b4631f6", x"0bb2b0aa38e1bde7", x"67a6cc8812e254e7");
            when 22988075 => data <= (x"79559e14e38a621a", x"51411022d027460e", x"ca655d6d917b44b1", x"b2e3a5a0d34463eb", x"fbbda398ad092312", x"009bf5e2c13b48b5", x"257b57a8ae3f26cd", x"480a993c9cf25430");
            when 19975322 => data <= (x"c569c1524c1b9d2f", x"28455c3914662f91", x"4f40af08b467d928", x"b302ea34cb3dd0eb", x"7f606389845b5512", x"6999e968ed408e95", x"1471de278af55aca", x"079cd458ce377fce");
            when 5921815 => data <= (x"1feb531f1ab88972", x"f433704ff5cb9fa1", x"d1773d1e75effbf7", x"75d15ad5b5f30bfe", x"32eec3e2c1efdd2f", x"6984cf80f3529d01", x"7bbdf2c322ed0774", x"8197b32f3d4eeb6d");
            when 14898615 => data <= (x"8139c1d7f2642e56", x"9650bbd8f1ddf0d8", x"4002c95fbcf42344", x"8c7dff4e0edebe37", x"abfffabb52f2cfed", x"0fe454ff7a3b6293", x"abd83b46942ca2c0", x"6a7e6dc2fdab1592");
            when 1778015 => data <= (x"1cfcdeec552d452f", x"82ec07183c136bb4", x"2ff94bcab33a5252", x"4c3c07c3c310606b", x"e813d8511c0f4864", x"15526a8111c07cba", x"014698ce79ea5b9f", x"fac054d1f22ce8fb");
            when 4850560 => data <= (x"3463e9a3bc83f14f", x"a34c31ef84b2f122", x"cff9827ed691ca64", x"4e5d446cfed63c3c", x"4faa75722df57229", x"30d492ff0fb26225", x"4d2d4f053336f4d9", x"1c439f172cd0c932");
            when 15478157 => data <= (x"054948673b75fbff", x"d6d900b8acc77bbd", x"a2559ae9e0d63723", x"31c4bbeb91213e4c", x"f4b521e7a9d91317", x"42d4267089a2032f", x"28b0b38325b93103", x"0f94e523aad7f980");
            when 28212951 => data <= (x"f9007085330eb882", x"a9a1a910a84f6904", x"9dccd86a78689c2c", x"1b393f817c790a77", x"f0490b9e5301ee2c", x"92bd235c30ea7eb8", x"b9e793cc598cab82", x"1289e80a3ea34abc");
            when 16189841 => data <= (x"180d20de453578d3", x"d4960d8e5902e79f", x"b7c7791fe825a1a8", x"0eaa245500e84f57", x"86f2ee884ce5a705", x"a87776979efe2af9", x"9d720c01a8a8564b", x"285cc0e7e1619bf4");
            when 15476465 => data <= (x"f15fa995d968d12b", x"25b1341d2b4dfe24", x"ef2a938f3a2326df", x"0194e0283b9a4bd0", x"ec77f0ed8efa9788", x"030fc50f17ecc259", x"ceec449a176e0b63", x"39f841c71616ff9b");
            when 30063269 => data <= (x"f58ec9c387fc361e", x"70f7093d6a014189", x"f61c5531d4da150b", x"fd40617b0354bb69", x"4d37af773fd4033b", x"f1410981519dfb18", x"105607e67411771a", x"af20a44aa3739250");
            when 4484630 => data <= (x"75b7421c05133ca4", x"cecbae1802a70a56", x"266a9ab75697c3b3", x"ac4f5cf486f0f17a", x"40467a2c8d1cd55e", x"8450f8ee9d668009", x"7219a6b455f92d4a", x"e446eb50b57e4ab8");
            when 21231671 => data <= (x"4db9989b349ecbad", x"18a08d276b82e436", x"fa4a22a70301c3e9", x"d4e998c84fdff050", x"4db209b0238fd03a", x"ac4f424d921501ca", x"dd2ad8137125ce2b", x"adafe5266b667310");
            when 4143990 => data <= (x"2abbb28f5f3018b4", x"f979cb15a463e4e0", x"d1ac8d8675d85c3a", x"252094de9e255c59", x"542dcbfee0a148d7", x"c18b916eba414517", x"2ae78c1a0ed96ef5", x"a3739944ddbbe47d");
            when 30261368 => data <= (x"1e059941747c9e4f", x"92b47f089e30a4af", x"94e8593c92004e76", x"d237a45558112d7b", x"78fa541756066a58", x"74eb6b3419e61ce9", x"d2a3dc4c7a772e81", x"e88eec3f9f7d4a5a");
            when 22432440 => data <= (x"0a676292ca8c70b9", x"9dbd28d1a7575836", x"0efb30470c38e0f9", x"848e25a519027883", x"81a696c2ce2f33a0", x"c51fff7d3e113c88", x"9d6cc748b86c930d", x"0e6f6e630595350e");
            when 14791333 => data <= (x"048c3c619eed7240", x"2e520dd3192c0c55", x"a1722869be7241d5", x"a2312ba95ed00f88", x"7a5ee66aefc16e8c", x"eb924aaa370841a1", x"12d220e54fac7b20", x"2c142c0738d4b3fd");
            when 8249247 => data <= (x"8aeac5a79a9ab8f1", x"be3cdd84a4829eed", x"6c5c19e053fbb9b5", x"16972cd3775164d4", x"5ab7ac14f7095fbc", x"21b536e50964efb6", x"62948340ecb08e8b", x"6c4332d708e0af2a");
            when 14320234 => data <= (x"327ed3581f0dbf95", x"ce8a4d2cc734a8bc", x"d4c42fdfd14bfafd", x"6880bc1310602500", x"00d08f4dbd13de33", x"e6c90edb904d5ffc", x"605ec99906936b3d", x"29427f2e65f281bb");
            when 28530195 => data <= (x"94f45df15f0aa575", x"c9c3f374c71f66b1", x"dbc2976f2d57c0b1", x"4fe76d472f63d7da", x"df7ff652544b1296", x"31cf636fe26d8b50", x"6bd00d1012fb3f6f", x"bda9e7ab88522750");
            when 27305517 => data <= (x"c433d065e8b06190", x"26bd8980103e1a1b", x"d5fb3e2bb2819780", x"44d61f3838b8c94a", x"ae5a39adc6d93921", x"3483fc20fc1e17c7", x"103e0efedf24ce58", x"8bb842be51e65ea9");
            when 2620272 => data <= (x"e352e5ea0523c297", x"9f34ea61da5eb135", x"2b4e16db21437e00", x"5e6710e6d15de899", x"d98cdf91b5f34bea", x"2bfd06c40681f595", x"e1dfc8c26f6fede5", x"79ce1c03b8014054");
            when 21158278 => data <= (x"66590b36cb58f063", x"284383172c18fd66", x"0cdda5074f2b2117", x"79f80b9ff008fc71", x"c68a7c3aa770ac37", x"21489e1db29163d2", x"0a78e6b6a080f637", x"637d634190a54ea4");
            when 29938533 => data <= (x"669d865feb65c938", x"e23a77d699b461e5", x"10606033613a678d", x"ffb8c5fcf3c1e24e", x"b3c6416830b68edd", x"0ff96b4a601f3cea", x"f44d3de54648cb60", x"576331c5e22fb04a");
            when 18806822 => data <= (x"a7b9efb9766e3d43", x"97990b94e67080fb", x"417a429878f03a16", x"665513b91aed6595", x"c2188771588ba32c", x"bcd5dc11b93316cb", x"aae19bfde7a7c172", x"124f1dc6a0e6945d");
            when 25650703 => data <= (x"2ca2e86fbba95edd", x"ce3e1c65e10bfe42", x"e21c3f6523a4c2f1", x"8cbf472deff244e8", x"9e87f7016d9491a9", x"893adb9e04e8aae4", x"4bf5217bcf8ef0f5", x"56596b41d593e9bf");
            when 14733298 => data <= (x"5b23cafc3536155a", x"605c7c604feac4b6", x"3c6b46c9f1856a0b", x"80481676e98f7262", x"bfed30c756e557f4", x"632fb9b609f5d267", x"83611cd014e2ed97", x"1af8d79340c61e07");
            when 4692942 => data <= (x"9b6aa95472fd22f3", x"44e7f9de1a88f35a", x"c1fc2242d5821904", x"c9e24d9b4bf8b3bb", x"8787c0634bbaee65", x"98f5e9d155731fea", x"7e869b73afd54aab", x"95fb04798648b488");
            when 24139325 => data <= (x"742a6e7c8c75812a", x"020693939ada4868", x"5ee0f3ff0aa7c6b8", x"94dc19179799f938", x"43e622df1f193718", x"f81ddd324811cc90", x"30cb6b935f306b42", x"5ca63a761dfefe2c");
            when 2329620 => data <= (x"9e90241bde7f35aa", x"f49de89bff0ad596", x"e0ca3cf0009475dd", x"116fe53221def32e", x"3bc5fbbae90cadf3", x"64464e70d909d2ac", x"bd89c070bc25b9a8", x"fd208e0f8f1465ec");
            when 9959368 => data <= (x"a2af66cdaae40fae", x"4ff7daca13c559e0", x"77db03b798c90f07", x"9ebc027b4eed5d80", x"53c2e91fc59f0b98", x"e6033b7214eef17d", x"b3ccc6c09e7a5d48", x"c4f98247b5c4d802");
            when 20370116 => data <= (x"79392076f5029ab0", x"177cd22ad564021b", x"681fbcb12c2814b8", x"8907e7524b9bcc6f", x"466fa15777bdf558", x"f17bf1bf2d0c7def", x"95bf4c7b046a8312", x"4aec5b017173a428");
            when 8698622 => data <= (x"15d983bf201b1358", x"34e21ed64353b6ef", x"f5037e609dc4afcd", x"9758ab8041fe0479", x"9853b52bc66a8709", x"4278cedab828d3ae", x"37815a0096e4a0bb", x"d7d76a19725e496c");
            when 27931676 => data <= (x"f0fe96868a8a0891", x"6797bcb11bf18368", x"5593e454ab2e0b6d", x"93134c900494a210", x"018884c041ff84dd", x"1db01d785e84734b", x"d0a9ae2d606b8145", x"4a1405188fde5899");
            when 19931885 => data <= (x"d3ee63fa5c67da37", x"bac4947e666097dd", x"3e79afdcc3a265c6", x"5b4bae7939880131", x"579cb33307f8da29", x"f33da057957a7374", x"95ea366e07f3c4f2", x"1723cf5a61d90eec");
            when 22587036 => data <= (x"8d0bedc290f44c15", x"5dfe82065a0a7632", x"7bf24673da244e1b", x"fd3d7a2f707d0502", x"afb2d1e48785186a", x"1f4f8939fe91ea5e", x"524ab2a375953e16", x"5111ee76eaee89b8");
            when 17281092 => data <= (x"e6a929919383b1d9", x"a499a0e13be8cde5", x"a9faedcd417a2ed8", x"56afda03cfff001f", x"fde560d66e6d3962", x"480eddbcc230b4fc", x"1bbeba03794ecb0b", x"dfac8cc9b3791612");
            when 5819649 => data <= (x"47f5751a0f39e265", x"18657e7dcfa666cd", x"fda9325090d8643e", x"bf36185c2b8be7ea", x"7128377c9c8ff105", x"4efdad92feee5894", x"54733053daafd6be", x"ded6b9020f192350");
            when 21520120 => data <= (x"6fbcb64a7b26a484", x"a4793936374352e9", x"4088630b8f158f3a", x"4984d1313d5e7c8b", x"5b045b8deb71251a", x"5b16c9075e656774", x"62907d9dde6fa3ab", x"f81cec6863b296ed");
            when 17971433 => data <= (x"8101ecbb4d51909d", x"dcf5e71c406895df", x"f674bb2f2c92bdea", x"3fe3b3c9d25f710d", x"19d6e71d1c30129e", x"7b27ba12b5464845", x"5957889f744e7c0e", x"63e1db1576732fd3");
            when 28442226 => data <= (x"26b4c2d51935b46f", x"2473a77400422e4c", x"11d83de0d3806e92", x"982785bd31e29f26", x"f20d9abc8388fe80", x"7ec47ff5aa732b27", x"41e95d5a16e172ec", x"6ec0500e695b0704");
            when 16730202 => data <= (x"b5b4156f44b472b1", x"50655d0b976249ec", x"625f90689367aba9", x"e612a957181ebf3b", x"c571346494ef1446", x"aea74f26865312d5", x"1bc880d4fa86f8fe", x"6f7eecb9d6c01e28");
            when 33138198 => data <= (x"4046d62dc511bbca", x"328497ba5e729a7a", x"57cd218cb47ae726", x"232d6a48671e8a60", x"e688bca767093174", x"6deb6894b53519fa", x"efc2532aeeb31a22", x"2dea5eaadd42b3e7");
            when 4303710 => data <= (x"1851c28a7b2983a6", x"84e49315e3dd186c", x"6124e45f146a7b71", x"e94b1ca3097b48b2", x"a08c236960886a1a", x"955bd701840ab339", x"7b3ed0c7273759b2", x"fec985be63acdcc7");
            when 31236494 => data <= (x"0bf373994db965a2", x"f1003580daa3e071", x"1470510f2f04ddae", x"fee2b69e5ee6d6eb", x"bc4fd4fd389f89c1", x"7cb3f0025e1bf67a", x"3a4a5792fd93853f", x"036ed2ad1e3aae05");
            when 25968760 => data <= (x"c26227a2ed7188df", x"e4f0beeefc2b8dfc", x"189cccbc2b181014", x"9738a0b56f29948b", x"285026405f23af28", x"0de9d7a7870b583a", x"2b180433c30d05ef", x"dcdeb89747bfb0f2");
            when 8688657 => data <= (x"5ea1b5bb9069bc8f", x"402587fc236779ab", x"1d1dc23d0bc59ca4", x"0b35db9cbbfbda81", x"0d7caf94d3768f64", x"773aa7e3ab1bab3b", x"9f94f97242c0a1fd", x"2bad68992b66a94b");
            when 17763141 => data <= (x"5626595184f0840e", x"be1559e3bd7b283a", x"673c84a7041c8ea7", x"f952194dc57eeeae", x"6fdee8c8d1713a3f", x"f6f95916f2306e3f", x"2b31829d0a9ea493", x"f03a7c0f013d0af9");
            when 8945210 => data <= (x"79de8c0f20144816", x"a985f86b5deb64dc", x"e1d8ff849eecd1a9", x"4c514a42f7a834b5", x"b92da453718edf66", x"60df558479fe9c5f", x"2fd6f02b276d1ef8", x"74b25fdc4f1eb412");
            when 19577361 => data <= (x"78510afc82424a87", x"9ea001c1d7a9fdb7", x"4beb39f50885f6ab", x"ef3c0d106dfd8d62", x"65f5997e8b115d50", x"3d7dbd4c93000563", x"bb3520e6a8b7fbdb", x"188b1df7d81ae639");
            when 11282543 => data <= (x"2656911eb8820b51", x"e617c926b200c0b5", x"202d660333be3903", x"4f3120cc35ae97f2", x"2f2ab9a576a37de0", x"d99474af2058e21f", x"d34313c39f800cfa", x"bdb8059a3d9ddda2");
            when 2796246 => data <= (x"9cc6258917991eef", x"cd2df15164b1a979", x"631b2f30f1f986d6", x"84936c544770b432", x"9cbd19820e248d5a", x"047e4c7720cb6a16", x"587e6fce95d9901c", x"75be88eb151150b4");
            when 27346566 => data <= (x"a13ffdd0b88f3296", x"118917f8d6023717", x"535059a6095e68d8", x"9d241acc08171c74", x"e5618d54b08c7283", x"66603f91de389eba", x"a77532dd9e6fe9fa", x"8292a2b0e477e901");
            when 9445269 => data <= (x"f5e0256d7beeb935", x"67e7fe43f72fa3b0", x"069383520a9755c8", x"e49eba367006db33", x"728d5d490961323d", x"246b5c927aa5b6ba", x"b4c017555bab717c", x"7ee430bd9896626d");
            when 28631567 => data <= (x"862afdedefbdf1a4", x"c311e32412603b9a", x"627363a1930380e4", x"9c9e708c64ad4bdc", x"6173974c17acb7e6", x"75553bed2228e0c3", x"34ca1278936bad86", x"e4dcbed6627ed8b4");
            when 3747012 => data <= (x"ddf4f11cf50f0ed6", x"612d6a29993b81af", x"99b23f19e7b8b8d6", x"443cfa8de668a13f", x"bdc6e5cda595987a", x"c14158946570e733", x"ffab281c318f2f62", x"55694710522cd074");
            when 25178916 => data <= (x"30e1a006738a7d4b", x"0995586a9eaa3482", x"2069da6f34760933", x"b2d244b8bd76cab6", x"67573b151c30baa3", x"08dd7f0d0866774a", x"1246b27cfaff5ce5", x"8fcbdad00d55d552");
            when 4146340 => data <= (x"fb27bf3239a524cd", x"2eff66c0882bf2ad", x"1c508f78d0b628be", x"ff7d9636bd8ce9fb", x"fed3c025839fa881", x"eebab8e9af23a9d8", x"f25704bba5d39895", x"11faaa29045e0b97");
            when 15079107 => data <= (x"7c22cf3354751e2d", x"0303342db594d8b6", x"4f181aa34fbf76f4", x"83ccd983862feac2", x"2bcb33560625232c", x"779274da68d623b6", x"a9ad4fd9308ac26f", x"2a25979f0ef5d5d7");
            when 16959522 => data <= (x"e6c4851af96d3cea", x"979ade6a5bf13b65", x"c78d3d2dfc6058cc", x"8d9f3833a9128d39", x"7351635c297c88e6", x"5fa626fddddf72f0", x"26c929e7ff3d072e", x"56043d2deb8e5281");
            when 14928503 => data <= (x"2c990d9c48484ba2", x"34a5a6d832017b1e", x"45f5a35e638b2294", x"476f3cde1ca7bafd", x"ceebb8f020738d79", x"035303aaadff43f5", x"d7e8caae20caca27", x"8de43e5a506726cd");
            when 25681876 => data <= (x"9f365dcdb9cb6534", x"9147bd55834742b3", x"877768f2cd271f9a", x"d0ac863cd9c814af", x"6534bcfcc3bfaa50", x"74395f5b2331ed5d", x"4355b60c1de8687f", x"bf404f35dfb88d98");
            when 2204459 => data <= (x"42a4e06fd724ca96", x"686938b75521057d", x"2e11f82c6c27897d", x"c2f125106d8162c6", x"e3cb5039f3274191", x"747ebffe0746136a", x"374cc181ac129f99", x"6f514d3f0957e674");
            when 11683902 => data <= (x"4916e1c5ddb6bdda", x"3e63d26b1231d8dc", x"be6f630db3049226", x"535af75e93d15845", x"d34c3b3a2bfd94a3", x"0c089a102d80122f", x"9867a8f81e946bc4", x"fda02cd4ba917fa5");
            when 21189371 => data <= (x"6330bce6f8ea5af4", x"7c122e2ebca2cee4", x"b6e32d27369e7a1b", x"6a6eab2aedb723b7", x"754467490a083b52", x"1bee62d8a278213a", x"68854cc622ff7721", x"a89aa8884edc30ee");
            when 30853100 => data <= (x"cc5471490487da2d", x"2216ea41672147fd", x"093bac9fefcbb606", x"a4bb24e052ccdd4b", x"8249d902597ad3ab", x"4cbdefc1c54483be", x"aaff8a71c172ac55", x"9700364abe0b3502");
            when 22890234 => data <= (x"8af8ed5405304ee2", x"094b326dfe6d097a", x"a4aa5936c673348b", x"a9a3c045e04b4bea", x"45e698df56a50518", x"e1d0adb4ecef04e2", x"95cedb4ca6f1a862", x"1adcdaa127cb24cd");
            when 29489883 => data <= (x"44e22e7aca97ac90", x"45ff43bf9510e4d5", x"4b70bbcd52c7814a", x"5c7ba0e2b1c7347e", x"9c95f3eaa0847ad4", x"2c8051d13cce1f2d", x"ad86377256b4098b", x"d7d390d253c583fc");
            when 23974339 => data <= (x"34d52bbe4a09caff", x"ce20665aa33527b9", x"c10f82c2206a260f", x"a38acaeb2abcc449", x"92b1b881410f11de", x"1a1926e27363a204", x"b29c33c51c6dbea7", x"a4683703f83eab0d");
            when 29305681 => data <= (x"8be917cfd46c5ea1", x"1587acfad4a9e0ca", x"5b99e210883e2f37", x"14eb53c8b45cc6e2", x"75f47cfad26a933c", x"7e3e44c86798bdc2", x"44704bae4fe1d8d6", x"7b5bb5da6e9ae813");
            when 30941391 => data <= (x"ecd75991d0a985dd", x"e7fc7803ee1f7a15", x"bd93d1c31dee2aa7", x"f05c847160dcf29a", x"9e6f36627d74b05c", x"aad0cc07ec8e99bc", x"da1d59a8489abfd0", x"06fc2bb6d15c4a62");
            when 8230292 => data <= (x"a6f17dd148837057", x"772df7f4b9333c3c", x"b02cc9441b368996", x"b648e524824b5449", x"ef36c195d649ed69", x"dd3d8f145185a4bb", x"57e5dba11af89d56", x"91ae8c2be2f511f6");
            when 1580187 => data <= (x"acf739d6cdec3c30", x"efbb4ed58b0beefb", x"6d079a34b0c66390", x"a87ede329d0c2106", x"f0e3a074ca37f7a6", x"9f3e7f63bf0b4d87", x"a321c8d5b4060b53", x"e67785f8a0013ee5");
            when 33344696 => data <= (x"2e5bdae48648eb4e", x"51566cc7e41fdf4d", x"4ea169cf4af07d0d", x"cd82aa5888e12097", x"a2a8d6dd2ef09f8a", x"cdce36c3f90eac99", x"f325251bafe56ec3", x"3221986e4d48046f");
            when 12876694 => data <= (x"24b550da38d3b8fd", x"2bd87267175eb845", x"9bd0feb655c613c3", x"eb8fb8a26029e822", x"5c43f06511c8acb6", x"e4eb547f794b14cc", x"b418c304d40ef9ce", x"0ebfa2b1e8f0c836");
            when 27806521 => data <= (x"3f9e97b565afe988", x"faa7b7d9a39875b0", x"3a5290e9907cb7eb", x"cae35a898126ada9", x"a55cd3b8672a47b0", x"083b41f19cca8cbe", x"8dfa4ffcf0e97011", x"8f74c1bc48a93364");
            when 21792499 => data <= (x"256719f4331cfa83", x"a031e2fa45ff7b0e", x"825e938797fdb9a6", x"72e849e2eec16bde", x"39616c7a815293ab", x"73753499e7bf982d", x"d04ac1247b91e370", x"7f07a84b957f9af6");
            when 18717990 => data <= (x"4fdae6cff04c1125", x"22889109573c54ca", x"a9eb538b8983e760", x"69902e90af018960", x"5db4339a382eee42", x"6581479bf68ef90e", x"0f2fc847df3728be", x"67d966d2f6ccb33f");
            when 10457558 => data <= (x"fd926cfaaa34aa22", x"1e089549a9a32430", x"101f8e1a61e1d06c", x"e7c56b518a3bb1e6", x"b49f18855de8df21", x"d2fa294c7a3dff59", x"b1912434930294ba", x"a8470b86643c89e6");
            when 7991422 => data <= (x"5dda0d4130a5461e", x"5c0f788f1509aed6", x"7a6be034ad05cb9e", x"b98d21ef4a856584", x"1a20af39ab1f5469", x"fa467b6098fe9f74", x"30ccdc983bcc97f6", x"24f585cc42e58385");
            when 11411505 => data <= (x"c4043631a921d676", x"8deb03d09e59d9e1", x"8d1037012e101e70", x"e5fe9cf85fc12a44", x"8a81f6d013ad4768", x"d4441244bba3df55", x"62b3a211377d80c1", x"54f6bd50ba1b3967");
            when 20015866 => data <= (x"7b53cad4999eabab", x"1ca9143296122075", x"76f51a5956b18908", x"be6b8597431a492f", x"f7bf9fe2626ffb53", x"b7c8dfe9dca78ba4", x"4fb23dc80e54707d", x"c249dd71c23c5f90");
            when 3974167 => data <= (x"71cdc7015b349044", x"63d41afe426fe325", x"48e82151c996d222", x"6aa3e655b86db633", x"a1bddc866dcd94fd", x"11ba2a8b4f4c9c66", x"7743c99ac6d15a79", x"d6feca410bf882ef");
            when 18203681 => data <= (x"c1fb308c31fa921e", x"038af6adc44b53f0", x"87fb509308ba4c5e", x"a81f940cb8ef4311", x"ac9cb9ba2b934901", x"1c52c82ca6a60d1b", x"68b5673234c33c7c", x"e9cf3759d2f6f21e");
            when 2214292 => data <= (x"f225510001bb2d70", x"00e3dfe07d8fe726", x"4b0f2d27f6dd237e", x"f1d61bf9a664999a", x"8ad6866b4fc3dabc", x"d07f218c6b14a8ac", x"19778704903c17e2", x"6630c70a85efe076");
            when 22761233 => data <= (x"e94dfecbdd7bb65d", x"e55ddce544f55007", x"4f48227cf19809bc", x"1cfd2ed12fc024b6", x"b7fda7dd64617e63", x"4c60a228413071bc", x"0dd4d7b658aae586", x"b063ac85800e7908");
            when 23112762 => data <= (x"ee32c4aeec84b47e", x"72b81339c72389f9", x"51cff445f6430acd", x"6b8d385588e37996", x"34bf5ebb0750ac77", x"96156e075d1a0262", x"1bb2f664195ce25c", x"d13433a590e7c249");
            when 29599038 => data <= (x"83ccf0569428bf0d", x"cc3389e8eeffc83e", x"df03c265a7b99f4f", x"187d1d02116b826d", x"cbb7707a25a5a16a", x"a371ef4c7d49f823", x"77f5d2c45225b751", x"ace2524edf55ad94");
            when 28421901 => data <= (x"c01e5a17533530cd", x"1ec4641aeaff62ec", x"18d21aaf64759360", x"7ef9b09cb6405941", x"342ace028d0fe7b4", x"21bdba6a8d7ea9bc", x"4964fe819fd270f6", x"289f54e89407881d");
            when 33250753 => data <= (x"a8c668bf211b0278", x"a12528e92c195e55", x"feb965b40ad53347", x"68fb4dd31db9198f", x"e73251cbb7a92015", x"2e058c91e5eb7441", x"f45f89d7570520dd", x"5537170bac4a8415");
            when 11700685 => data <= (x"d0a5677b708d39ad", x"e1aebc302c479bf0", x"cd3ca8cdc62033ff", x"0d140f746a0e6676", x"fa7699dbd8dcc45c", x"e3235a27008c552f", x"7ab1502b4a428dc8", x"fbfb567bc78a877c");
            when 5004036 => data <= (x"ad43cbc99a023a5f", x"268bf147e6e15f13", x"215c5d07d8aa6f35", x"df8429dce7dfda2a", x"d53b19c03b508db3", x"16f454c3aa11ef7c", x"ca8cc4c173ba1935", x"1b74a2bac48e0d19");
            when 17608267 => data <= (x"6954d862b65e6bde", x"c2372c91ae29d545", x"01bfe4a7be6d0741", x"c315cfd06b4bbef4", x"e54628e5fb41264a", x"77c8bcf4c0d469e9", x"def06b98ef1ad787", x"21484d954982ca60");
            when 10365569 => data <= (x"4e451ad0e517f499", x"e646ca2e24f43e63", x"d0de301540628783", x"19e45fcf9828dff2", x"e9647ca1727f8806", x"dcf3cd8424290f44", x"521e488477d9a221", x"4c0863a58a9bbab5");
            when 17109301 => data <= (x"5affd17544e250f7", x"c5ee7912c7995fdd", x"7f64bd2d45ae3a3d", x"71ca060b5defbea5", x"a13e0c0eb02b8ab0", x"852624a7ff33027b", x"29098769910b3601", x"c039be452079c96e");
            when 17433370 => data <= (x"c20db4cc53e75df8", x"1facba5ebaf03e11", x"cc8c30a43de143b1", x"231fa6ab06041aeb", x"ef244d7ac4a8c7d7", x"adc66e0808e9cf57", x"54a024a5135dbcf9", x"79da702bc666cda4");
            when 21238213 => data <= (x"df41008c3012a012", x"6fefd56cbc566265", x"6694fedc836d2c19", x"972d3bb12d3df8a8", x"e83f7d58f658b8ac", x"d7f15c4c0aba7ff9", x"edafcc87396dfbb0", x"736c279f3fed41cc");
            when 4897868 => data <= (x"a919238e8acb87a6", x"b631f853e0c82306", x"742a1344652f1122", x"3b2e4f6f3328b0e2", x"4a98e613ff79c450", x"1b8267475894d25f", x"01dc5aa9798eec6e", x"eb75d868be8b82da");
            when 17311609 => data <= (x"0d4c1bff49363fbd", x"55820e139d72f269", x"2c6bbe065832d6e8", x"bcf70258a6c357ab", x"9c0f6c833a982cb3", x"1d8c3e6862fa03d7", x"e6639850a5abd0f3", x"64406d6f961afc46");
            when 7221517 => data <= (x"2bf1f172b14d47fa", x"c46b49aec3753054", x"4a82a5bff94360cd", x"41626d7973e69570", x"6d880ab1ce4782cf", x"94f5e74f7cbd8dcb", x"a133dcfbe500b0a8", x"199a680b9fb7deda");
            when 28127957 => data <= (x"3978aaa2a7328b5b", x"301f9bc94763287d", x"07abf8944cbff780", x"1fc21de517df1976", x"d5b569d85dbf9594", x"cd2c8ca0c587ec50", x"d0e8ae52721614d4", x"c382c74e41b77724");
            when 15627891 => data <= (x"a5ff133a69e6f825", x"e120068a6adb2e5a", x"20a92dad855c217b", x"0194ec6e06b443dd", x"5c6fb0eefcf4156f", x"3f346dc8294a8b52", x"de3b8b01b2166b1e", x"1fe905d499d90998");
            when 13455912 => data <= (x"58ecc0d8716d4c25", x"1c4bdb99fd87911a", x"3763e1a0afe76dc8", x"f30f0bf9c59c2d00", x"b97675fffbedab6c", x"704c8cf661f8cd51", x"e85c0894d1edcdff", x"6b939c098fdcc387");
            when 9827801 => data <= (x"6ebae2e34e7381b7", x"63743d87cf6989d4", x"d06961b16dbd04eb", x"1ce2f340ec6ae4e3", x"0c19bfce1158831a", x"076ebde56aeadb2c", x"c17757e58574e7ae", x"6f67a46ee81d9a30");
            when 9182350 => data <= (x"98b29affcbe1655f", x"48f901924086fa23", x"6e6ef77652b226ed", x"d2bdb75c9ee2e639", x"19283a5f6a14238b", x"7589f389126bdcf0", x"b7dfa8f28adf8462", x"4fd6e2a0f2dc9a9d");
            when 17175856 => data <= (x"cada05a87861815f", x"46a5f07067b375c2", x"d0a3c970e0b121c2", x"59ee1d9f0b45a6f5", x"cba723ac0e7b6ce0", x"26abdf64d56cb709", x"77706b905fc2f0bb", x"5ac4eb37832cdb37");
            when 6505459 => data <= (x"049f25865013c824", x"8b77c9e822788620", x"3c26dac19da7ce88", x"22360538ed09a8be", x"15efd5ad96bf1313", x"7f47957cfeea7240", x"ca7990e33fd764cb", x"e81ded5039ac692e");
            when 26838293 => data <= (x"589db2a342bf8271", x"2763293a4d86bf88", x"eb6546c3bdaea84c", x"198c14af0e0b89c9", x"fbe81591d1ed7d83", x"0f1dc41eef9badb8", x"1a8b4c602eab5463", x"1101bbebd9a22459");
            when 11260915 => data <= (x"0791a030d46a5e8b", x"3cf9369eba6b8681", x"9eb3fe080b3f7ef3", x"2d974952366c43c4", x"348872a6f9e886bb", x"6f7bcdcc2629f59e", x"1010ffcc4d0b18d6", x"63c662853b0a5394");
            when 13216863 => data <= (x"874de0cdf879c833", x"30f6d6ae37a7f0e8", x"713bb0e3285bc5b8", x"6de2482dc7884ee9", x"1bf9a533a1dd1e27", x"bc5cd4d0e7c29b2b", x"4503a93592f54996", x"6d2a6a2936948be7");
            when 5211522 => data <= (x"8955132e644f2d19", x"60068ff12fcca214", x"c9e6145c6214535d", x"ec90660fdd34062e", x"643fb33413247ae3", x"863be9663b05686d", x"079f679f061020d0", x"5892a3ece262f073");
            when 7988861 => data <= (x"4108e95ea37a32f1", x"3d7532c0eb1fc9ef", x"89435d9e19841a34", x"a0fff4e22f14662b", x"375d298ca0725f34", x"effed286f109d79a", x"57b2abfa424f927e", x"106146d788ce3e6c");
            when 27827510 => data <= (x"f327433631c05fae", x"789a9fef0f682322", x"f18a0bb58818900c", x"adb0307c72920207", x"004ee6a706505c70", x"7c9123346c5f0cd2", x"ae4ff3b1881d5178", x"2c7d22db331d360d");
            when 11200591 => data <= (x"c70f030ddeaaf12b", x"8d8c5b2e2a6fb124", x"b542ac28a98adad7", x"7bb4fc2c5e5d5ae1", x"54bd32088f13ce52", x"68cab9601896fe8e", x"40c549d408dee8eb", x"73d515ac711705c3");
            when 9038835 => data <= (x"4410b59fa6d2532e", x"04d9819e372d0e6a", x"0252d1b421a0645f", x"a874ac8d0786d760", x"1f0b51fe887c1444", x"64dfc9a1b0c4a19f", x"e082ca9f3328ed82", x"7800555f8fa91134");
            when 15902038 => data <= (x"a0a7821f9b2170ca", x"a2dec32702251a9c", x"bf0ca193e23e4e30", x"8edc5828f2bc90e7", x"65e59114998a08f3", x"d082d6d81c6f5430", x"f2ef6c48ba7b87ef", x"09365d316c5291c7");
            when 33028293 => data <= (x"46e727b0f97f2c30", x"c1feadaa0c60611f", x"b71a28a2b41f681b", x"616e1f9915aa1db1", x"fa4c502ff8168b84", x"60ebb8970e69b2aa", x"014cfb649f17e342", x"1714dd7b932955c8");
            when 31648827 => data <= (x"63777746e5cac85b", x"3f1f237806bb01c8", x"f6c3deba34bf5ec2", x"85052e96cb4938ce", x"6fbaf99913545692", x"4dd95e4f372de1a5", x"2a86f3b6cbb710de", x"c6081602b7e2d6e0");
            when 17106038 => data <= (x"25b00866f286346c", x"3afb992408432a41", x"a835d79ba5f60bf6", x"eac336ed929d7968", x"ee89870b42a0ae0e", x"bd544e247c19e530", x"47a3534e91b9230d", x"ebccbef2ff76caa6");
            when 1964256 => data <= (x"bf0e08288eadbddc", x"fd5ad291fcbf8680", x"0df43ae9843a45d3", x"a9eb61250e4414a5", x"cd3f17b7812694ac", x"807d9903f48d30c4", x"bab89f03b4590a60", x"597abccfe5cb3cb3");
            when 8668677 => data <= (x"c6fbef65ee8b18ad", x"0d4279413f75994d", x"4213a2cf246bd1ef", x"221f6257b3878d33", x"7cbccaf901819c6b", x"8ea1c9a5c8b2f6f6", x"a2c73e195236358a", x"543544283b64a3b5");
            when 6456409 => data <= (x"9ea5b825dd249c14", x"1e052f3e157f73e9", x"f71d5973631c12c3", x"250404f2fe6d869f", x"bbb6e9cde5fec0bb", x"216db6cde7d01c69", x"ddb46ba3da3d0ff9", x"e906ec54918b218e");
            when 3110646 => data <= (x"1f5c0ace0a566a8a", x"c569d1f9d807a700", x"7b1c12f8af92f82d", x"65d76ee458176b13", x"5a437cf090eef034", x"2f62bb2c3d5a5435", x"0267f29d82ca1452", x"62c2a1c6303d8955");
            when 33669514 => data <= (x"da080d745851d022", x"de2ba1b8ee824386", x"13edcefcf1d6cd68", x"e8db506cdb031740", x"a61e4039f762eeaa", x"1803d0fb419719b1", x"db5b8a98d741aa6d", x"b33be6b3386edc2c");
            when 27447652 => data <= (x"c52265ff3f28ac4d", x"739492a5b8105b83", x"cafd7919868e785d", x"47de7b03a7adeb8a", x"02c3d885f5286486", x"0eddfc01ac1d0365", x"7fa11dc0e7f2567e", x"76588a200353ed47");
            when 32188339 => data <= (x"03e9a54345800a18", x"f661775b456355ab", x"2f2cf244809a1e15", x"ebdcb1dc49f84e9f", x"e77edced1d01fca3", x"184bc2679c4fa57c", x"77d19348ec1ccc33", x"1de386a00a3268e7");
            when 29353962 => data <= (x"f1c89dce2f80781d", x"4b3a7fe7eecb9ce1", x"d1f21223e9f7e430", x"0f252bb390ca6bb5", x"ca29363b81b646c4", x"16323464c6ebae00", x"f52704274bc73095", x"a088ddac3e45c118");
            when 29095690 => data <= (x"afd7ced763435e75", x"e423e0b383c4fa4e", x"92bc37bdd8ca1524", x"d052b8a5e3834e36", x"b3877e520b23c4cd", x"ab4365a56599e2d4", x"c5fa843e046226ab", x"5a6f4e3dad9bff48");
            when 29827645 => data <= (x"c1dded44229cb104", x"5ca9b696fd40309f", x"24289f75fcfb204a", x"2f245dd5f4d866bb", x"b5d6865887743066", x"fe075ed4ab14e3d1", x"6d9c711eecbd1759", x"3a919c6505cdb5d9");
            when 12027031 => data <= (x"5c91d53e36b1b7a5", x"737e3bef4fc44ab3", x"52f6c71c8cd07581", x"2ce4d02609dc0d39", x"291853601fed3d31", x"5b755f27c69a173d", x"f9e30b0f523a1731", x"ac2cecb87e2dcde1");
            when 29803056 => data <= (x"6ba3cec0a0af43f9", x"8a7f62d352433367", x"f39f7589053e644e", x"d145470e13da65be", x"187e71141ca18611", x"67bc8dab39ee616d", x"7c588e11cee7898e", x"d1e5d733011a55c5");
            when 8250474 => data <= (x"e694dea5c920e340", x"27480b8b701794ae", x"dc534ae8e4bce1bf", x"e4a735f23f4bd3d1", x"b842e62661cca309", x"728fc33ce9f22ea9", x"f3c1e4e62bf4bb9e", x"2229815131ff317f");
            when 20363108 => data <= (x"05c46bce66d48271", x"b752e6712f8be699", x"669351b9cc405529", x"8453c411c931b2c4", x"e0f3fd76e0a0506e", x"497d77a2cf2e994d", x"36c7b5ce41721dfb", x"6db27a53625337c2");
            when 5768099 => data <= (x"5d071a8d2bbf0e40", x"0d517a62428a5b66", x"3fca32d86c7ca6d4", x"cf15418d0bc2f8d6", x"8c50dd6e880b27d1", x"28c11dec3eb10c86", x"d9e5db6020e19842", x"924bb4f72ffecc9b");
            when 10383324 => data <= (x"91cdc89050b90bdb", x"1a7426ee6f0cd5bf", x"656a49bad100b6ad", x"0c04f73556de5a9d", x"aa56ccc98404336c", x"dc495d2021acee7a", x"dfec35d0c69b9291", x"5f1e9570330f48ff");
            when 7982281 => data <= (x"534393248f443593", x"5136f8ac4422f15f", x"bd260531275cbad2", x"66e691e7fd3e9494", x"5b28c609f264b204", x"038e79ae4bb7847b", x"2778e64825b61b64", x"0de996640ccb4359");
            when 26224710 => data <= (x"a402ef4ba261ff34", x"917a4ed0e27c98d7", x"ee53b0d04558aed1", x"e85931a72c02b6bb", x"09c8871f34b41033", x"1922c4291f585b1a", x"e7930591f5286440", x"d4fc1a3ab6093d38");
            when 6302232 => data <= (x"96df4063e2fad89f", x"c527ec1bab0405a7", x"c1f7b1b8696ffaf4", x"db74a161835d581b", x"435f940b57af8ec5", x"df4ff9c742a5c95c", x"9e144ecb7bb2dd19", x"99b1d86e9d9475fd");
            when 12602633 => data <= (x"22c9f7a6c464a752", x"35a1832d21dd0904", x"b42a98b12fee24c6", x"ce9fe19d34d6d0f3", x"09a41c9adb342bd2", x"e07f3b6a718de384", x"38d0421751573efc", x"8ca93d5c4deb5ebf");
            when 19977370 => data <= (x"ec67697e3586d0f4", x"69c110055e2ea13a", x"fbdd822f3abae5dc", x"9fe8f475b6335899", x"adecf0bb9808197b", x"ceff9f988a75eef3", x"6dce3ea962f21a25", x"17c8de00eae251a1");
            when 6811069 => data <= (x"b63960be3685980e", x"a5c72b9126c24dc6", x"ee43a6c6f6e11cda", x"91225b419a5a97a6", x"2d7c4b0c5dfd30ff", x"c71d4b2e973db5b1", x"674d66714794021f", x"bf3ef7c02cf53257");
            when 1091994 => data <= (x"a032eb56b0708da7", x"338f23e579d9f172", x"3932f29e2f7eed83", x"d0cbeab81c409f81", x"2896bb38a80b5e2d", x"75fececfe687da2a", x"564a2dfb09cf6f0a", x"fc85442dfaa79acd");
            when 28139469 => data <= (x"561993db1b563e17", x"507c0ca6cd1566dc", x"a70c7aa9b599c7dc", x"3501c4d5965b8233", x"e981031102c742c1", x"64f88c89fb0dae46", x"5d80bb2fc3ea392a", x"91c555190e08c853");
            when 10380853 => data <= (x"fb5d6dbe6c79b9a8", x"3a8b514425b4cf45", x"191c8c11bf7c1fc6", x"d6cec7483bb756c4", x"fd753b438d545aba", x"9ad630a5c41f1d75", x"99b8c02bc82d2491", x"08549ecd453e91e2");
            when 31493972 => data <= (x"6e8cd3bb1546824a", x"30fdbe47ee086a79", x"12d2520c6feb7560", x"d19ce8486111d4c8", x"35ea3904962a8d4d", x"105b1e18ba0dd93f", x"dece5942eb36516d", x"9dd256d15c6a59fd");
            when 8692408 => data <= (x"3207156893435a8f", x"e8527ec480976441", x"cce7e208c50b101f", x"96f4a8bd55fbd77e", x"cb1013ab904df3b7", x"ad976a754cad8c85", x"fb274f4e423e0bbf", x"e53c7a4474d76961");
            when 8233287 => data <= (x"163b39fced360feb", x"9407bd8339d28c40", x"98aa71ca0cc4bf5b", x"1cd6efae311bf25e", x"1706959752df0df3", x"4e8ba84a406b37ea", x"c74521aaa0ad376c", x"2b375ed074f1a212");
            when 26945922 => data <= (x"4c4d7fd705b3c8df", x"bf2c8dbcc257f7c8", x"bd3ab85a769c31eb", x"ace24dde8707b128", x"d201d22384280678", x"b0a46f7db82d742a", x"e89dc66f67b53b4c", x"44012c47f802da93");
            when 27035495 => data <= (x"211186d3824c597c", x"5f9ddc60969c1aa0", x"cfe284b5c5fc168e", x"3fe888d92b8d7875", x"917174b289b71e88", x"3247d9bad3707046", x"ae0a387c4c77d75b", x"ed56f5942c5de18d");
            when 14942174 => data <= (x"2ceec82a2289fda7", x"d9965fcef48f2ced", x"ad4256c1b4b3edb3", x"320d2f7b7272cc11", x"29d931b2f1228549", x"a6ecb6c5289cc30b", x"bbea858118ff96a0", x"9eb314ec36614973");
            when 33842587 => data <= (x"86a060e54a80336e", x"da5f40d16accfd9e", x"d96c68bd76ce909c", x"fe6620e9fd7dfc2c", x"0c7352f26f384804", x"52020bd9a3ad30ce", x"65773441f73fa2d6", x"e99ab1471969afc7");
            when 18120636 => data <= (x"216797ab810b8529", x"5d14e4688ffcfd85", x"823839eb20bae5e4", x"64771fb3f0a3b75e", x"ed3a21e70c44c361", x"2805c6014d2773f1", x"69480b0d392271c9", x"b4b0d77293e087e2");
            when 21687987 => data <= (x"ef7ea4a304dbc91e", x"10c0d54abf3b889d", x"f4d8fc479c5c2c02", x"aa5b041c869520cb", x"ee60d365ce9b934e", x"ec385524f9c70263", x"2c74d0cb9d995b02", x"236bb42dad0aecff");
            when 21334380 => data <= (x"05237d0fc36e6517", x"6c86751d26a8452a", x"5cd7691815516d38", x"e7ea226939afb771", x"03c5ffbe0d5861b3", x"7f8ec60954efc666", x"70653a625003d2ac", x"70aa37bb27c7b1af");
            when 17055584 => data <= (x"46ce94ce1cc057b6", x"b0b28b832f49b682", x"bd869e19133ae18f", x"e45229f4ba4b6ff3", x"e231d484d5f70ba8", x"3e82549d5ad7800d", x"c9af8382073da1df", x"4ea6d47968b9b6d1");
            when 30699934 => data <= (x"5d05cb8f2d8ccf6a", x"e444c27be2e44e30", x"d5d7a25b82ff2f9f", x"03d784a10c3bb2fa", x"70458fa2cf21b7bd", x"fe695a6ba4904ef1", x"06819d54f3953ade", x"78860baa7602140f");
            when 22720957 => data <= (x"c2b0c07762130e1d", x"a57e34497c5477e3", x"3be340859bf69c2b", x"30966e710c431d83", x"c3180306bd3eb3c5", x"2cf4b2142bb57a23", x"5a3944da16d3b0f6", x"9c6279f8b1e2d86e");
            when 6806884 => data <= (x"3e1d713fa2a0a58d", x"eb01dbd65d0722d3", x"4768bc60f813bfa1", x"6b7e2b24977a252e", x"ec2bac7c2aef28fa", x"2f808b88ed120e72", x"7f24f46b07ed1df5", x"c18ae6ab510b16bb");
            when 23855428 => data <= (x"32dcfeb46ac1126b", x"efb86d0b6d3f5a3a", x"549815c233aff47a", x"26a4856c862b7957", x"cd2c6bc7a507f0e0", x"4055f096a11b4e97", x"9765e4ad80b8450e", x"2f92554137bc737c");
            when 27290014 => data <= (x"cec79e1524d13401", x"123d8c381c1fa421", x"3365d28469e3bc75", x"7f795af922fe8b8d", x"356a0a1412bf620c", x"a48f936f077e4415", x"c5f18bf0ed3e421c", x"e0b4260a518a791a");
            when 28179373 => data <= (x"9e73002858fb788c", x"9bdfecddfb03b13b", x"cb93a968f3b0a69d", x"0414dd1c6fcde08d", x"2f1e05c1f944bbe1", x"ed85c71f712ade31", x"33ea272f62d4053b", x"715efebb4a216a2a");
            when 10802121 => data <= (x"22ad9ea972b505ce", x"f0accaf7b361dc06", x"42af91e38de6d8bf", x"480eb5bb5213ec7c", x"87223b32758affee", x"f719d917cad22167", x"09e51622524e8546", x"ec86310b36a894a6");
            when 30077342 => data <= (x"dc86222019b9ed70", x"4f595af61552c90c", x"cbbc268cd443200b", x"e4b1a74e7a8c440b", x"94ee600f04859dba", x"21e22f8e413b2e45", x"41a50f21bf0700e7", x"992331dcd353a71b");
            when 27460502 => data <= (x"e0025dbdf3206f18", x"9e62e1024da9d717", x"12fea1168c674a55", x"67a0297dd3c0cae1", x"7697e3f548f8f345", x"2c549041a3a2a969", x"2332d7d90b50960e", x"18dc55ed53711cb1");
            when 7430648 => data <= (x"7a91bd54d2f7a658", x"1472736dd1a8560c", x"2d8c73d604210bb1", x"44a8a3d2d0d08c76", x"62c3f163147c5464", x"b655148e3f5a28a8", x"513a3592a42a6d13", x"d2df27a9cf11fa85");
            when 10624456 => data <= (x"772d64bb07c9b4b6", x"1853a70bfc04c273", x"65db800006faf300", x"7ccf2cd6d3fa0d76", x"5aa50aeb2510370e", x"3070c2facb88bd34", x"bd777ef387a9e4d1", x"f9442fe111b00c3c");
            when 23279025 => data <= (x"0c3bffc79a64fd0d", x"df35cf31f819cfdc", x"90931380167b6647", x"ed6efc665f064b0b", x"7e150267a599e477", x"4916ea0c776a9306", x"6bca87b6b590770d", x"86d852b3443acba1");
            when 27524468 => data <= (x"02d8cafb7c501450", x"66dbdd2b03cb128e", x"0f1175dfd8af8f02", x"521861c28029874d", x"6bd66c4996ccf54f", x"889a4e904bac5a3d", x"9692a78f91fa9371", x"ebaf36545a86eda2");
            when 32796405 => data <= (x"2170b714fa80d443", x"949c6c75345f8470", x"a2d295e24d81f1d7", x"ce3c6ae120f3af26", x"81a1996975cae3d3", x"ae54fa176a346633", x"a9de546faae53e32", x"b7e3eb83182915c6");
            when 22259667 => data <= (x"ee8884b0d9df53a2", x"3645496f549f88bd", x"eed56e062af0ca8d", x"34cb58d720a3bbc3", x"e09df28874e43bd6", x"32be04dd42a0b8d6", x"8822ef719d0d25c4", x"274975964e8888e5");
            when 23605185 => data <= (x"e47b3cbc9376c41e", x"8f95c4657b1cdc49", x"ecc1296dc869700e", x"3109feee015819d8", x"da71f984223434a5", x"7afde9d8ccf20a78", x"5fe997a8087b41f3", x"4536ca57f796fc81");
            when 1913676 => data <= (x"96ebda8f6e860fe6", x"4c1569ccdb0df9dd", x"246b3cc837bc179e", x"e4a1c60e757d6922", x"7bad2f7db69041bd", x"138496983fcb8920", x"b6453681e8b14d46", x"b801c18b2c88dffd");
            when 15005827 => data <= (x"bd37c18e754fd7e1", x"e5342219aac4edd1", x"27c389e0f360706e", x"2006162f8d4f2f22", x"3da4412f60b4a707", x"10cc5f5b6513c43a", x"2ba93c29a1653add", x"bfcf59cf40d9d8c1");
            when 14476418 => data <= (x"d37a5d10b2e4b7d4", x"065e55355366639c", x"b02bfbd3d72d00a1", x"76a33b1b3e1875f1", x"637fc80b41fb977a", x"279d062c2ffed5e8", x"ec5dbd8e525d03bb", x"c873569d22d67e7d");
            when 5879584 => data <= (x"8b51c3a50a2deaab", x"50da5ef31caa6223", x"880e593cb106bcc9", x"724bbe0f47664cf4", x"f8e876f17ead8e67", x"4cdbda2f67bbd3e2", x"658be1055bfad70a", x"d9c5cf5ed1011d28");
            when 1197177 => data <= (x"f0e021582abc6928", x"8e64ff1556a311c8", x"9c0236fb006093e3", x"f8eb98296e4e4514", x"8bdea7ec0a78f345", x"e26d95bfacb61233", x"84a4b2b8890d5784", x"2e41f3e686da92d3");
            when 17565791 => data <= (x"6412a33d5610dfe3", x"c55952dbb532fbfd", x"2e7b742750002013", x"120898149fa374d2", x"bf591587b69e8662", x"198108992b809bab", x"9ae4304f785ec92c", x"f69b9e608d71394f");
            when 15768654 => data <= (x"d8e110a127705fbf", x"0ab0c4d4d821432c", x"c7c78ad0b6172934", x"9e65b2bdf75377fe", x"a7d0ee2dd88866da", x"319fa26c13ea9e7a", x"719bcc514000ee87", x"f206336b53e4ceb8");
            when 21043743 => data <= (x"d4588c8cd8e94033", x"12720113a572af4f", x"458ae3cca6c27c0c", x"6cdc170f0d2403a6", x"08e0d9fa6e9082f0", x"5a2e251b891852b2", x"37d007f400240c45", x"cb8ab8bed9cb85c1");
            when 18120937 => data <= (x"3593e1ed72172a59", x"fa9825d0fcf1a811", x"c330425662361afe", x"d0274fe39efe14bd", x"c1651f26cdf1c22b", x"3aafef2847e56ad5", x"90468ef947ba230f", x"96d675298f805569");
            when 20391807 => data <= (x"90cdad0560e1e2ab", x"2afe2be4a818af7a", x"a80cdaf3012421b5", x"db04438e1bc446b9", x"8c72c0f8be9549cc", x"a32e52f6b0ff0aa3", x"56d331dac378a71c", x"9d0b0bbb15a4469a");
            when 31950887 => data <= (x"f03a0cb4992c1027", x"e75aebc9b8020c8c", x"5e8fa35fdc3bc025", x"8195e858db04e03f", x"797722d10685e542", x"7ed2503b58f1fa14", x"fd2a7022a85785ff", x"a35df67d853eefe3");
            when 33459001 => data <= (x"c11928e29fb19f4a", x"869ed0053ee25a60", x"07f5bfd21179abeb", x"927b6f8bf99932f6", x"e9c8e0f17da31e8f", x"081790330eea004b", x"a7a76f7d4f7c5e34", x"953a6dc53e661598");
            when 14012510 => data <= (x"1edde1b1096180cc", x"fe20792bd815ed5a", x"b403c94078ea94b0", x"dd931b0a2bdae581", x"b1d7590a9a21bf71", x"a30de23511be4788", x"201324b3acc9b88a", x"2d6a47d1c27499a7");
            when 31558765 => data <= (x"9a75bec3f58bcfd2", x"8f0bbd7fb0840916", x"365b7fb9f205c27c", x"7e71e15fbb51b400", x"fd5d88cc36442145", x"c8158c1dee42a8fb", x"58deec2ed156cbcb", x"45bb57847f502cc4");
            when 18026440 => data <= (x"a37f2decac27ba93", x"cd72282e86cf22e2", x"96e500776846a46b", x"a6ec4389136926f6", x"d1f6a8724d947cdc", x"5eea5ebb42d5bf8d", x"05fdb86222b06370", x"13b9ffcedea6820f");
            when 3302876 => data <= (x"0516c8906b4c3ada", x"99287cd8a6fd870e", x"62e0c7148863f351", x"5ae0360c07f38a8a", x"139b0b360ff33e2b", x"e0fb3164c23248c2", x"810251bfa61b5556", x"fa58882dd368dce3");
            when 21614701 => data <= (x"aa20b7abd7a3357a", x"91e93f86958bb976", x"da3cf3cfe856d35c", x"03c5005fcf7ac446", x"8aef9302abb24eac", x"9ee27558b2d33f24", x"a65d537b49dc6ac8", x"2df7a3669e3865cb");
            when 18363868 => data <= (x"25f6707cdde9722c", x"3974f95eb625001b", x"98321fff4e0c7d45", x"18d6891b5cf50c7e", x"2625e292adeb0c67", x"8a535d17a9ef8d91", x"80b37a0b667792bf", x"03804feeeccebbd5");
            when 8093135 => data <= (x"b9c23b170bc3cb0a", x"65fba38ba639b92d", x"fbca56eb4c50dee7", x"1f324196b7786410", x"6ed897d90f666492", x"2ed2a95c7bf3f483", x"9802b7d9a418a168", x"22e34d65dc9db9b5");
            when 24457168 => data <= (x"7ea64aa855cefe6c", x"14ae3f6049efe310", x"747930e4124065f4", x"5aab1b959d8a1ff6", x"2f5a445c4aab599e", x"d11a30e717dd0425", x"79b8d213ba87d53d", x"6a2f70450c8a7937");
            when 28106105 => data <= (x"3c59c13d041f024e", x"c16d536058758bca", x"c4bd90e801baceb2", x"30bfb7c3265aa8ee", x"5336bb7b38ce01d2", x"8d72234cbe3a702a", x"80afe7a29d2ff3e7", x"f4fb86b9e57c04a5");
            when 23829273 => data <= (x"4729564cd034b068", x"5552f473716d094d", x"50bb98c60eceea23", x"d5f0077c34362d97", x"02e7e7e5724191cd", x"77a75443bf552710", x"0a3dbf1e93c9fddc", x"1b99a3f9c346bdde");
            when 26206171 => data <= (x"a8481a6f12d91f4c", x"de2fe2be097ef9cc", x"f883e3389c00a078", x"7593a31742e61d5c", x"4583af6f43148044", x"22aad6a29eb76c94", x"9f7595155d10ca83", x"aafb2eab308c0687");
            when 29108479 => data <= (x"16afe94f0ced3292", x"0188ded2b6dcd24f", x"c7eb74021e5f070e", x"96919ef73f37497a", x"768a37ba15af67d1", x"b409062d72b45d5e", x"b307b4e613f45a64", x"78b53634e2649a12");
            when 20583661 => data <= (x"ad38c036fe993f4f", x"71d383e91e4c1cc1", x"1e4ef98b63b3bff0", x"a0d9151e3c197641", x"cd65474ae6e675d8", x"8c460ddffa650938", x"fb51690c43017207", x"20ecdb19f29e0bfc");
            when 32594464 => data <= (x"fbada3500cec7ebf", x"c2655f2454bb6ea8", x"c75ea33fc4b4440c", x"bbf5938b183db9ab", x"4c7bcf2409bdd9e1", x"fc785f4aee0c482f", x"4f1202c96ec4b978", x"4acecfb6dc00c404");
            when 33575945 => data <= (x"aa0aed9729c1e265", x"e41dea1f6a545481", x"576d86bd88c1fe7f", x"6dd802be60717ce8", x"a65702c871dc1e8e", x"97604c1d8e145a94", x"fe39ccace2f1882d", x"3753af1f045c0503");
            when 22347259 => data <= (x"66974490c630796f", x"c9a1df785d36ba32", x"5ea5c113be52f13a", x"b0807086a9070a5d", x"3719eb2b96945433", x"1f5f7706a6447ab9", x"50c7b56bc3d13f81", x"a7118fb328e1b5dd");
            when 29514437 => data <= (x"993aa8d74f0eaea6", x"c122c80c4d931aa4", x"62f62cefc7966084", x"0d6b932403ddb020", x"a90737b4de27221c", x"fde44f84861d1b9e", x"8281ea12aed3f45a", x"8808725d1c94c80d");
            when 13663119 => data <= (x"79b3736ad1ee7d2a", x"f452e29e05b5e2ee", x"4b2472f31969824f", x"f663022841f68b51", x"7867af66bda83976", x"2aa49222d062aa6f", x"94d00d9e3e42aae2", x"83e38b1b50ce7363");
            when 20056798 => data <= (x"3fd6920501f029b4", x"b317fee44564ded8", x"15cde291d16c58f4", x"a82cd135839f3326", x"2a2056771b308c41", x"4971e72b3d87232b", x"1cdcacdf6c831520", x"542f7791356e8941");
            when 31670306 => data <= (x"83b01682c557fc8e", x"bd58b3be141cb253", x"d4dfb92cac0fd7b8", x"c23f4784e0010f24", x"ae7ea1bac80ca876", x"af2c3c35f1d8d550", x"e4cbf50ffdffa230", x"7eaad7351683573a");
            when 32828189 => data <= (x"4d4794099eafdb5d", x"b26053f29baa70ff", x"b1c3195afc279652", x"62c4b9fb58f6ad6e", x"faa8b7a933a3c391", x"fa32fa7b94db4d29", x"efb5385e13191ff0", x"e87879b9ad1eb792");
            when 30095037 => data <= (x"5b66858ef57acb96", x"4b425b90accc16c0", x"82206392b4e19051", x"1f9324759ce6303d", x"cdbe8de4c03eee5c", x"b96d7682b66af97a", x"def7d2c703a84817", x"88527e0319cc8d55");
            when 7425204 => data <= (x"1ed0f49ffd3ae9fa", x"60b953d493e54a6b", x"2235082743933ede", x"4253d09058409a0a", x"02348078fea93436", x"887247706c982829", x"3ce5d93c3ed11911", x"c772c057c52e695a");
            when 13131189 => data <= (x"8a05760591648541", x"bf84c86df71a1bba", x"ea061344a2e08aaa", x"b6f6fa1f2ba8c6a9", x"f0af0ebed8b64cdd", x"faa67d55648528f6", x"16941bb654a4f700", x"fe68a2a0a1b06229");
            when 21869338 => data <= (x"dbe8559e93723023", x"2cd7f87dfd598375", x"a5720317e5616d21", x"e38ac86c308f6dce", x"95ea0e34e3dcf82d", x"620425779765ea7c", x"2fffe687c5523f1b", x"6cb521f09a1b1f95");
            when 25946009 => data <= (x"32066044c1c5373d", x"b2065d91d33b9798", x"b7e25f19eea5c94e", x"6cb5bc5ae87f6652", x"02bfa3c393f6b40e", x"fef12cdf32265e96", x"70ea1df4baf28319", x"1ea6a3fe619c3cba");
            when 5952280 => data <= (x"eb3c3f8bd789a38a", x"ac7db7ccaa5fed8d", x"b8bc746a9d60c815", x"f858d2ac6051e045", x"a8a997cb1f6273c0", x"af5102abbadd92a9", x"6b295a399177bd31", x"97da054eaf30e33d");
            when 6880823 => data <= (x"29ee2f974743b8ea", x"877ff34fd812611a", x"44e3700b7e6f9dec", x"51bd15cefbe1f136", x"e5254feaebcf5bfa", x"4e2bf8e2752c65e8", x"182b15f5b556ddf1", x"fd9f88a6c18e9355");
            when 33815075 => data <= (x"4b3f0476860bb0c7", x"406610fdbc999983", x"82f2d5c5a0aa36d8", x"4a5dd3a605631948", x"84ef0a31d43accff", x"990eea641aee3734", x"b5949c1548a479dc", x"ed72f93fd2ee7709");
            when 15666906 => data <= (x"d885d615ecef0d2d", x"0e9c224f6397bd6e", x"d281a866b3997dc3", x"ced951117a4734b3", x"19f78271d822742c", x"3312cedcf0b94c53", x"420f6c11a5ac4272", x"cfb5093939bfda95");
            when 27346086 => data <= (x"d5feda90f53e5dda", x"370cb69c7ee5177c", x"caa0a13066838ef3", x"c6b96fa6bcc5a737", x"c7822145da972911", x"0b1e9322ece1eae4", x"e896a124b6ff09f1", x"900991be85a0e978");
            when 24771838 => data <= (x"0e2afc49385b7773", x"f3e9a5e19b424b34", x"2a05bfb3fa9e69bc", x"43ac0ae7d2c12876", x"fadf31d2bc534d8d", x"2651e6615dab69fe", x"3e39aa5e3755355a", x"e5b0dcb42735edec");
            when 13110672 => data <= (x"d9e202ca50079b5b", x"d15126333999fa5e", x"00f2c80f4eccd4e3", x"d61c2544f527329b", x"b2614d8e78907e61", x"97783b66c7cf4059", x"dea0c7f06ef315f1", x"60985f593483ba11");
            when 2052100 => data <= (x"52330057f7c86ab3", x"5240cf3d08ad6576", x"2971df3ea8babd53", x"fa7ae469e2b0c0d9", x"e43a198042128682", x"ccf4025c7103b044", x"a9701c2dcba34be3", x"2cc088138ccc7956");
            when 32574421 => data <= (x"7043ca9af83bb05f", x"80addf332bb0f090", x"5753ac481c22a2ec", x"e977636369061311", x"7af9db07a4e771fb", x"74f9449426e1eb3e", x"aed6b3c797a8eb12", x"d5a5f4237baa3ab4");
            when 31234921 => data <= (x"a3b4c963d52a2f20", x"504473ce7c12d4bb", x"60eda0ed454a5b25", x"5b3566132ed2b181", x"aff44d1c4312f20d", x"0624e49e1cd3e499", x"7c111c645348ff46", x"28d4a208c7d76208");
            when 32592171 => data <= (x"180d5eaa477efc50", x"bf44d0b2afc52c0e", x"a591f48514d7a0dc", x"1c1d778ac9419c59", x"632155f989027d91", x"9bf9eddccad9e7b9", x"4ef9d042548870aa", x"3860303520a40692");
            when 17571725 => data <= (x"2214db3b44fbe4dd", x"9023c880685dfb33", x"6afe4cdcbf4c43b8", x"9bfba8c28323385a", x"089609b151e82006", x"729457102758f82e", x"eadaa2c7c41c9223", x"9802c4c44c0279fd");
            when 8792920 => data <= (x"3d91abc70a661e2e", x"a1fc4c3631acc021", x"e0528b30a10fd667", x"d3b5d9a7abfb6d3b", x"0fb5ff338859112e", x"dce8ac4cea637eae", x"598b9b04e6c81492", x"fca3de2ade69579e");
            when 15575243 => data <= (x"a8024ead68a4b235", x"ab4ff040d258905a", x"2cfb494c430a077d", x"02c92f93e14484ee", x"30822b11e8431394", x"207009163ae47066", x"269b36c9d36d6d1a", x"8decf52919c2d8a8");
            when 3799157 => data <= (x"65c808d26159a1b3", x"9fdec580f5f90802", x"0653a5a9443d24d7", x"c04ffe9f2d0071ba", x"7202923392b674d5", x"f3e657702c126f9d", x"9ba62ba0373419ad", x"9fadae0e5b110d62");
            when 2641937 => data <= (x"5be500117e9560fb", x"1a0da397e04bf796", x"e0711812c1fde1c4", x"1a6ecde8c494cf49", x"4930fa091a11e06a", x"89f8d52a8d7b6ca0", x"2145bbed5f2e2ee0", x"fe2dc4d6972a8c11");
            when 16771274 => data <= (x"69e98086d889c58b", x"f5c901d801cf731d", x"c484f506764d1034", x"9553e070c4dfd1e0", x"c4a10b9d8d64ea7b", x"0ce7a9749d2d6e90", x"42d174ed8d3903ae", x"ec8946c162c0c736");
            when 25482256 => data <= (x"ec4a41e7b465f7b4", x"44258b70b4effbc1", x"34c9bb749adabf3b", x"c44deea88cceaf08", x"5d8b41f6ba62bbb1", x"6d6694cfa1880b3a", x"b72548f37c1fed99", x"3bfe979c69bf36be");
            when 30622587 => data <= (x"865d8c6769c77d0b", x"a514092d6ff88314", x"7f5803340cd59213", x"1517167d87a4fb90", x"ea65969c3faf0318", x"9a091ca8d170eab5", x"26812a08df5b1acd", x"55f7797bf918dbab");
            when 22408643 => data <= (x"6ce376ebb872c50e", x"f27397a4862deae5", x"2453d44bd17d185a", x"ba380d025aec614d", x"71caf4f3efdeb13c", x"e9c9e5083197c066", x"408ca0551f0b9d33", x"937a52f544d665df");
            when 12042307 => data <= (x"1ce7124aaafbf56a", x"67317c6db0004abb", x"10cdde5355f3ae00", x"6ed520ce3281e683", x"f6795ace3a9a9459", x"3e73c30d80541764", x"a76e07561ab8d5a5", x"d3cc8580ac4a17f9");
            when 13635576 => data <= (x"ff517fd2f5fef9ea", x"64bde2cb70c4a949", x"60b765f1ed65816b", x"7fbb2a2964a77f84", x"70ae3a598b1d473e", x"dd8135d224850d80", x"1567f32742cb5cce", x"0d5f91a37376f5e8");
            when 33415296 => data <= (x"78a891441728784e", x"03158f11627b10c7", x"af7567cec9f8d0ff", x"2d096554ffe96140", x"1796692cd5bfaff3", x"e3aca2c49c9b5a7a", x"1aa502cb15a55152", x"f8b2d2b8945a1428");
            when 15043753 => data <= (x"245f5c798f99cbd0", x"2797a74cbb0a3548", x"9b0b06d2c8887dec", x"8fd530a0f9a0531f", x"72ab73b1a45fcda7", x"060184d3c8b0ab1c", x"34c577986bb63ca5", x"9192952491f29a16");
            when 19316714 => data <= (x"aef1f8cd8784161e", x"c63d85b30592342a", x"fa95e6ecf152a64e", x"28c2900bca2d3003", x"a495eb94260e644c", x"0af9378a0832f79a", x"7ec99c7a17e33131", x"808c6bc1a32db505");
            when 27255371 => data <= (x"9d33c4ceb9359497", x"9ac5724f1eff7e5a", x"8c861a4a14b4ccd8", x"afcc3121104aa2c8", x"db2a6be5c6e9a402", x"4d2878f03b482f95", x"efe66c8c90f4f4f4", x"c90833edf6875666");
            when 15479944 => data <= (x"b03ad1f4eb874c76", x"9c9730fad5da5c42", x"1de8ad19623c1496", x"1fae668d3d04f2c8", x"a0ebe19304beba72", x"24bc9e4fb889396b", x"7e36f6bf7a4db079", x"625bfaeb61897312");
            when 18178509 => data <= (x"239fcd43ccc2085d", x"ef934e2ab4970454", x"93acd2956adfb6cf", x"601b6bac7a997735", x"df805dff0772304a", x"da79e51b97c396e1", x"61db6a68755f8f42", x"d4d811d64e2a53b9");
            when 1420207 => data <= (x"b4558e5eae5a54c4", x"6d3ad5072f8555a8", x"5d25d542cd3200f7", x"4bb1754a1f70bc8b", x"971060d34a1470c2", x"c36bf019b3857dc6", x"dea674de83177d81", x"f56aee347d71e77b");
            when 15767183 => data <= (x"76e6fa0e890b4ee2", x"225848731e87a70d", x"a936de7e03b50b9c", x"78a2febfa88c43a4", x"9b5b976bbbacae53", x"29ba04033a92d6cd", x"ad5d0566bc6407b5", x"22e651cfb46e0029");
            when 19277129 => data <= (x"94a625e25a8e29ff", x"c5563de3aca83986", x"5d031b828004be4f", x"2f13b3e9d1e3352d", x"e67c4b455b791a35", x"28f0a3b2b075faa9", x"8d1525919cb8dcfd", x"3287256f88733f42");
            when 25714898 => data <= (x"01907fd85d06250f", x"1bc1e16cde418fde", x"9d4d98eea9580090", x"1cb2ebd9d3c4bc94", x"9d25ad9851d11f02", x"625d2fca111d96ce", x"76890173409cc843", x"40fc8795d8bd78c5");
            when 14918289 => data <= (x"4436879c1e660e87", x"6edc0419b3c352c5", x"aada83eff1e3cffc", x"5c60e8dc4f8159e0", x"75f4e19181a97281", x"b0dea3de89519b8c", x"9bdba513c6e2b979", x"c1ac7667dc8fab0a");
            when 18083492 => data <= (x"ce273ba03cbf2a61", x"e56abf612e03dbba", x"032be389ed520258", x"e71f57ef8dde04ff", x"4714818a9516a3cd", x"4a3896bddf83f0fc", x"687a767e87d2ac91", x"944a5a3cb9f79062");
            when 16625019 => data <= (x"6f8e9a63a97fe8d5", x"85e79257ac14ad5a", x"6ba16b635ae59238", x"06b94bc527ac10aa", x"ab0d98bfead7de94", x"beec315a662fa982", x"040f1d8f39081405", x"68eec2682bcea245");
            when 28893781 => data <= (x"09b40033bcd2ac51", x"e7e575afcf1517a2", x"72ce439c17d19697", x"195aecfce7add4bb", x"3491d21b8d7f8ac4", x"ff922b3d318ff8de", x"6aa5762a743a8bc6", x"f55809cb6ee94dd7");
            when 33531381 => data <= (x"4079e6449481059f", x"864c83fc09999833", x"3a9cb3d04f54e931", x"aa7346705cc9b15b", x"6fc191c6e37de822", x"dcd8ee70fb7c3166", x"0fc7081b0f4f4654", x"89b5d7eaadad9c03");
            when 13194685 => data <= (x"486357ed5d936c5d", x"d744d2e4f7c47a35", x"ade951d63311f717", x"1930c28fbe40470b", x"fcde7ae889e7a3b6", x"92516c5c43c96921", x"3e228141050560e4", x"ca1a56d3002c20a7");
            when 11310019 => data <= (x"ff3f505d7bd75a3d", x"beba9c431ad92d9b", x"9ffda048237da6e7", x"ebd05ce531ce87d6", x"26977e89574d9405", x"df6c8c2e82cd5ed8", x"dba2b0a1639589df", x"bc49a1402a1f5bd8");
            when 723981 => data <= (x"cc683fd799c9c71d", x"e85ca443d6a60f13", x"0c415b4fb76b94d5", x"b7513aaf72d3c8c1", x"693cf5cc3a1d92d3", x"b61837af4f93b7d1", x"4d674b582a05dfe9", x"f288b9fb5a4b4f0d");
            when 24394593 => data <= (x"b7b4395627609cb1", x"b23292bacbabc638", x"725004669e9a4445", x"ad1bac07b9da5a53", x"dc5095de8b8e4cb1", x"607a196e65711a48", x"7a18d7a44ff78936", x"2776380968f7e8de");
            when 24326958 => data <= (x"12521c3b75d9563c", x"311302ab31d041e7", x"24d3d26a5580d990", x"c4e7e91e7817730d", x"aea70023b34ce366", x"e8fc01c121ed5219", x"59e90a27c68cd24a", x"62ad6b21f9726e83");
            when 8544035 => data <= (x"352294ddcb3942df", x"fcad50c115765066", x"52f41ec0ae4fbf3c", x"4f25458051a6d9de", x"9c78382140540766", x"76cd636641cdd76c", x"cbaa870a6b41878c", x"b9069222e9f2856c");
            when 33834845 => data <= (x"9e4722e521a07f2a", x"146a6e2e70dc3105", x"e9f20048912e3a18", x"a503f1424c3b0dbb", x"b72190fb6b8aea02", x"bcb2543b1f73d704", x"fce268a0b9b2e8c8", x"a847145ea1418f98");
            when 7559611 => data <= (x"15a397ebdfeba869", x"d8c3c44d222bb109", x"ce135a0143d78754", x"f1bd717761390662", x"cb509f5feabf16d6", x"62e2740a3fcce950", x"83c72a8a9c0cd690", x"dce2f6dcbc321dc2");
            when 741007 => data <= (x"a9950b7324688243", x"8573bcb438f6becb", x"77a5e6bd6013a611", x"3ddc25834c225935", x"0c9b298e45b5d228", x"3eb26e15ff0b8b9c", x"610afe7cac643b0a", x"e9cd01d33f5795ed");
            when 11227845 => data <= (x"2e09f95d5b0a4e0b", x"5fa3dc5ed75ccde3", x"19f4330615e61b03", x"93719911bae18465", x"78b16d15b730c4a3", x"1018dde9ab9c20c5", x"82edc79cf370bc3e", x"a8c84330c60cc32b");
            when 8078402 => data <= (x"acb14646681dc15c", x"ebb431485fad94e2", x"0a8e7a765fe19804", x"77bbe48b8dd78de9", x"4faa3fae03e1e52f", x"99880ec42cd2ddcb", x"b52b392965abddef", x"24494e170463e42e");
            when 6538979 => data <= (x"b02ac83166b2bd41", x"7e8dc4c1f93c172a", x"6345e8b83dc9df81", x"8039a93b7eca2d30", x"6fbbb40c05e6ed8f", x"086db014410119c5", x"7166ee57ef1e8b6e", x"b2fee17e05b9d72d");
            when 26863818 => data <= (x"7429d593a5bf44a1", x"74fe310794408759", x"1748680defd30344", x"71a127b6a4744079", x"2dbcf953051aa936", x"1aec11c5e8c05241", x"9e262fdfa5a79f8c", x"86dc9c9a0d718910");
            when 1214807 => data <= (x"0db7e7bbeb94a96f", x"5b865a95cc41b858", x"ea54de80f8670fb1", x"c17383a80b441693", x"68542053b385ad54", x"b7bedda612cb741c", x"0d82af8c2c48bd29", x"55f302dd0b019368");
            when 14528404 => data <= (x"0e0b2cb19382ee0f", x"1f6bfb21a97aae18", x"3fe7a66812ba8198", x"d0167ec6fafec1f0", x"24d86338c6f8f486", x"7a5dca746d462d09", x"8a735e7a39767113", x"56b3ddfb585b5991");
            when 9946341 => data <= (x"1b96c36fd76ad991", x"dac71e6fe70476bc", x"542d1def53795c23", x"b1f50a8e0de100cf", x"3b2181f8f80ee61f", x"e3961f7133a43a71", x"e36a490e40a3b654", x"f76d498ed910ab54");
            when 1360345 => data <= (x"16ef9cb3f44d2808", x"08b6bf27821efab8", x"47b424d1613ec5cd", x"1ee8adaeb01918b8", x"7216a8aa3681c7c5", x"c29ae50cb3347f3e", x"28738e00f252621e", x"1fdbfb8e973cb76e");
            when 4140641 => data <= (x"1881d2e730d72180", x"90b4463181ea446c", x"866ee65520fc9ec8", x"cff7c4a3902c4d84", x"b576a154fdf990b7", x"835681c97e5ddcbe", x"55c14cd63845ab42", x"6e16494cc4128716");
            when 846200 => data <= (x"07747f78a8318bc2", x"a30270c303625210", x"7b50d931597c415a", x"c06537412b570937", x"e42e11dad1343114", x"0f894676cad77a13", x"e9e29dd14e0a9542", x"c254eff02379c49d");
            when 29325578 => data <= (x"f95bf7a7eb8f7c6e", x"0daa2e38917b33ff", x"8f98c023107ef6b4", x"358a2dd3e1a6f6b1", x"7da3b25c7580318c", x"f2047a32e2b28224", x"9a571f252ae2f280", x"33a5f80409de68d5");
            when 2296082 => data <= (x"d31662842046a59b", x"9501a73aa0c32bbc", x"b5df0cf72ec75297", x"5dcb163bac59e95f", x"22a93338d330ae6a", x"5798cacb802b9b54", x"25ba4482a963a2f7", x"b1e8576a8ec34b35");
            when 17809698 => data <= (x"c199ca62362eb936", x"5331d2a490b5f94f", x"e45fb3e20c8f84f8", x"ec95413cf1180836", x"9c7c8b4527b79add", x"f38b454056c0ecbe", x"f2a871317f21f0ee", x"b997f356c01fc9f7");
            when 13724359 => data <= (x"8e62c55ea40e241a", x"3ed7de010a019691", x"ea9e3f982867e188", x"5e384f997501fa5a", x"a6b72c91c11216b7", x"7640f5d4302d3526", x"b3ce4da1d8519ad0", x"1019282baf4ee35a");
            when 2249073 => data <= (x"3c22be200911fadc", x"72d7511c882aa1a9", x"11938080ef1bc472", x"e74bff19787b6549", x"8dd7f177f3bc3269", x"3dc715e85b655e76", x"84a07c7f45db8ad7", x"a8bbc1eaaeac095c");
            when 20514181 => data <= (x"09cb20cedd220532", x"6b9bc4aa8c7a60ad", x"2cc0d0cac73b3296", x"de65ebfe915b36a3", x"6d057d474f4bf34b", x"a24efa3b47a0953d", x"22f913c8e77b869e", x"4fa6561059c163be");
            when 3795614 => data <= (x"958a10c42d6d2ddc", x"12f756a4c069f44c", x"35549fd6e25082c8", x"ef32a779e762e37c", x"ebeeb1b46cbd2c1a", x"4f68a7938e8b22bb", x"656596c2ceceb7dc", x"bd7eb1b2cd34f5ed");
            when 23694150 => data <= (x"b13f5e461adcfbfb", x"b2300abb5662e607", x"a5f8bc3e97986b02", x"71dd792f4c5dc09d", x"70a4b4f5628cc636", x"37ac43c32bb1152a", x"a157466f05e81785", x"327135b7ce668cbf");
            when 18503068 => data <= (x"8632d35abef93929", x"1312fa34d822b7ad", x"2963ca8faae8938e", x"abdc5101aa80e9a8", x"1f926fb5e5cad09d", x"646b4d05204c0bb8", x"9e1b938fe7650d04", x"544b63ef34208569");
            when 29091013 => data <= (x"474a06ec094d2de8", x"1d3e272b3226393d", x"127c8932588b66e7", x"b41948ff3fa23a78", x"595c207502d8bdcf", x"4ffbf54331332813", x"4fd04256ed821972", x"d6097db0c4abfeaf");
            when 9912711 => data <= (x"8290c0865eb7bcb9", x"be1ed14b7030d3eb", x"a10d4c764932f4f8", x"549744d73ffde8c8", x"17943aae246b8dcd", x"a6ea8cd4d6c967bd", x"282fad64661aeb5e", x"b36635d6d6f85b66");
            when 21653916 => data <= (x"ef7c66d798c8a962", x"ee654c3417edc9a6", x"cbd189887c27e6b4", x"e7b4d31a36f25b00", x"4e40321c8ff8e28d", x"59ac287ab7d381a3", x"6c52d540e9674304", x"f700a93be5af5c23");
            when 21864677 => data <= (x"6f74db25763e6d0f", x"d24a41a5dde80964", x"5cf08ab403d052a1", x"8e9bb98868489929", x"ffbd45d767c19201", x"a1117dc31d377034", x"e628ef2780554ea5", x"ae5eacc9d9eed52c");
            when 8555639 => data <= (x"fc04911a154cbf2d", x"b46de860a8de29ce", x"e1031b0e66ad32f3", x"23cafca1ff75ea05", x"e32bb099dbc9e00e", x"1f8386f34152be0b", x"3e6e8663cca6c7eb", x"020cb2ee189a41a8");
            when 1384542 => data <= (x"447fadd7b8bd29fa", x"b3e3202b3ba6a412", x"d8904f3790dc09f7", x"2677c65aa914739c", x"acc83664fb8caeae", x"5cfdbdb9296878d4", x"2cdd5f9b6e127e6b", x"3bc5dabc73ecb8e3");
            when 8149842 => data <= (x"5747cd3461b4bcab", x"b10214901a478166", x"d1733609a95cf856", x"81424df5acbdf47b", x"46257d0e837d5a55", x"d92217ef9fe3dcc4", x"7a79e5b3b21bb77a", x"0dedf6314cb5d34b");
            when 6719357 => data <= (x"5b03eb8b5984b7af", x"d583b3d45d6dff69", x"0d8b8862ad5668ae", x"42ac10dda76fab2b", x"fe7a9c431c7fb4b0", x"9f686385d73804c8", x"98cb07c0d7b47bd5", x"5f76c93704e9a6e4");
            when 29818217 => data <= (x"b0cc87831ba85a45", x"a697f0ac2ed4e667", x"c6a2bd97dfc4b674", x"eb57140af0fff840", x"40ae5496e84e519a", x"37dcfaee1b33b211", x"1457970a8a07ad62", x"d57c8bffdcff7feb");
            when 10384367 => data <= (x"a0f53df66d76365c", x"cb05550352d6bc6b", x"ee77c9d160b2bb03", x"eda5d71050963de1", x"161906a1cacf829d", x"d12b8f4018048fe2", x"28992b33bb6dc2ba", x"800eb21cdbff3b47");
            when 31129953 => data <= (x"4abd09a49e3f9fda", x"124846e6f7f14649", x"eeb6e6ba1acdcc9c", x"11ad232a16c7dea9", x"35cf008c41680a56", x"4c9440693ad8dd86", x"cf852562a9fe1994", x"9e1dc9a97bf466fd");
            when 30685252 => data <= (x"282941911a3659f4", x"dbf608491e7bcff1", x"e1cd9707c7854005", x"1765387b794a5ffd", x"89e14651e4fc9dfe", x"859ec749a8490f66", x"9efe4aca634bdb21", x"ac31cb4a7c9f8110");
            when 25609636 => data <= (x"b404f5f5fddf62e2", x"6477a717f0e6104b", x"cacbcd53c6c6441e", x"854a812ee90b1a31", x"0288c88a5ee8ef8e", x"9fff0844ffef8dae", x"3ec36257376e3259", x"e62a490fe33c39cb");
            when 1046604 => data <= (x"a418e1c11ec924ee", x"02a40cbf12371a66", x"0c60a672cfd4cdb7", x"ba14819458ebdf05", x"501557eb281e2847", x"071ab1bf4a16e59e", x"48d55ccb0a1e0eee", x"c4b2f794c6c65666");
            when 20744827 => data <= (x"2f075ab9b9e34c45", x"b9b91f75e49c5796", x"e255e63611a627ec", x"c0e543b7f5fd645b", x"445cbc640c6a74bd", x"dd3bb08f25635d09", x"c45ba0ccd129568b", x"119f86a81bff7d64");
            when 1103753 => data <= (x"0c29fa54b695b7c8", x"b648a9451360e304", x"a1c04d8371257499", x"0fa17e2d8a859e26", x"d9dfb491cc8bfad9", x"fc40373b00c0effe", x"a33918e8ec265add", x"fcef6809061647db");
            when 28110477 => data <= (x"e67f17d7d091e805", x"418f4488355b780c", x"63828fbe9ac53e1c", x"9d3d9588ba6d92bd", x"8cf2209ed96a4f61", x"aca0e22df838fcdb", x"0bbc1db10e483c56", x"f14cbb152f2742a6");
            when 26397405 => data <= (x"b194daebf35fc4cb", x"a35f08901c0c1566", x"4c86c484a424a82f", x"d5b413609382e78e", x"38125dd0d38c77e1", x"5f727e747e3646c9", x"a78a98f8e5f359a5", x"eabfdf2568a39066");
            when 8504798 => data <= (x"42065fcc02f85fd5", x"a51cd97391ccdd5a", x"c2848c4e9cecad6a", x"86861e47fab31f1d", x"1963920353434980", x"d8e19343dcb956d1", x"145977fc559001d9", x"ca8d3ad29dc9ccdb");
            when 15429412 => data <= (x"4e6cac0351fda4e2", x"5b61a2c866821f9f", x"829cee9f56f0efe6", x"c813466a29376785", x"c8acb32968ca036a", x"fba85de0a3952973", x"34d12f5ecbb6c843", x"0f723f02e1ba024f");
            when 30777390 => data <= (x"89d74028db014368", x"8307ee07cc4413cb", x"988e15d0d2f6a456", x"73917acd8f084232", x"2aa34e05be365c1b", x"2cb10ebba15414eb", x"d18f1a3080dc9fbf", x"b46dad82b06bed05");
            when 9944242 => data <= (x"cd9e945c15948c49", x"71fd475fee840551", x"91d9941499ae0174", x"48c29736ae9432e4", x"d8109eacc874f6b1", x"3a2a9f5c9a7e2ef2", x"ab773e640f5870e0", x"ad51277dd3c071b9");
            when 19139741 => data <= (x"99d40ebbb95e07de", x"eefb1e099391bbe1", x"cd6b4d2cc68a288b", x"81df1bc4be3360cc", x"53eb0ff03727a285", x"8b418f4a690ef3b9", x"cae6ac8640573de6", x"8546f572eba3f6c6");
            when 8274329 => data <= (x"d4bc27b470c5093f", x"c81c97b259e0780c", x"61fc5d53ac578769", x"b64f0bfc23fea575", x"c247017c847220fe", x"32dc476297ca7bc9", x"e4ee650177681397", x"d44181cbcc5ad0c5");
            when 4804052 => data <= (x"cde8508dff26eaca", x"d64b0503232a5fd6", x"c5121d86821e7aa8", x"3194d70bb93639c7", x"6ce995cc534495be", x"5b65267772c58b68", x"259943a4332e3eab", x"6696616ac6e7cdd4");
            when 1662695 => data <= (x"dc8310534ab58447", x"acbdfe8baccb5203", x"4296d8888db733ad", x"56cf934cc213a6be", x"958889cbeaae6a1f", x"618d576c54f220b9", x"b8f17e357d9845e9", x"49610abd29a48813");
            when 488305 => data <= (x"baf3f11fe770048c", x"a279f1bf80468dc3", x"607f4c64b8e4533d", x"98ca58208454b9e8", x"d2ed754f36d43510", x"9f40fe76abab17e8", x"529d7ed72713383e", x"8d18e90ca64910ff");
            when 11122762 => data <= (x"556fbac1766674a2", x"e1ead26e453cee15", x"2356dac22415629b", x"85396cb6387c7350", x"d735bce660741f2b", x"d74e669d29ae7b4a", x"260cbcfc92bc099e", x"63e283b48800ebaa");
            when 33333011 => data <= (x"d2e47d1f5e6b9bc7", x"04c9cb78a5a6aa4e", x"41271fc67905b07b", x"139cac9b741b3e66", x"146cbc72fa6d0a90", x"32d3b8d5427dadfb", x"b2e529c6d8c8e754", x"c311ef06ba8188e9");
            when 8064373 => data <= (x"c9002bf563ffa46b", x"12f488225f10209e", x"558c03573592e289", x"75beea733a15d0c9", x"28e2f9f40abbd199", x"4a64a9365583a21f", x"e4ae5527f804b49d", x"75a32af61160ff0b");
            when 17563212 => data <= (x"b5b30b4c20ef2502", x"0213ff243ba24742", x"09f0f4a11e3d06b0", x"360d6878484165f7", x"c815fd17fa00ac2a", x"e396bbb5c1d4e825", x"b5cbea694329de85", x"ae820664184e4eff");
            when 16142394 => data <= (x"c38769678b958a79", x"eed90b4720da2eab", x"c1b4501a3533d961", x"fa76718875f937af", x"2082d32a7db1c717", x"3075e606eb914f83", x"329971c6997596c0", x"6180d8803038cdde");
            when 23555098 => data <= (x"32354e875ef77ab2", x"6746f0388a03b2da", x"f63ebdbd58725dcf", x"87e668ea3b6e9f27", x"9852f4b9a0563254", x"ca3db0a28ccb7b2f", x"f6fb45ae4ce061d2", x"4a04d222ea9346d6");
            when 21437663 => data <= (x"eeb5712030bdf6d3", x"a5910b88043b6083", x"5781d1a39009ced7", x"02e8cf802f99410f", x"3db8f72c3e400176", x"67b9b56c8950e6aa", x"cf6ade983c54d246", x"b4fbe07519b351b6");
            when 15715942 => data <= (x"579753c04f5f267f", x"07538d95afb4a24b", x"9aaba74ea2257f99", x"985bd9d4d8152f47", x"6a884bdea6f1177a", x"8fc16274c71408d0", x"06a16a76e2f2e645", x"4b39e9624e57e516");
            when 26674072 => data <= (x"7e1f01a267db9450", x"14029eabcca14739", x"1f8b6475ca7efa82", x"4db3486f262a176d", x"2a399523c550a60f", x"66a4751261db1331", x"9e9b179a01f942ce", x"52e2d0174336ad10");
            when 22315005 => data <= (x"6c78680e51aa6ee1", x"223dcd727ff4ff45", x"9ff6f27a06a08c8a", x"143b6bf09a46ae49", x"bd5cc8097cfe4c32", x"20c601c8582bf8a7", x"bc8b2a9ad83fa419", x"0893d6866bc60d28");
            when 10583341 => data <= (x"dad3336690e44c2f", x"3d2bf2773dfe9b96", x"97d0319831eae950", x"90a28336eaf08d80", x"f5c7b2480c584da4", x"8520680faee75878", x"456f2922a4321003", x"c64bf176174c0abb");
            when 26461260 => data <= (x"838a3dfb14398555", x"f3dbee55bae455b5", x"a5facc0600040760", x"078674a033794ed6", x"3c6960cad443e34a", x"daa27ff1e72ad84f", x"81a6474977eeef35", x"071420c662cf49a7");
            when 21833960 => data <= (x"542ee7f907e2783a", x"041e3faca253b9b5", x"36bf79b2cf74945c", x"c69ad60f0f7abc87", x"2a2063a7803bbc50", x"38bac5de17d5870a", x"e2a4e25631260095", x"fa96ad528df8a4a1");
            when 11789454 => data <= (x"ad11022e7ad0ff3c", x"2031018218906d61", x"bff8cc5f5e8733ec", x"0f7d96084deebfca", x"e88489787a9aea78", x"0b55f1b850d6bb2e", x"513baea50e377be6", x"9dde6184087ee0e9");
            when 24625508 => data <= (x"2f4b7cde43b24cb6", x"4372bc9271ef5095", x"ec32f0198c141d8a", x"1f62b110503c8ed4", x"a3e792deda527c7c", x"756701cbf3eabef6", x"ec435ebb56169133", x"47434582ff0e8d23");
            when 31160303 => data <= (x"fae4e3445753d572", x"1f20be15405bf408", x"a0d711cf20962db3", x"8df9712ced3a7137", x"d9fa7f1e6def40eb", x"7a406e0f95e6617f", x"a98c552b1a933390", x"d85621dfe4b1d733");
            when 30060542 => data <= (x"456c8be67332cd05", x"fb30b5482246dd94", x"5dffcb2372c01e02", x"2e756d6f3a54d2af", x"6ed5636bad01ef6e", x"d28bdeeba8dbd481", x"33d25b8892600a07", x"be02798d70524989");
            when 14567377 => data <= (x"6d44cea0835fa24a", x"fb109a11256fffd9", x"5c923307985cde8f", x"3dc83ef744217e7c", x"7a51c7f6f8f48ff2", x"ca37ee45fea7d448", x"8c0bfce1cc991f18", x"d92149b3577954f8");
            when 26060933 => data <= (x"fa3d0f92f1e4c53d", x"5c3c097f29b86b8a", x"bfdb4fc1fa7d0d8e", x"f89d39138588074a", x"527096460b038307", x"e193da9077425adf", x"f2e3f6401ad75899", x"3f8fc23ab1dcc84f");
            when 25017249 => data <= (x"7cb853e82b2b3b93", x"58c7bb8adcb0ff49", x"ad71e16a3f3b29df", x"f42614f7b4d24cdd", x"4748f388dfbdfbb5", x"83afe6b75578a358", x"879e9456e9b5cba2", x"dfdee6a0c6751635");
            when 29161107 => data <= (x"eb5f1651e51bac4c", x"9dbfda315c357fe6", x"674a54947665d851", x"62cdb41b4ed28195", x"785e5e19d74651a3", x"02129175aa4a8cdd", x"512221025250388f", x"cf2eb469b9ba589d");
            when 23813018 => data <= (x"436e95cb7e92c707", x"b220f8a743455c5d", x"a5bcf81016d42a9d", x"7a2909f4de46c2bc", x"1227efa669164564", x"82268f5784041447", x"e0995460be5751a1", x"337959c03232bcdd");
            when 27822704 => data <= (x"2ccd7109f6c7740d", x"4ceccb3a2910a0e8", x"36612366db656201", x"827cea224b38f658", x"73cad4081cb53129", x"ac261e57d168bbab", x"9587d6d0441b1fa7", x"c553f52990847c3d");
            when 30708718 => data <= (x"2adb46673f6d839b", x"f3f39ed39fb76728", x"2a354593d5b43ed5", x"dfeaf9679b754b93", x"a810be77bfae4bf5", x"ad91992df3855417", x"226d290173ee2e9b", x"4772ef434591f476");
            when 27194331 => data <= (x"1346cc93d62578eb", x"b9062b5b266fa57c", x"da99eae1aa2bf3fd", x"b7d7e9a91fdc69b1", x"d324abd2eab4434d", x"5b3ec0e3cd44d3a2", x"2f3a76b962d2817e", x"445efe30a44b914e");
            when 18612442 => data <= (x"27576e6da867b425", x"7b08924fd3b19c17", x"933e00e3e3e1e4ab", x"80463672838bd02c", x"956a7de2de33ef9f", x"a1f3e0be313de574", x"00984aacf05f080d", x"bd39b7a0214baec5");
            when 30585086 => data <= (x"caee19c8a73f4dee", x"19ca24196ad13f8a", x"c0656ca365cfd5a4", x"6f8b21160e189797", x"69b6d4f204e2e72d", x"a9e831e245f1af0b", x"9fe748fb0d23ba9d", x"5af7028c44e68d54");
            when 23036731 => data <= (x"6f02ed591f7638b0", x"d6ed52c7ca0953b5", x"9e17be16b401337c", x"9a2b17ad0785b556", x"bddbc34a63f61403", x"4f3cb0beac21ad20", x"03003e2458c5c93f", x"c8b2c96fd216bea5");
            when 26064830 => data <= (x"5fa96487bd37fdf8", x"416af3cca4589c85", x"dc3c3f33db6b96f5", x"e6068c0d6b4bb041", x"c4045a62d92a58f7", x"abacac28eb6904b5", x"7b70482643302a34", x"ab65ab105753f451");
            when 31690957 => data <= (x"742fb50e8a1d8190", x"c17aa1a6554e5542", x"d7a090fddba3fb97", x"e386f7ea9c576aeb", x"23597c68634eb831", x"74e4c4ac68ed2d3a", x"7de587bfa5c60ea7", x"ba0125e41a88f153");
            when 13095987 => data <= (x"dacfb456eda015aa", x"de3e605702b826cc", x"c92d102a5aacc037", x"92224bfdf8743325", x"4928779df18f50a7", x"62473536561dedbf", x"d993287521f701cf", x"12f9c573e2975888");
            when 24097907 => data <= (x"84bdfccb0a8a0771", x"30dc0dfaeeeda94c", x"858ed59e44c545ae", x"25fb4fc0ebfea3c2", x"d191a4a5d2f3db75", x"2986e8d9d256ac76", x"0787978e6b0ab2ba", x"0b7b72c1bdc51475");
            when 32983731 => data <= (x"a54d9f62a49029a9", x"5ae1209a3ac6fc04", x"c0bf6a3df357d10c", x"0f38bc85366afe03", x"f2b2a2a1d8011dce", x"9e8f7a9ae7b6c0b2", x"e9a6513f6753c151", x"a2fb2c450b6629ba");
            when 27574483 => data <= (x"a5edc0b16eead330", x"ea2c7a49a5662aee", x"77195bde79673138", x"4ec9a0cad1350a25", x"413152d2c2b0e7b2", x"67ed542a0452006e", x"b9049ba491f80a87", x"1e16a635d1b5cc34");
            when 12950330 => data <= (x"5fb096f2362061d0", x"ce882aea8819c06a", x"fdc93e72cd532ecc", x"32f236fe8d66c07f", x"e555d4cbe0b56175", x"99f6c714dada9c78", x"506c9ffa1500e001", x"9f8af046b4e068a8");
            when 16852888 => data <= (x"d80d171b55bf3eac", x"e87c462366a3a167", x"aee3488badec33ae", x"da12f5c6d3493266", x"4e6b524f815da052", x"8881fce54daff2d2", x"45ac38a07bf95bef", x"7401d29c4c368113");
            when 30707361 => data <= (x"5926ccfe95d6ab04", x"b54646ddb2d4a5af", x"8d08acf1f5134273", x"074289f448aabb32", x"1b7cd7dbbf6735fb", x"5d75ac4c5cac4909", x"33dc08112f2ee017", x"8b2c5f0dfeef3165");
            when 8006759 => data <= (x"83fa462f30e69dd9", x"5b38aea7f41dfe3b", x"278bdb2b86667d13", x"3be27bbd71ad651c", x"5b4f9c503b9e0de4", x"76a1f2b349b13de1", x"3ed2c5224db5f0bd", x"f8a8cfcbe4c5be9e");
            when 33925965 => data <= (x"208bc47f61cac685", x"49044eb10859b11b", x"c2d2058703f328b6", x"ee56cb9ab3e30137", x"e6569c6a252c086d", x"94ef7970079bd20b", x"fa6806787d596bad", x"74525c2d9ba828f0");
            when 19178210 => data <= (x"a05eeb4e2476a07a", x"fb0a43b2a9f5ccb6", x"6a97d53faa6ea40b", x"c6ddaf30ab9fc25d", x"67315c1c114c0012", x"77bfef2b93653641", x"aef07c47f170e3a0", x"8f1e387672572126");
            when 12440858 => data <= (x"04ebd311b69d4a2c", x"272e85290e24624d", x"434c9ce2cebb6dad", x"47e4609122dd3be5", x"b8ada055f2cb69a1", x"bd89e00a397d994a", x"aacef4c8104d6920", x"3184679f7e3a31c0");
            when 25927747 => data <= (x"23a48e7e4fd2123f", x"fd63fd9f3a736fb2", x"b9689ff74d633ecf", x"90b86633f6d3a2cc", x"26966fcf99ee30e2", x"48c83435dbbd1fa8", x"a099c81a083f1229", x"187d932df2f39fe4");
            when 19606792 => data <= (x"05eebf3883eeab03", x"7070fc916baafc47", x"4923eb643c5e90b7", x"809cfbf1ac9074a9", x"a049ac06e73ad557", x"c994b9f00c47a3da", x"1c5a4d2086c0a039", x"f757a5ebccd78be8");
            when 27350143 => data <= (x"89d9995d4ce6927d", x"6ad26e3845d2d779", x"f4576ba405e4abcf", x"51e8c318e2314196", x"9a7372dd69581657", x"f3ec3c92ce057779", x"d3053bb75fbf0208", x"aae9c5f9f2112e3b");
            when 3601238 => data <= (x"a198843990edeb06", x"699acbc4516cbe60", x"ffb9d1886b770e30", x"8a016ea605313d01", x"4434d2f696fff572", x"c84969b17e59bf69", x"6b8ecb2dff8fe031", x"f48770c5bd22cdff");
            when 32811514 => data <= (x"86ec485161dfbef3", x"805db35dc1049452", x"05f0fa3eb21b91af", x"5fe934f4b63ebe2e", x"57567b736df32841", x"230a7faa90ff220c", x"74aa7a5845cfc4b5", x"85185a4f410676ac");
            when 13723430 => data <= (x"48ef138f1a6fa3e3", x"692ed6add578a2ae", x"39d1d7f9cf3c4545", x"92ed83199ff2e553", x"da56d41f38455074", x"8c613120f80dbc35", x"bcf331663fc23cfe", x"fc7b4171acd91936");
            when 16907635 => data <= (x"29011db26f1ad622", x"88b180d21e1c4958", x"fa05ed6ef4254067", x"fb767626ea4d8207", x"6bc425bff6839d6f", x"c440f01fa383c219", x"db9b93027ef75c01", x"7291a32d3b3c1280");
            when 17124167 => data <= (x"821d1bcaa99367de", x"ffd1511fad4aa39b", x"d53274775550a9c7", x"3ca25756213c586e", x"05c4ff6146bc0ebc", x"6c6c8b63bd4c3429", x"02b0b59b230f130b", x"e0e20fe1ff0b4762");
            when 7423330 => data <= (x"aad9b644129d6b9d", x"2dc52c69341f41fb", x"3cebc0161df2b095", x"81b5bbc3c6d8418d", x"a04c787d7d9e66fc", x"9554639c3eba84f2", x"6afbea662790e319", x"7143e25d16186d29");
            when 30565862 => data <= (x"8bdcdff8b2ea8b69", x"08580cafc77d6010", x"838d32f7f3997d0b", x"2ab939af369b7bf3", x"dc638c209b579e05", x"eccbac63195a0e61", x"6508e7c43327bf43", x"2cfdce738ab140ce");
            when 17280023 => data <= (x"099958e8cc73c5a3", x"2ecbfe9a6e169680", x"01518298b8dccc84", x"a0e0ac5840ed38bf", x"d6cc3b30ee42d66d", x"795a83f70f027a20", x"ba5139e5d61c246d", x"72ac80f4573dee99");
            when 6318643 => data <= (x"d3cbc452ad99be5f", x"eaf487f9d4ca90db", x"2e0272b2e7724a82", x"6bc8c3c58601ba3a", x"ad8430463c60413c", x"dce3552642127047", x"de68a74a8e4e8ba5", x"6598f6dfb723fc7e");
            when 27387156 => data <= (x"939286156c89aad9", x"578997365987d058", x"eb99754f0c2f0b30", x"5026ace09f24f6e7", x"5a7fbba21c0ad160", x"d85d053bc8a70ece", x"94c54ca18e447cd7", x"9c4ffd6a40b2cfc4");
            when 7347702 => data <= (x"ed8a0e77dd2e2efb", x"3c3cf6f2e5dfc4b4", x"46c86bd47efd5507", x"473675b240313a23", x"c85a37668c14be16", x"fb76c88178208b61", x"fd83c1cda67a4cb9", x"4ad734b6b772a78b");
            when 29276280 => data <= (x"5fdb21e2ff008812", x"e4c6740438b85210", x"69abd4e023bbdd79", x"9ced7674e217d23e", x"7e9b80fba6781cbb", x"15998d399fe47926", x"db25e9dd44d707b2", x"5256c8248e401fe8");
            when 15839464 => data <= (x"5c60220ec8f81986", x"bf4d632529ac5191", x"f2629be0fd189c16", x"33013638e257969c", x"fe58d0133dc39529", x"72194cb842870a82", x"2fc89b1a3cb77ed4", x"d28f6f5fc27a0193");
            when 21677377 => data <= (x"88d7496117f7daef", x"b01e6e3d6e4cf4c6", x"bd02a3ea6e09d2be", x"12851f29bc2c7c44", x"5e8a4e2912eb1eb8", x"6c6c2d477a08e005", x"f325a60a115025ce", x"a9ba11653810b8bd");
            when 32118315 => data <= (x"d3cfceaccad73719", x"805b078195525afb", x"3ae4e07ddfa3eadd", x"0b8169e73bd20491", x"96b6146131e96593", x"c7f6da11b2278a1f", x"2f9c174ca853fc0e", x"b6e6b8671050ab2f");
            when 2667965 => data <= (x"69957e36e05b90da", x"e6d39012441cbb3f", x"5b4845ca673a0ff6", x"e8470ece0930ca33", x"43adcd17829bdb49", x"2d6a41f9e310caf1", x"98ca1cede95cea56", x"c6a2dcf0d559352c");
            when 16814232 => data <= (x"d26e3b715caa3f8f", x"dde54c61e174ae76", x"aaf684052df9c4f0", x"61d984aa5d712a56", x"0b87330502a719ac", x"7dfb2f805761e3ed", x"cdc2582d8ce200e3", x"112b77b133d20e19");
            when 25719715 => data <= (x"4fb972d01206fb5a", x"416f793a7a4cde11", x"23ba255d61a2fe1c", x"4ef0c56b54790819", x"f2fe54947c661dee", x"fbf15240d9dc8b04", x"56528d631a48a749", x"a8a3aa0e2346c07a");
            when 16184243 => data <= (x"715ea077a2ae50a5", x"72c45cc3591752b7", x"c59fde1dcb346966", x"44aaa953465e1f0a", x"c6a97dabde0a48e0", x"848d8bec3ed077e2", x"dcba551a4d39eee7", x"8d0c24f26104f951");
            when 16352961 => data <= (x"30fadff1de2a61db", x"5751cf2d6fb873f7", x"e4817e9b7c453da1", x"1a44494eda66e506", x"f33c5159dab0edbe", x"e03dd8acd0503008", x"e3bf2916a017b081", x"4edfb09b00ea0813");
            when 1637022 => data <= (x"288085034c7c50e7", x"721b43540a099d3c", x"dc3e382aab4500dc", x"0055ee113b4f8b24", x"75e3c8611549c076", x"b5398ce7147bac9f", x"5fcb1a0b24af8a54", x"be1a1c6b117cb7cb");
            when 1655190 => data <= (x"3eec50a1c336c90b", x"599570e10431359e", x"c0824d99e46e0454", x"d848ccb3c1163057", x"057c6da6661dd823", x"848ad9c727daf18b", x"fde7e642e9cbe73a", x"323621449103751f");
            when 29206664 => data <= (x"4cb48087041d7840", x"e413a01a5d0b0ac4", x"599a3f24f89d976b", x"25a544f9c8cde704", x"2a14a28835c1917f", x"302dfae250239b48", x"e432bae0608dd388", x"b5c6e7ca294f2b02");
            when 2104420 => data <= (x"8d08ec89dfa1469a", x"e1d46815982555ef", x"3d580cbb85cdbbaf", x"8672153052d36429", x"38643a0786c9b648", x"bd8a8813a4a42cc3", x"855a1541355e21ed", x"f5110ecba94b0f65");
            when 2237562 => data <= (x"2feae9d2e04d8dbe", x"e16d605b820d2e3a", x"61c6fa9231a4328b", x"dbb13a01b938ebae", x"65aeedac97a6a935", x"a00b63ebfd767721", x"e7b9389543d7603f", x"ee776ea6273aeeaf");
            when 10939535 => data <= (x"f128bc3a9935d7e6", x"7d08dae35d606365", x"c1f82e3d75884755", x"2b1c0cbc16e84446", x"75a2f1bfa9ea9c2e", x"0e0037a5aae0c732", x"8ec06c0af1e909da", x"9808b0275a868c12");
            when 27603299 => data <= (x"5b24b82ece72f157", x"ce6d0b3fd291bbc0", x"74bae11ea0aa8b43", x"e33aaab16bcfdeda", x"8ab4e329326286f8", x"3ac019b2f4bd0dd0", x"d1aff4966d974464", x"a2c63640d5ff76da");
            when 11743432 => data <= (x"2dc3b5736eec6c2e", x"a5065d1928564345", x"1a37807cbbb2c4f7", x"b056487490a0744e", x"b71544f79b22c87b", x"25ef8dde94ecd271", x"0175c4330ff420a7", x"534c80fe2050f46e");
            when 28774651 => data <= (x"8463f5b054b0f0cc", x"08178e6e19def517", x"6da4f9fbc7ec02c3", x"30df6a28a66adc4e", x"8d92d3701e7aea6a", x"c164c3e0de75a7b5", x"54e328784b8b5ed7", x"c672e0ef04fb897e");
            when 12353712 => data <= (x"ee578346e68f44c9", x"fa6fb1604dc5a8cb", x"a5845b84789ed51c", x"3bed3cec3bd3dfc9", x"2cf5cfada6edac5a", x"ea177cce8ba8ac5f", x"1eee4049e9729e03", x"072ae05788d5985b");
            when 18698398 => data <= (x"a2b043a98e3001a2", x"9b6573e72c1a8837", x"0460a41d69856137", x"35f7d41314a48c1d", x"b3db501b9db64a4c", x"9299373d7c59ec18", x"dd4408dddc7668b6", x"ebd8652fa886b2c2");
            when 18667435 => data <= (x"55eee07542c2fb0e", x"6d2aa4ce1b5734ee", x"9b8ce1e5ae2d5a40", x"51e6ce8a2331adbc", x"ee841166a563c0cd", x"59dda689fa006431", x"91e45aebd0dfec88", x"0d671413a4920d1c");
            when 12476288 => data <= (x"a196fd1c22332b6c", x"a07873d3fbc7b606", x"21bd048df7d110bb", x"1f71809ca6e8bba6", x"cfe4564ac37d399b", x"935b2ae7a5217470", x"2cf70b257a5245f0", x"0b77da12c2a718a7");
            when 33053539 => data <= (x"bd8857ac1b887dfd", x"6e4562ea5da887ff", x"c02e7eae3fafddae", x"d19014fcf0342309", x"067a5d504aea010e", x"ccc9edeea54b4b02", x"34c4711b475e15f6", x"0d1ba9cda2698b7e");
            when 4379060 => data <= (x"e06c85cd171024d8", x"c4c5e203b53e9627", x"ce11619b1aa66e4d", x"a7945ae71fd42818", x"635765fae2d70752", x"4dc84cb2a824d0e1", x"b21abd7c7a73d5eb", x"b96908fe51282e82");
            when 30013201 => data <= (x"dde7e4d654777de1", x"9ba191dc9d35a392", x"f02b5a1a5de24fe0", x"9cbc5acac2840503", x"5b5ceb6b11ef782c", x"1c7adbf37565c492", x"6b70cfb627efa8ea", x"813823c1a63231b5");
            when 24753965 => data <= (x"379449fc055ccb9b", x"6efea25c6a70fad3", x"3d0c851b3927d1af", x"65496e0ff67b98a5", x"8ecc3ae3e8317f85", x"9b3422d6711630f2", x"c2fac6beace373b2", x"67d234ecbdd25bc7");
            when 2648512 => data <= (x"3d7abcbbcc1c2bf5", x"8f578d89f1d27bfb", x"abf79946e6e247f3", x"86b9e071c40cbcf5", x"04a12bc958e8292e", x"8d1aa245e945b991", x"aebb496b5cc5ec1e", x"e1cf0f564506c765");
            when 20847342 => data <= (x"fa761e4223545c15", x"6c0d3f5e95824d07", x"5034b1f85588ff75", x"0bdc6cc031b3ecb7", x"a8c0421e83db7cc3", x"b1ec6b2f48cf8445", x"6227ad8a71a93a62", x"9c07f1a961f1a93f");
            when 31721812 => data <= (x"7af9636369db2631", x"07d58c80bd4940c3", x"32d2334e6ea672e3", x"01a4415046cbb7b2", x"94c32a74db2f0c22", x"87a67b6b43cdc989", x"baa62a3b0844b112", x"d4135a3418898eef");
            when 2254298 => data <= (x"c5e1f7ab684b5b34", x"794521e3abb88b4c", x"47a29733b6f7f983", x"55c00096ecc974d1", x"a827ab5fe4fa05e8", x"760933a79ee483b8", x"bf5766cae16fd81d", x"8af0d93d1eca9411");
            when 23226381 => data <= (x"fc94a05a51a5a46f", x"478d0b8db644026d", x"9e8c92f5bd967d48", x"5d716c7b8d61e5f2", x"e0b0b30b425035fc", x"887e038bd6dc5200", x"1ea725cd45d06543", x"400898b813d3f31e");
            when 18305145 => data <= (x"5490d359d0f4db46", x"7365e101404b0bfa", x"ce9f833656b6fc5a", x"ad665300c8489bde", x"45974e3c7bfb31db", x"8fa6b7e01076da9c", x"a322483c875cb32d", x"4b0135019f8126f6");
            when 29048619 => data <= (x"3d69baa934c36f01", x"d046428f33608110", x"796ede560402d1e3", x"5fb1f2bb86b4afbe", x"68e8dddd01f6e36a", x"b5786fe27ed25c0f", x"bf72bad1185d6a8d", x"9abdfa693385dd8b");
            when 23128882 => data <= (x"3da4d80371fd4eba", x"25a0cf2ea6168bfa", x"011e4acb50fd86f3", x"eaaa152d5b20a8c8", x"418738fc34274988", x"caf7b4cd50e9893f", x"c05cf13677132b09", x"f54ba29ee887e64e");
            when 9539044 => data <= (x"4f77419f51d1acca", x"51c7474e560762fe", x"39b2af43a30fbf1f", x"a8b464bbe2f91e4d", x"7ca72b99be69b1f7", x"bb982f70d79065ab", x"104a4ef59486df61", x"c66a24deb7a5f959");
            when 7855112 => data <= (x"eec00de48832dc0e", x"ac61e19f5cc8bad3", x"27f85e4225ff05cd", x"d5fdcd313b4ceb28", x"086931454dd91b74", x"e7ebf3e447911d3d", x"0e5987ddbc659a98", x"644338c47dcc7069");
            when 22919281 => data <= (x"45a4260b35e4f6ce", x"8f489f5251c4aaa3", x"fc1d06cf50f91770", x"e609e39c152bc560", x"c0f16e894d5c7a65", x"b04751765beea6c1", x"f452ff57436ec071", x"d65dea416b21dd0a");
            when 10309824 => data <= (x"44486439fe04bbe7", x"02255cfe7cbff0be", x"2b0a9c7dfd0d4da5", x"a0a939d26e83dc79", x"9a025593c9d4e945", x"634ab6936dbc04a3", x"3c116d2f6950b9ec", x"e27c7f827bff04fc");
            when 9441377 => data <= (x"192bae740762174c", x"139a7b6fc596a4ba", x"b2eb3d1a3d8017a9", x"2424fe8ec40b1731", x"be0294479d17cfa0", x"c6d8fb554570c022", x"08451e0a92b8c92b", x"81c741c1ba26fffe");
            when 15067748 => data <= (x"8ca6ed84613c7ef0", x"1f244354f7cc9db9", x"e951b17d87391cd8", x"9ac4f12b5994a1c1", x"a33257817e28ab26", x"a268ef9d7cd004fc", x"bae4d9b883a17e3a", x"878d61bedb50f48b");
            when 4815170 => data <= (x"b3e3ef04577c6522", x"a2112cb777d48ae4", x"cd1ad095d4a8c7f6", x"dbd460d2941136dc", x"dbb0702cf826b36f", x"4775726f6ab9b64b", x"f76db82cd60bde61", x"eb375ce5e6787e12");
            when 22626657 => data <= (x"70ad749d7d35a552", x"e21e5e075f6479f7", x"acfb17e18eaf5b43", x"4abfc57e685538b8", x"9bc692b34ce29117", x"8c7c73cc22b9562e", x"4794bda6fa407966", x"458fe63accb1f893");
            when 2268491 => data <= (x"17b74fe14f70e02f", x"86ccc7640517ac10", x"1b5ef486e78e6b09", x"c607188f9038fcfb", x"e52b23cc6317f02a", x"e8d2b7f0bf96e8bd", x"b40fa9bc0f3cae2c", x"033ffd4b4d8492ad");
            when 21238280 => data <= (x"3389ffb49a55f92e", x"ea0454b725b794c8", x"f0f9b044c32fa0d0", x"e60baf9e1805006e", x"5699867dbc686720", x"d807377d56c9add9", x"611fb62f0e9ada39", x"d5ebf7896f5d8ab1");
            when 33797793 => data <= (x"ea62b6911a7c93fe", x"60b0c067bc5e28a6", x"ee3e15323665b255", x"bafa0bfe3fe76e6b", x"5bd93a7c0478268a", x"adf7bd762d862321", x"7929a9f665289f0b", x"0cc47c5cf39c32b3");
            when 19310576 => data <= (x"987144a70ec8eb4f", x"f38f79e99eba8c8b", x"a53babe8b82f02ac", x"9d7852a6f9ed35d5", x"1932d999414cae7d", x"e881a123291c4144", x"ddab764823d04234", x"0b7bc2d2c5b2ff1d");
            when 9484671 => data <= (x"9a4d0fd2325aafd8", x"74277d821443829e", x"0d66a89170a95e79", x"987ba167bc51d6bb", x"846c7b0c20573d91", x"22eb6566c223949d", x"5247781b332ddc7d", x"5f7d581722531df3");
            when 4414903 => data <= (x"29c46c0f9b2ce037", x"39d9bbea10b7f61c", x"a95e7b1d8b30088c", x"4838a3bbc2085a3f", x"daf9b8d5de194b7d", x"e56c1a1e5c9b10ce", x"4f752b9e04b11938", x"482b5965cebf1036");
            when 12614246 => data <= (x"5364e529a0a2e464", x"26f38a65044d9779", x"e0dca354a27b13a9", x"c21f93c38306994a", x"a915d55fa1b36fa3", x"952115fc44c54405", x"3f0850909677ac77", x"2e1e782721792080");
            when 15945253 => data <= (x"a5ab35d5f54e9a2e", x"1507dec0a7e9ef09", x"127bd55cfa9504c8", x"6bf49a17ddbff5fb", x"807411315df060c7", x"61c99fe57209ae5b", x"9f4a5948a58825c5", x"d71884f9a7651048");
            when 23408289 => data <= (x"0f5ddba1ab04da05", x"aac35d821ffa6e39", x"f8834b84252e3508", x"4c649e475e9dfea0", x"6e6026ba4dc73de3", x"5c116f19b0f74282", x"9d5ebcc574a51375", x"e618339cd0b409e2");
            when 29015054 => data <= (x"22e044361a7ce37e", x"dd033cd854931e02", x"a4591d3bbcd313b5", x"afa88b9e37b9380e", x"7845628de3a92f55", x"aa5880a2f94d3647", x"1516a0a2cbd58492", x"a6b34dcf89206661");
            when 12684767 => data <= (x"ce671e0860d72460", x"f2c655559dc26133", x"9eb2191717ca4da2", x"c39f4fc886627f79", x"9768e0b69bee0885", x"e9cd651f93d744c7", x"81b97c8e950563de", x"44196f90c4f6fae6");
            when 28463303 => data <= (x"5813c6d5c5438acb", x"a49447639d07d3a2", x"120082c5d06ae817", x"56c05f637b797cd2", x"e8de06220a42776f", x"0891f020c502d550", x"ad251dd060ab4c79", x"9681da3ded8d6384");
            when 2167672 => data <= (x"a39fdea3ef1880d4", x"7763e60d55a4d0af", x"5a2ff1171cd85b6b", x"a162b0c329ab7e54", x"f19d1ec84f535aba", x"7bd3ded8fd3b6ef8", x"434b7a8efd69b9ea", x"efbb9b953d6c1011");
            when 10001704 => data <= (x"61a0ce849083ab76", x"c9944c234397008f", x"7f70aabb9c0ecf9f", x"d8369fe13b4c7abd", x"4cd01a0c0fff0d88", x"7211b9cc5e535fb2", x"3f6ff0427ab25f5d", x"a1ce17b362c2af74");
            when 25712050 => data <= (x"036bc87b29171246", x"507df15b2967e1ba", x"e25d90beeb4fdc15", x"76cea82ff5c08ffc", x"f409cabd2cf109ba", x"2f3fb22f0afe2d4a", x"6d4a633ac3e293fb", x"22b86a5cb7521b89");
            when 14145968 => data <= (x"d3dc85ae8bcd4190", x"de4516bf961a6ce9", x"d4b2ef1b8279c93f", x"8b93b0dd10f7e0c0", x"dd79e89943e76f7c", x"433f7ef9c6b8e685", x"7310d10a6c6f5e54", x"d33dfadad88f6802");
            when 25281796 => data <= (x"76e2145919caef82", x"1de547c1354fc14a", x"bcfa6ad76fa9711b", x"b4daa2dfb611aeb6", x"923f16b4ec4822ce", x"b97f00d3381900af", x"1a94f9761438adb4", x"390b8b3c1b00af50");
            when 8742031 => data <= (x"db5090f6b871e474", x"994acfc5ed290c95", x"c3b74c1eeba161e0", x"39ac18463747e11d", x"3b7234e9ab61283d", x"2932075cbe67956a", x"99dfbbf76e8f6eef", x"9ae3854dc79ad38d");
            when 21316168 => data <= (x"b8c0b6133b7bcb3a", x"bc52ea8fa9b2efc6", x"c2eabaa34eb17d09", x"eae82fd15d94dd3a", x"fb2d309e5a621921", x"fed2ba312f3553fb", x"555710d08809a202", x"0aa6b95c36630297");
            when 29545730 => data <= (x"40821be9ed6e0e07", x"d05364ad8c218a51", x"acdc7790c9577291", x"157dbee4e204eaa0", x"5355d6d59dc11d0d", x"798d2a116b64a24e", x"f4c85ac7951235ad", x"5f97f15b4edad16f");
            when 8795235 => data <= (x"bd23ab8c3a40dfc5", x"e435207792b1bb94", x"011099b31795b547", x"4b83383b4d83d754", x"2a888fe44d968e30", x"f4ec4c2e5727363e", x"ea5092bf6a240f53", x"9cb9ade05b105547");
            when 23249837 => data <= (x"a1b2c2cb4999ab33", x"c9fcb3ab0a1719ef", x"4393c80a452e4262", x"9dc1bfe3e4971427", x"93dff3ba0de3572b", x"47246d7d1f2a6846", x"3bc4b9f7aeab3f7b", x"5ae27f2a99def398");
            when 29946837 => data <= (x"2b890b3bdf7a1232", x"1096e710e78dcaba", x"42c2d22ea8c9a93f", x"afd20909762e98ee", x"16f39c256e7f3c5c", x"36bff58a0fd16ca3", x"2b259f840ee4e6dd", x"e89ac955889d9370");
            when 2885303 => data <= (x"b6867e7c959a30e6", x"f456305eea5edd55", x"b0c53a6154232933", x"9531881e6d8ae2c3", x"976f2c644a9368bc", x"e647272290dcb894", x"0b6dfb053b29aada", x"c1a9a9eed2088e02");
            when 21383978 => data <= (x"8b2029fe79ab5751", x"4a3f511d2d4dae0b", x"c01cd035a5db1b03", x"a810c4c3b72f5679", x"7e3553ea4e02cd34", x"e87ec0e93aa4efe8", x"b1dc75c19be0cfb9", x"4773246f45396e72");
            when 3127101 => data <= (x"1821b3568f57b01b", x"4981df80f5b9ad2b", x"7aeb008a9236cf4b", x"6215d9cbb2d5c4d5", x"0404e26aee9ea48a", x"622690bc6f7efb1f", x"bfb476f48c222a50", x"c5426b7221adae5e");
            when 3424214 => data <= (x"7254a0745e79061e", x"c0d9ff36cda4e7d1", x"776b1e4411890e32", x"5cb1d7c4bc91e689", x"95b6a6b6bf4880ad", x"b1ed994579954888", x"44a1b0e5c4e45bc4", x"e7176aedd9e4bdb5");
            when 14731957 => data <= (x"10e6262cae422f2e", x"f1bda84d49311166", x"c07778815d4b1b89", x"b7e781c903abdce5", x"13b6b9ef183371f7", x"c5b70da04ddca91b", x"10bd6588c7ee5f63", x"8dd2b92106a7a120");
            when 21748008 => data <= (x"2b49ee28515379ee", x"4bc750fb8bb05957", x"30595bde796b4a19", x"00371c17bd3c60cf", x"34065d9f21ae76d5", x"141361a3efde9d93", x"5fa403c494fc4ced", x"8716b6809724b7e4");
            when 29098175 => data <= (x"fe029c8f9ce1872b", x"ab572e6220c40cef", x"c30703feca955600", x"990233bed7d7b33e", x"e226fca56cb3b373", x"91cde0c7591f7733", x"1f29bc9c67e1571d", x"d0a712bce48ff3a0");
            when 27577434 => data <= (x"e65947aef476e38a", x"35b402bed468fecb", x"e558ed8b7034d874", x"f5460c08e809cea5", x"1a76ffbd6a1c093d", x"38da78fa58beffff", x"bfc40d6181cdb151", x"1c4001535924a5f6");
            when 33827778 => data <= (x"a11443b75df1fb6d", x"c1b5acc189651723", x"018b252b4cce2772", x"5ac5ca8fe5bbedd5", x"6e79babb9bccd465", x"241bad643a17d5d3", x"9badc64024c91a2d", x"f9d418b4c892e777");
            when 13948538 => data <= (x"bfbc568cccfe4622", x"f64fce027ef834e7", x"9961e8d183fcea7d", x"206f94dedcfca16c", x"08b0087e46cf81b8", x"f4701aa374194f4c", x"cf39edc78c4492c8", x"0cf435439ed5f0e2");
            when 7598325 => data <= (x"919d1f7f64e03016", x"66c49ec9f416ac5c", x"e54c5f1289b397ec", x"8aad7f5f63f43e36", x"c987c354b35910e0", x"371257003dc6cbe9", x"ee28115550b21b84", x"9f76fdce1fe6e379");
            when 16948045 => data <= (x"c17e905453d4782f", x"c000d682577daf3f", x"c0771dd5125936e5", x"6d942d3b5642438f", x"f393b3d9e5179593", x"73b06480cbfef416", x"8d828c451317c644", x"c6b08b6167dc6f05");
            when 22985938 => data <= (x"913fe62f5a2c6a0f", x"df83448b59a46dae", x"2fd7c6305c28d094", x"d07e51a0c55e8689", x"80315915c1e0dc97", x"498b04520b3058cc", x"32654841f1e67581", x"d0069b9bf7af41b6");
            when 29065408 => data <= (x"1e9c8fd5d1c2de5b", x"131897fba584297f", x"03b64aa05caea301", x"7d8fb39ac7aed14e", x"d110a351589c6f7b", x"3c49947baf5b6ff9", x"b47717ad4b0e168a", x"49b4a2fa44771a20");
            when 1660169 => data <= (x"67f8ea2f9a297709", x"be03d252111dcf3e", x"de4e07cffa904d46", x"d8213e8b161b34ed", x"41f3d4c238d4fe1a", x"6a196ce935f9392c", x"01581754d2286a95", x"d56ba59eaf05db9c");
            when 26056635 => data <= (x"f34199368e0456ce", x"79f2bb198f9e6a25", x"5090b5b232635b62", x"3a971fa6427a8e72", x"688bd319475d420c", x"2b3b169c1e8c3edd", x"c09dc999b14d44b1", x"5364d177559c0a29");
            when 9265273 => data <= (x"180ba160f60a5237", x"04fb1f88332cfe33", x"2af43577f453034c", x"377c4e9550f2e427", x"837ab3c027a20d79", x"8b62b4a7c70f5823", x"4c2c2645b44f47ab", x"e14b7eff3a46f9d5");
            when 20379023 => data <= (x"c7edc6738de13556", x"8b6b4001d60e50a1", x"9d7bbf9de53409d9", x"272f918ed526117e", x"3293a579e870b4ce", x"d69b21dd3ed17bee", x"45c7ffdc1bbc8e2e", x"0d5b83da4b41a2ef");
            when 21192244 => data <= (x"3696f2ae2757d742", x"df6ac7958c4fc331", x"dec55f1efcee0481", x"283b1b5abbb092c6", x"1297d9123fd6c5d7", x"3cab48770cb2dce3", x"360c98ae87aaf354", x"f9d960864b92cb66");
            when 25265252 => data <= (x"9c90e97740d57c1f", x"296a78414d6c2afd", x"4643c4038268c772", x"ba2a5f3c04f003ae", x"1452df55a073c1d7", x"7a23d58f9c9278cc", x"b7f73ec16e6185db", x"a53ac79362b2fe15");
            when 14062819 => data <= (x"e028a1a36e2e4ceb", x"49c5e4bc897fbb13", x"907eec6655a4230d", x"14c73a67bbe350a3", x"be7832c0cb25bef9", x"aaf6f7a183944ac1", x"2e95839f8a170f53", x"29a5d4f79ebc5666");
            when 32971273 => data <= (x"49b23c682913f88c", x"604211397fa5c1ea", x"fc2f6928d77fd15d", x"6e3f67945607b3bb", x"5849c21fb640c42a", x"abb25ad01933dee7", x"f72e82ee285c8162", x"562398161e58f403");
            when 4175271 => data <= (x"4cb08ba1e66fc927", x"2bf9401ad5216c8c", x"b4dafd29b6a3a1b0", x"b740cf867a12509a", x"b5419b0a6a5aa4c4", x"10a4808eb72746ad", x"a42e00c4306a4d28", x"a105496132de9a65");
            when 26713435 => data <= (x"0d3264eec96e2331", x"ca5e37ed2f44845e", x"a9b850604f538b35", x"ff6f721ca536d896", x"a8e1f0006937ab2f", x"ed2e837d3f08d55c", x"fab74e833f8feed3", x"b2c5aa618248eeb2");
            when 24235671 => data <= (x"a9f67bccc975a681", x"7d3900277c824349", x"a204a49df5ce9982", x"c10e888ccb44984b", x"b5d60a33a574618c", x"6607fa8c049f3b80", x"a0729f1d610d063e", x"f249b7c3b3d8af96");
            when 9161127 => data <= (x"5342546c8a8df4ef", x"8e7b87a2c417ef6a", x"3bdce3c9c32394ca", x"76eac66617561085", x"f4c0d18d52fc039b", x"65b0854a87728a2b", x"4b206b59110c2a61", x"9db7fa40bb901e21");
            when 9154019 => data <= (x"b5ee478995c34b9d", x"21f3823f0126e4d7", x"dae1285874da98d6", x"c553f9c8bf2a8cbe", x"c808bc526898bf3c", x"d65e9c6b8c3ee189", x"786b7337bce59759", x"afff74ebb9ca2085");
            when 29826431 => data <= (x"54f5d4a2f6a24281", x"56a2844d1b111410", x"6c5bf6779796c8dd", x"58d10062a7f571a4", x"28edbc72782e73af", x"4e86fdff3acfa361", x"803d70f3c11b51cb", x"8515689e9f56a4a7");
            when 9531420 => data <= (x"87fea6e4f252ce66", x"5233e0b8338f4afe", x"f955a79c305367cb", x"4be75c4a431cc123", x"ba20ce61815f06b5", x"57d10580871a4cf4", x"398c355209b5b2d5", x"1fc1360b5f82edf0");
            when 15563613 => data <= (x"8bafd183fef0310b", x"820126349d145dc2", x"c5236c6b84f9e27c", x"c2484f1a28ca8215", x"1794262f3d0fbd23", x"e022d894ba1d6bbd", x"b7362635cf9d1359", x"0fe895afe4c9ed66");
            when 17595768 => data <= (x"02ce2289b9af6845", x"2cf2390e6ef9c166", x"57272464491399e1", x"322c6ae9407d63ae", x"6c53f5b53f86dd74", x"18eff6041a19dc99", x"bf5250d846d03df9", x"265cb1d2231dc533");
            when 24239097 => data <= (x"36d8143e084f2b6d", x"fa09ba2f5dddbb47", x"f01008b6e9855f67", x"733638f678ede1b7", x"ab9730f0a899f4d5", x"4254975a96b04e00", x"7ba97c173889171f", x"d024c19c54e3cee0");
            when 14979348 => data <= (x"9e631fcfa41755f0", x"e4e098296240f742", x"b95c2a13f5e6987d", x"44140d36e24c9b25", x"d666dd95840e340a", x"73197304b14861d5", x"6576b45542bae741", x"0752caeadd53345c");
            when 13155134 => data <= (x"6ad439e7f58f9746", x"118cc16dfd16aae7", x"f0d6d61ed4df276d", x"6e1d37da6b16f714", x"1fd1c2e9ac2a9e79", x"6eaf315e149a2757", x"9275a96ec5a3ec0a", x"8dd0d157d1e39ed5");
            when 23125022 => data <= (x"ff1e897b17b7ac46", x"b174f60d1e019e69", x"c98826dbcc6a5edc", x"8804884709d1573a", x"a356fa7681054bdb", x"b30e13b9b3160b98", x"96d5693ee26ef4e7", x"49db8ccecac490d0");
            when 31326107 => data <= (x"fec6aaf787c06e8a", x"c61d9b42eb25e557", x"3df04145ab06a1f7", x"c2627b2156ca0230", x"4c1fb6136b53a0d1", x"8cf78edb2262b69f", x"8ced83bba9ddb88d", x"25bfbaf808424619");
            when 29876795 => data <= (x"d82855b5abf04181", x"75d62b15b14aae0c", x"cdd3de60903263d3", x"e896cffe3963564e", x"a98685a8707a3f70", x"cd5a61e3640f546e", x"7a04ce27b7ebb483", x"4e0a14e399031ec5");
            when 31256383 => data <= (x"0f2fbb2676fd34f1", x"0045733dbceb763a", x"1f217befad918f1f", x"84d08ea684f9fc5a", x"e29ab4fee1237c9b", x"34dc0b728e3438fd", x"a61a0f6fb578b156", x"b88480bc79339819");
            when 31874759 => data <= (x"9bf1dd598d42760b", x"2aa7a3a2e1d9d28e", x"27c9706188ee30e3", x"c0fbb84b338bd2ba", x"93d4c199c070eb1b", x"fc93b5bfa5eb2b5c", x"691ec6250b796341", x"fbd2a959b1e88538");
            when 17833874 => data <= (x"56e2068c2ef4e009", x"94ac9830c81bdc33", x"60349b3336980f76", x"7dafcf6efe4b43e0", x"0d463ff3769e28da", x"22c0f4c0c0d3a3b1", x"54704b8eb280bcb3", x"7915edee2e1edaed");
            when 11058265 => data <= (x"a1e7b2b6675c0bb7", x"3af7c6913abd000e", x"b0278cb1423ea83e", x"fa10c6d6583bebe0", x"0e75071b77022366", x"edab290d49abb728", x"24b2786199fb13bd", x"731dcf0eb79e6f7c");
            when 1971125 => data <= (x"82f958999f0d8557", x"ef802ab5b3c09c75", x"dfe69031e2184c89", x"5de85da8197a329a", x"59e4a620105cddd5", x"4e94a4c4f6b942da", x"26e5b579474a685b", x"6abd702bed903433");
            when 28800024 => data <= (x"1e535d71f662ddc3", x"ecba147c027b5eb2", x"3875b0471bcc81ec", x"95666671e4d288cc", x"b74eab795c0d3d57", x"30e5acfa8392f38f", x"f2034eb902e7b924", x"9c91962ed6a9cd33");
            when 24875312 => data <= (x"fcddc6ac0d47e113", x"1ab0a637690c4a91", x"0e99ab546d0fa95a", x"83feb81e3ecb9a97", x"7d8b2dae4d866fed", x"6c091b773d57bf6c", x"e880f44794ca7e04", x"76e6648baa100d5e");
            when 3409780 => data <= (x"3be0c04f89ec0780", x"c2cb53e3604388d9", x"a3d12bda42729b0a", x"1273143a323e2e19", x"c5efa5f2b211a979", x"253e7205f5894bc4", x"84f6420200e3bb7a", x"d3a4f47e49e95f84");
            when 27064352 => data <= (x"05c8a709f2b1d6fb", x"96e7b92c9c0cd05b", x"87601780a9d922be", x"873e16c0a0352bc8", x"35b557be22f9d4f5", x"9f5c6cec11f84df0", x"3de19976c5aea6a7", x"6b66840b95c301af");
            when 4421992 => data <= (x"cc3ec9ee5b09ff77", x"fe44ca3178aa31d7", x"e4468e26e3814ba2", x"13c5a45acffb0962", x"c2981ee37865fea1", x"4aad2e320223f564", x"988a4ecee47408f6", x"bab27e6bbe051d48");
            when 2346053 => data <= (x"2cbe806c9073021e", x"8498a6c787fea0e9", x"13a6d68b66d1d4b1", x"e39428e59a606850", x"d11326f86887265d", x"0ff6a554b9e8e7d8", x"3799cc357b8241ea", x"8825cd68753d460b");
            when 28945747 => data <= (x"fca3c31a474c1460", x"d6f2c864ecfa7a59", x"b1be81c1b84d695e", x"cba9ecf7565a7d04", x"a72e3d61b0021fae", x"776be9b144307593", x"73f2b2e5baf537a7", x"c756ba22d4d0a5b3");
            when 15965733 => data <= (x"adc4121cf2685aea", x"24f13a5ea2b467a3", x"41a592572233ee98", x"869c1345bff83720", x"537e4553c62bfc83", x"1e81a704d90c1ece", x"988cf08942b87b4f", x"dbc6f0a34a39939c");
            when 10342153 => data <= (x"19b8ad7dcee05854", x"58ee5d980109dccb", x"3f8b85c9cfb1b79c", x"db44a43fc1b025a3", x"0686078d7dd9a3ee", x"e8e31591055464a0", x"608300178fd17ddc", x"a931599db01bf834");
            when 3167632 => data <= (x"a88df69707bda97c", x"72ba54117993f055", x"8b1952c59daaf4b3", x"4763e0fe3d95f90b", x"4b96d459a3428c15", x"db534bf78077a752", x"3c4306a06cb94310", x"21ce53f72d366d75");
            when 15423551 => data <= (x"95c071f9b5e3de3d", x"ba2d45237659ee8c", x"240836aa0ff2aa96", x"5f22a45cd43df4a9", x"816be38972e1e159", x"3607ca438599842b", x"9481137bbf8ade58", x"88a3a031b0805d04");
            when 32967838 => data <= (x"e4507cf8d1abd085", x"ca830c84490d250c", x"ec32131a4a672287", x"046bc68013d510f5", x"8f71da46a6368fa1", x"d7b33bb785a21881", x"e18966d6ee6e588f", x"a8aaa32c7d8875f1");
            when 22510876 => data <= (x"f1330a9b36520ff4", x"97e74b2892ab6840", x"238d2dc4bf0e8391", x"485356f796d0f68c", x"276028d4217a352a", x"5514161c6ed6e879", x"1fd068b62b7ae452", x"fdb12a1e74e53463");
            when 6216067 => data <= (x"9555c6bde49deb6e", x"93de4ec12ce1264b", x"d1586a0ac98c68e7", x"cdcd0581fdec615e", x"e8edf6600d675158", x"9f87bf29b0ffd698", x"6af0fe8cf268699c", x"215cef8c85559316");
            when 21493591 => data <= (x"dec83edb502af23a", x"c751e13c6fb075e9", x"4199ccf2aaed9c34", x"f16def409b8d1002", x"6e5d363133b1cf6c", x"e5e985cfe1527af2", x"79d418243bccdadd", x"03e5d67532cd8f79");
            when 6432999 => data <= (x"36cb10db2c488ac9", x"48f84dc03b81fa33", x"fcb8615ab681fdb8", x"34f0d4b5347cf448", x"05e2d06706888034", x"420c4181a358fd8c", x"210e9285fe51b29e", x"ad9d4b4a3e67e859");
            when 32601525 => data <= (x"7832efca7971e44c", x"075078c62610b203", x"274682c23346f310", x"49f4957b43fce0da", x"aa98c81ab7f6cb18", x"03d00cea7c67a9f6", x"a36e6816bee4fff4", x"f63555ca542c7c9d");
            when 26837863 => data <= (x"fcd13f5af379e99b", x"71bdc56994630905", x"05af2b7113bd6e27", x"4217abc6fc3f1e75", x"a987bc6055a12529", x"d7288c0b8afb3f47", x"89b4d58a31a068a0", x"07c19054be70e4eb");
            when 10302078 => data <= (x"3ef9d2f724818f9a", x"5bec9a9287f9b8f8", x"36ca6f29ea822283", x"e8bfd489d3ba312f", x"177255676e1c606e", x"980748d01b1fac68", x"cb330201ed2090a6", x"cbf5b88995fbef79");
            when 1826076 => data <= (x"3c1af80921b8c2a3", x"f07c3e046319cd0f", x"5fc04be8346ee093", x"0147621c263da594", x"579d264046b2661c", x"21b5555a8c011ec8", x"77a505e6b5e36e0f", x"0434879dc29b3a26");
            when 18451199 => data <= (x"624594a0ac5c438a", x"6643aa8817d4a209", x"7ece472854e1ad6d", x"867d131d269b5847", x"46f218c9208d4218", x"228e498e2cd030a5", x"b24477e827795701", x"f3e9319fee97df70");
            when 27292975 => data <= (x"7d3194654c26d732", x"c65e37ec4e22bdea", x"e3db046f1b5e8582", x"9aa894d22fbebe1e", x"cea71351c50f150a", x"b8d7fcecb42dc963", x"6f5c55c0f4446e6e", x"7b86beb7a8df1a13");
            when 7405633 => data <= (x"d29425a9eebb858d", x"9e8defb1da2e39d7", x"5119c31a10d0af70", x"50cb74c913efe3c3", x"2ddfe667678774ec", x"322b87e82822bae5", x"5c2ebdc9cf46b0a1", x"cf2a02cb3f797b97");
            when 31353087 => data <= (x"7d9dc244c19181ef", x"8b3eea4096209a2d", x"43a794d80bfdcfec", x"993c17c0d73e7615", x"d260cf47dd42e39f", x"4e374877efa47a17", x"b12e31b0f510844b", x"eca7fc22a47109fb");
            when 13419992 => data <= (x"b371adceb29b4476", x"a095d51414afc9a9", x"c332b10b80da50a5", x"7404fa9173545597", x"b718024467ac3d89", x"ec1a1b288b3ede2c", x"047a61ccc16c5ad2", x"303c53ef1610b7cf");
            when 15961203 => data <= (x"9524219e83228aec", x"cd1989d24d0f3b5b", x"dd22ad3fa54f996d", x"ee835bf722e36e30", x"a8b86e0c16ef5c30", x"3d6fd01ec7dfab23", x"24220ed8d05c536b", x"586b022cd9cba522");
            when 9591585 => data <= (x"76d62f13dd4235ff", x"ba7377e12d9cdc90", x"fca9fc59c97be95b", x"f379bfb033dd03ac", x"6d7b9cd5376396de", x"a22542e301223aca", x"09050b89ea783962", x"1dad92033a06187b");
            when 10850600 => data <= (x"e651f68191afb64c", x"06f779f33019310d", x"7572169ed23102cc", x"257eaa679554f184", x"3fba945108d75f7b", x"78d3eb877109da0a", x"b55bb0b9ebff168e", x"1a92107a18bdc106");
            when 20888630 => data <= (x"f541784fb6160399", x"0b93590af8f45e80", x"a3dcf3203f979cb7", x"2355cfdd3383b95f", x"0baaf2a46e986cdf", x"7811a3fd3a5f0319", x"b1fd68d2892bad25", x"f6704303215f60c9");
            when 33320666 => data <= (x"2c48df77652c02dd", x"5ffeb0a0e68ad054", x"bb7010cd34721556", x"e4e02883d8d9e299", x"00fdb45b7be4327e", x"12a9c500e83c97f0", x"f749f9b2543a4ca9", x"b0380b516981690a");
            when 15698932 => data <= (x"9024ee7074a76c24", x"9759182131d60f97", x"9c2a43f8eab886e3", x"52291ad35ab97a81", x"57a9aa91d1476d8f", x"b263604bd59509d2", x"61dfc5a0adf1be42", x"92395133edaebd59");
            when 23728509 => data <= (x"f85d24dcc9cce94a", x"ceac1174a7761c6d", x"439823807ab5738a", x"30c6dec3956d91a3", x"edf5e2674aebd389", x"6f42c0f8c34569ca", x"625ec0a2b681edf9", x"5e16fab58c0fa59a");
            when 17473659 => data <= (x"8347425a5ff74227", x"96c40be8fd2b9dca", x"9aa6180129074ac9", x"3179e100bfc88d99", x"f56b7882a91be50a", x"a60c0adf99814016", x"6f6a4913e50153f7", x"0ba7a58fd3f89039");
            when 29852339 => data <= (x"13c8e31396a4c8f7", x"ca9b23b70992ad5b", x"c64f4d3c2e7b540f", x"ffd783a61b2cc775", x"20dd9fbb750a449c", x"f0d0034c847f5019", x"62324dc16bf6b2e2", x"5cb9f6fa3968f492");
            when 3565114 => data <= (x"84475234ce80a8ea", x"b475525487f32bc5", x"5fdec8d12e4520cf", x"67def6ba9003d0e3", x"4536e324c7a48828", x"b39a00343891d36b", x"d6bbac7b79f62eaa", x"e20c99d1550b2c92");
            when 26720785 => data <= (x"9f959dc26d1703fd", x"9f625496522e5d17", x"c4a82de3f1d501dc", x"8a71382cf1fd3542", x"790aff9349472c8d", x"27b36cf23ccb1b39", x"d61e62d4dd12126e", x"e1fcf786f67fcacf");
            when 9038285 => data <= (x"011aefa86172862e", x"eb5809861055ea54", x"11014c1fcd8612dd", x"786588ec001c90b9", x"ed6dfa30bb7582fa", x"68fcefc4699e2b3d", x"9e9323067a3a0f61", x"4b3e314a75a6432d");
            when 15466337 => data <= (x"6a1d6096b1640087", x"e5dd903ffaafe8a7", x"7ebba4900ce8ea32", x"e04e68062b85de44", x"c44698b9f3e27ba3", x"1d0f0096b1800976", x"ee8c1a90df7d6481", x"a0757cfcbda30a77");
            when 3947312 => data <= (x"345208e8df688c26", x"2a3ae64c3b7466a6", x"499fdb4cce752c8c", x"4574b6a5e0d06502", x"dded17bca7c14ca0", x"ee17fd490ead676b", x"58a0361c4f12ad13", x"ce518149c61ad498");
            when 6821362 => data <= (x"baa1aded8e624890", x"ca5be0a6e3732331", x"c6c77a2dee105683", x"9eac087d4a17ee71", x"49a76d1dea4ab487", x"deba958dba7595df", x"f8220785c41d4770", x"d08800903b313562");
            when 11540140 => data <= (x"e2d1bea66a064a0e", x"c8c0723a9748c668", x"4f5d2407b098bec3", x"26bb4b7dd10daab2", x"26c0264242bbeab7", x"6ac35ab81a4f41ee", x"64387fba8e0ab365", x"a6d01a1dbc2ff7e9");
            when 3392005 => data <= (x"1b181a0ba7a72561", x"b4db2ca634fe7753", x"b4175b74cc0612a9", x"6380929cf02ba22d", x"b1428d004fe81ecf", x"238e03ce09d45bae", x"ad71ed79253cfb07", x"4897d57d2f85ebbf");
            when 15689356 => data <= (x"e7839e382da55553", x"a6711f4dd6d79da3", x"16110240f20efce3", x"a0041c5fd80ab995", x"06275517f7c0d929", x"9c381cfbc39c502f", x"cec3bcec35b331c8", x"4ad59bf23d111464");
            when 7995407 => data <= (x"39f1d07668473469", x"27350db2fe8c62f7", x"c3efa2e77d43ecd1", x"d315c4214381ea18", x"a828cb2bd6732d41", x"67adee43e7db5457", x"9606edf7cc3fe190", x"68b341490284a4ec");
            when 6881003 => data <= (x"6b10ea9d674e50b8", x"01cf1c692acd43a1", x"0ad1cc43fc5beae0", x"3cfb725c8b4082f0", x"2906a9db6d13c965", x"b497d0ea9a81758f", x"341d3797e77cdf03", x"24c3f162760cda05");
            when 33643391 => data <= (x"8a6a39d4d3b80a2d", x"1c57cf12cf327b9e", x"d9f57b577ca30ad9", x"7902431fb36bb8e9", x"3408515a76425385", x"b0c7d731ad5e3d36", x"10c8573bcbbb4220", x"8e16cb105d40cb78");
            when 24074164 => data <= (x"f3930f9bfc5f6634", x"93f2b7a3e5d2bc14", x"7711611204b10dce", x"940db2cad20f0c71", x"7e9fcf0a2159a9f1", x"7a99ad645d2fa9ba", x"15136bd0b96e1d0f", x"cfeb73d5b43a8c8f");
            when 4512648 => data <= (x"243e5459edeec1d8", x"eaccd8f4adc05517", x"5f9a4947187ce421", x"0c96c1c5f0ce0bcf", x"c73b97d5a8ce34a6", x"a7a1b66ad389025f", x"2ee42c426fb012cc", x"01f4062edec6b726");
            when 31865193 => data <= (x"3473882323045f1a", x"a59ded284b863b60", x"d2b87bcadc1f2e5a", x"1c74be561688258b", x"f4215223c224d3bf", x"dcbc5d6f0891b611", x"eff9e950335fd8bc", x"d830f393ba83fb12");
            when 24503523 => data <= (x"1d52fea545a50c5c", x"74bcac1645fb115d", x"b24b60371a4d95c2", x"5276448b4218f646", x"484301178d2b520f", x"0b52dbe4911b0479", x"55c6b995011f15bb", x"46dcf698bcfe33c1");
            when 17855027 => data <= (x"d0779eebb20d4a91", x"6a3c5a4f21068237", x"e9b1171e84f78d02", x"7361fe4c615e62bb", x"c48ba70498313884", x"33095901c9bf25b0", x"1ab72de91d0c30d5", x"f8dbde947445a070");
            when 14752592 => data <= (x"99143a7e51f125ba", x"2f857ee013b6ac1a", x"a32657dc832e320a", x"a44336c9f4ac7569", x"8c6b3e2480536753", x"c2464f18c0df040e", x"0199f2f0f117612a", x"debf14d43be00e19");
            when 7691492 => data <= (x"b0009fa0ae0cf022", x"6d3544aa1a317689", x"b512fcffa8735194", x"2d1a418d4b4031e4", x"6bdda06b3e8cfbe4", x"1f8fb413eaa3f131", x"27d3063e1b1d9a01", x"4373a66478ea5a9a");
            when 9228092 => data <= (x"43e6b17182008907", x"a42334c8d9d18eca", x"9906540a555a363e", x"ce5f89e85a8cef15", x"f0ac9b7cb45359a7", x"33b83d6c1e4f2e83", x"ca54def36551039b", x"364e5b3ac644dcf3");
            when 8267652 => data <= (x"c5f02e52e5b069f5", x"e1fada49873be917", x"866e95cf8b750655", x"35d1177a43982cc4", x"16b26b8480e3bffb", x"f58bfe2a523799a4", x"6897baeb2f0a2b69", x"57c54d1a084711da");
            when 26133499 => data <= (x"3714c00f34f76b15", x"9fe661f957ff1042", x"6714416593e4c98b", x"8ad7e8327cfd18aa", x"0f5cd88487a545c6", x"a45063fdc1424acb", x"bac938666b18cf72", x"8eb23c013af06971");
            when 22893208 => data <= (x"8b6ab4752efa1efb", x"0daa043c0af185dc", x"ec69d8da5217454f", x"7614d72fdb19a566", x"7c6352e0bd5ab380", x"b7448b263fd73236", x"dd9cae9a691e86a2", x"819504ff45fc6574");
            when 27292400 => data <= (x"7159d4c13cecb6f9", x"c91414717768c109", x"76c7dd498ecdb159", x"e05dbc526f862af4", x"7784297690e0859d", x"daaad1f9685cca36", x"ad0ecdba90f3e41c", x"24fb752eab681c37");
            when 33669949 => data <= (x"d9d654a2738c8819", x"a621b4f2d6f2721c", x"8c2febb9525be956", x"9a9498ee46213cc7", x"ba1002a810941431", x"d5b22220e5d887ce", x"53ed70d94f32aaa0", x"d23ff475cb468434");
            when 21735737 => data <= (x"15f3af0c4d7fe093", x"d15fac4cfd94867c", x"c443f9830cd79828", x"c46f3933c0496e78", x"1796a3608650bad7", x"53cae933bfcd63e5", x"8ac52d9454f964a7", x"820298c7f2e75a1d");
            when 15387615 => data <= (x"db393a3f62c39d5c", x"67eecb792461e8c1", x"82102b92a26d7ac2", x"bdbb2f3e023da6c3", x"5c98fc8be0bffcf7", x"195e1ec777d9d63f", x"7e9f0122106b8eff", x"60cefc9b36818c99");
            when 32423094 => data <= (x"2a9e1ac486327f49", x"ac8e43bf6f8e3c97", x"a4a4bcc8960a75b3", x"3e49594bdce55d36", x"2f812d59ffd2d470", x"0b1f9f5dfb98cc17", x"4bb25d25ff3cf4ee", x"2eb991ede8458f09");
            when 10013604 => data <= (x"5cb13158d4d8caa5", x"d50c16e9fee7f1e7", x"843457e49755671f", x"e133eedea354b007", x"f79f8633478f42d1", x"7af4c3090f2f9e24", x"a9f7c07ba8c2abe9", x"3100af3b327536dd");
            when 15313358 => data <= (x"a0eb287c08c24a72", x"efbf1af45b721c27", x"1423e6375e99704b", x"7aff802db2862624", x"25abec90ee537862", x"ebabf269eb5e78ac", x"36b8d05efa89e21e", x"2e0f23538a28cda8");
            when 8300105 => data <= (x"db83c0be2eb8c9e8", x"49016ceba0327e91", x"d90e24622126f084", x"7ea0002f1637d991", x"42d1fd0e318256ec", x"5973a1562995043b", x"780f9b10878f4d27", x"63a5bd28db6650cc");
            when 6462855 => data <= (x"53af2eafa254ff36", x"acce097ec2a089e9", x"2c0ba3974e6d7f74", x"760e2d1c6f98d17b", x"790fe4dd81509849", x"f36ec7a573a94cce", x"cc093dc3f0ed8e50", x"b29f096033ca4942");
            when 30152002 => data <= (x"198c0d623e7bb813", x"b6a75e2b1031f46d", x"e1c597e18b1d1001", x"385899bafe1e48c3", x"fe188fc5560bc228", x"d79348e8e85c60a5", x"b48f35f0d9095217", x"6a6655ea0561acca");
            when 15363101 => data <= (x"c3bfed04c0d22b73", x"9613b3b4f5b80619", x"ec0a6200bcfe2d20", x"80cfb63abbbb67ad", x"6fae298345eb5b60", x"95a049b023571df8", x"88fa7e5e2270f88c", x"7c8046b9acfe0eaa");
            when 22723101 => data <= (x"3a88aaa2de21a805", x"92752efddf1b69d4", x"80805574b61897d9", x"4bd84f2442f537ee", x"787a91a62cef21e0", x"39bac595c91eff67", x"99a25d1b612e0c2a", x"40f990e136bbcb88");
            when 32183485 => data <= (x"51a9252087d9e2bf", x"0d6206a1f3f9268d", x"872625eb75f10c39", x"75504d9e03020dbf", x"5b6a7da2563d49b4", x"3c25004721383b4f", x"3d5c8c831e20605f", x"80b67ecb043502bd");
            when 23277207 => data <= (x"1bc00e1ba871a649", x"6d8748cc5990692f", x"b9a8046b8331da68", x"d7ce5aba215d9e85", x"fee0ea02391ced78", x"b65c0c6d9b9344e0", x"781dc8e45de6fa27", x"6e72212937b98d2b");
            when 13894948 => data <= (x"08384df2ad82b2bd", x"986278651e6774c9", x"240954b24cece2b7", x"556cb3f31d6a7d99", x"3dd38c6ba28ec1ba", x"99ecb0c6abe0fadc", x"aaa2947e74afec66", x"5093d5d4756ee5fa");
            when 31683371 => data <= (x"a028751df4dbc556", x"27e87132a0c499f8", x"66e542993b8db272", x"00059732c3540f6e", x"b6633854f3d4f954", x"b992f5e2c068b09e", x"449d99b676325ea7", x"77643c1f40855072");
            when 1114787 => data <= (x"7dda6dad6298948d", x"45279b2215c752e6", x"57fd0559a637348d", x"518eb4b8017c6443", x"cbb45515178cd64e", x"fd81da5e26f946ea", x"7b53465617ac7e83", x"387866b9f45c4e10");
            when 22263107 => data <= (x"ca8d0a79af8f71b7", x"bee979150b32aaaa", x"82a5224601605414", x"1f188b455e4d4b59", x"63b69c961be7c13f", x"ce9add7936cf4dbe", x"40fe785abda6c827", x"7603150deaa56b4b");
            when 33259228 => data <= (x"34934421a6f5e799", x"b8b0b6565b922077", x"b296556b59d7d033", x"a1872ee3986533f9", x"ecebb8bc87634850", x"4841a821dc035891", x"de4eb449e7f43da1", x"225863211137f51a");
            when 32847117 => data <= (x"d267a88846bd5aca", x"1b9388882cab2b84", x"2de760b7f1142dc3", x"639701942bb1a2e2", x"6cf0a877f2f08bd7", x"c68084e31cb44018", x"3b8ac4553762d96c", x"6d53cd92766c8b46");
            when 8993742 => data <= (x"b2423a3ea9332ec0", x"d6b42ca63f244502", x"541c1926242fe44c", x"2bdd212188b4d2c8", x"f65179af1b7ef82b", x"90a576642479de57", x"d7594d722a49549d", x"6388f4b0c5b1403f");
            when 1034529 => data <= (x"9fb788dcc530539b", x"f98ecf6258800292", x"552870b8b20f3a3f", x"166547233a120914", x"10d84348b380e10a", x"1d81b4340ca1888e", x"e6891030007966e0", x"108adbd15062245b");
            when 15719976 => data <= (x"16e0a46421bea54f", x"d4f33f83fc8ceec4", x"1b682697e452c6ba", x"1dc54cdb0c97c3ff", x"e5c819e8654e9b07", x"a0c2c605ea47d682", x"a046cf68ff641484", x"941174f4d1066fc1");
            when 25464892 => data <= (x"523104ec32f79b24", x"8cebbd67b6fdb985", x"cdcc9e9289fd3290", x"0bf8514fc52a6b8d", x"a28a4e44b398b33b", x"f70cedc5bd1da9be", x"d3b03293b7cee893", x"f8ae4df247d9a332");
            when 24813071 => data <= (x"a05ad1b96cda17ea", x"8afcc4b8510cccaf", x"a6e6431ba85d3f15", x"c4e362791f46fe0b", x"0460e7ed2eb1e4f3", x"ef7110df973b43f3", x"639db07f10fe98ce", x"d1de4d7f99dc874b");
            when 3709870 => data <= (x"72b13090ddc8d1f1", x"08eee469e2d4ddd9", x"1917e624dc43ef17", x"7b141917dca5f0c1", x"9d61a256bc33444f", x"c1ea3f854ac03eab", x"20b136ad7f08614c", x"5d5785adf8f18bd8");
            when 2113219 => data <= (x"ebddcaf0534f984c", x"1676cf84b72c5b1c", x"340d2d4b0544e186", x"5dd50e6807d674ef", x"47514cbf5d1ac0ca", x"fcc3af5e2e3fc26d", x"15661d9fbd1cfb91", x"a80679ce48c56ca6");
            when 28995174 => data <= (x"73c658867d012b4e", x"8e4312ddf5b5d0fd", x"52f231c6ed918477", x"04c6a3c44841e8fb", x"d17d69f86c1d64e9", x"c82a65ae3f085126", x"440fc9e62e886129", x"10bf6cbd37367b7f");
            when 25618265 => data <= (x"2d1caecb37f271b8", x"c40fc57d233768d5", x"19c40a0ea293ff95", x"2714ad6e1ed0a141", x"eebd5f5c3d5a176c", x"c4ec4491c90f34d1", x"4840ed8871536f4e", x"90be51d2a957167c");
            when 10065804 => data <= (x"7af7adf30cf9fd73", x"4b1838d220f7f1e1", x"de47d4c2fd83b8f0", x"0059c6e3b06d17a0", x"ff4c8baed1215a27", x"a8de51ba55eaf206", x"da838ef83926150d", x"04647d7702cbaabf");
            when 28608045 => data <= (x"98c9e4588c07a474", x"9dc27bc92f99f54e", x"e916a2ba6d3fc316", x"0bd33f6ca3dd9467", x"4342c88d0221b677", x"0c01029ab6d4f4b8", x"cf32858575b2a4ba", x"38af681e660569b0");
            when 19138269 => data <= (x"6d10950dd1e009f8", x"71c6e5c6d48bc786", x"3af1135bbf8c1a9a", x"c983ae8d845d7cde", x"02ad32ecb3fc702c", x"fd568eb749b73426", x"c00083efa690e5ec", x"911ed416476427e9");
            when 5667207 => data <= (x"5031e6780521d951", x"58d230d96b7f92b5", x"1da62dbb482b5dab", x"50f30b13a62b94ad", x"67ac01dea962d4b8", x"2e40b1facc235123", x"3c256a15307b06d9", x"53a0b07ae627d5c0");
            when 15970691 => data <= (x"7f72791fe7dede0f", x"6211067cbaa41cbb", x"31b073bc5746742e", x"56500d2e61ac3bc4", x"706e9da0c49d6251", x"1e563be24bf235f4", x"999c0087fc94640b", x"328790b0e35205ed");
            when 21626339 => data <= (x"43f1dea5a41ae780", x"74fc7f00a39fc628", x"a64f8520b67d0829", x"1109c88c12d6f7d2", x"eff761f5078fb6bd", x"d7cdf99f1c25248a", x"8a8444d5718cbc56", x"e0f7381c05907ee4");
            when 9077485 => data <= (x"af346f60886c2e74", x"882be9a5d296a387", x"36d1032cf1460e55", x"e72d28b640d3f144", x"871eb4950c7a045e", x"6c3d1ec210fa674e", x"f07df8ad8c26fcaa", x"c8dd084e1bea8bd5");
            when 22571911 => data <= (x"664760cec3303f0a", x"1a3ce1e533f374c9", x"27f505f54946fe92", x"0f610c242b113214", x"6165962201543674", x"3609abfdf95d0cca", x"c2778c6566b9bcc1", x"562ba265e48e59f1");
            when 27015297 => data <= (x"0d6ae8f0b58c894b", x"12e29d4106c45820", x"f56e7301f13b857c", x"437211b549ebaaa4", x"2fb2de029765029d", x"463c362caa3858be", x"df19c49df2d9da0a", x"aa88a57ed3987086");
            when 9985112 => data <= (x"d9c64fe6f2fd4388", x"205417a8c58da6c8", x"d6657a0ebda01b5c", x"6b3a50c144c05fea", x"2f541eded91460f2", x"2b1d5542c096570d", x"61a1c3a7b9b048ae", x"4f31534fe0668842");
            when 6797746 => data <= (x"f3eeb8379e77bd5a", x"752e502a844a3c11", x"75015d97e8f22320", x"043c738022b11761", x"1eec22ecf5961e2b", x"e58d28bff70e8325", x"56148da525fe7aaf", x"7dd3df0224bbbdc6");
            when 1521450 => data <= (x"05b570587cab6c1f", x"7e878cde12821c04", x"32d2d432690b2c38", x"41fe2997e3006d00", x"41475ac5f88070cd", x"a8ad257918a0b17e", x"754141692b0556b2", x"61d6d431aabd156d");
            when 20745406 => data <= (x"a7483c11da3dd5d8", x"830143fe58b94967", x"b6d96b62124a983d", x"f8c57839601382d3", x"0a520d7dd3835575", x"528052b3a0565f41", x"ef8cb011a90de1bc", x"8abc383cd7e58ba0");
            when 21972662 => data <= (x"32446d46ecfd8511", x"356d51dc3e05136b", x"5c9c579473fe3463", x"eaa6c512384b95ae", x"a1bf88e8e9a79183", x"753f9df82ec577f3", x"e3ffa2129b398254", x"8f33ef194465d0d7");
            when 16670325 => data <= (x"c17fbd65d3880941", x"dd2c5ba3e8086990", x"f700b210bd7eca1d", x"07eda4ff3b02ad41", x"e2cb1ce357a9c1f5", x"b13f6a4d8cd0af4c", x"8ddf6653432821cf", x"df5dfde23203fc5f");
            when 22586731 => data <= (x"3933f463ba92e1ca", x"b15bc4cea99962f2", x"420e7428675a79db", x"49f1b16a153ce6b8", x"2b6b1c0135484c63", x"056e8f571f0e8ec8", x"ce2547539e68be57", x"378eaf1e0fbd642c");
            when 6276761 => data <= (x"65e0ed22460b1ebe", x"fb34277cd5558cd1", x"86019bb6e0867c9f", x"8e406aeb891d7f69", x"b1befc5a50ad4e6f", x"0120a0f19a758d1a", x"a6d66ef32ab06bbf", x"09048bb9cce79c75");
            when 27288339 => data <= (x"6df27f893c9af406", x"a6fffcd3bcad44e2", x"5315870f80123080", x"a82d6dad8f29b2ad", x"baf2185126f7d9b1", x"884465a14cf1e4de", x"1435fab515b52a56", x"847a81d004157b3e");
            when 486471 => data <= (x"fce0017966d898d4", x"8fc09267bedd10f8", x"6ec3c62bd9ebec40", x"06c09098b3494efe", x"4dad4fcf7528170a", x"3ee4d8951af8702c", x"ddc12f35e2a405ff", x"5f48c26379616bc8");
            when 5827771 => data <= (x"bae280cdcb743022", x"c864ad499dc74b8b", x"389efd94f4231f8f", x"17dfea8e5d747d25", x"09bd2983c060ea94", x"25411e82d323c285", x"1ce98ae7def80d95", x"060e108b151feb94");
            when 31993837 => data <= (x"8cb39d65cad08923", x"029d4eaa5e33ae62", x"c59b8018519799cd", x"5603097fb59f9ba8", x"f9bde406af1c4c46", x"2df43aa86339ba3e", x"29284fee769688f0", x"5d0773a3d3d7e7da");
            when 23922218 => data <= (x"d08a0b28669f0861", x"a30e6663bedd0198", x"02cf1763bb7c7c6b", x"f3bf2d13a18d5373", x"73a46b19fd63e395", x"daa68915e518a1eb", x"6f9f5239cfcbcd9c", x"f67ef3c77d119e2b");
            when 13474770 => data <= (x"3b209b9f915a1767", x"d768c55a3c6e91d7", x"eae488295ba8f5c8", x"47e1c4df305b9827", x"a200bee113f6ad4f", x"e62a23498932eab8", x"1df7a8657167cfd6", x"6e1e2898d48ce99b");
            when 32025699 => data <= (x"51a354e9deb824f5", x"0839b6c73a4a2c2e", x"b6d1742886d0915b", x"5973e431b2cb05c7", x"daea16eb7c9b34ff", x"933392c837d33159", x"e51dc6ecf693b30f", x"933f8d480580e1c1");
            when 10004258 => data <= (x"d8dabaa649830d4f", x"a060914afa57f6cf", x"3956c9551c36b51c", x"e0aa448701bf250f", x"57090db7673cd009", x"e74fc3f2ed02817a", x"45f044e0e5cfe7da", x"e9bbb9f92c26703e");
            when 33612935 => data <= (x"8a2bf72b6eea2fe0", x"8ed2344c888e8ff8", x"1af84a610477381e", x"3860ab20065798ef", x"fcaaee79183c02ba", x"e9f4c6a04060d9ba", x"b8ff08f23fe340f0", x"3a3f3bb62f6f82bc");
            when 5059349 => data <= (x"351090ba820499ba", x"4fc2839a9768c4da", x"c0b1a1039e9de42e", x"7c44a327e5cc5911", x"2177cc3b81fb1538", x"7e8ca321842e78c2", x"05a04978877e9d5d", x"6b9cfaeb7721124b");
            when 2411680 => data <= (x"d2c241ad05df822d", x"bcf47bb11ca28648", x"77c35e430bf0f6be", x"d25e6cfbc4f61f2d", x"aa8013669f6bd303", x"8f8ea9f293ec4d54", x"6177831cbf08765d", x"ed5311b90a6c1955");
            when 22779932 => data <= (x"e797a931f7714f88", x"653d47b69cc89b2f", x"00c3d07a0626cc7b", x"9d92c1248d443920", x"84d916b3b0ce881b", x"298d40750a1c74bd", x"732c8da3dc2b7d18", x"fb30249558ec0493");
            when 10133859 => data <= (x"2c787bfb11f9e190", x"b2e38fbe3dea7d78", x"0aa8c30b09bd1d49", x"f2d3103802cb5a0c", x"4436c145b4ba0a89", x"4a650f79de6540b7", x"7696996a2245465c", x"4de74a5f7c9f7c81");
            when 25240152 => data <= (x"798f2fbcedbd16fa", x"23cc1bd9c2548564", x"95d0735a2539ad92", x"bb46d7f9618fbd69", x"254c359b1ff99ee9", x"16bb7239496137ad", x"bc0c7a71a7b9c09f", x"1a5030b6c6f09058");
            when 32723438 => data <= (x"957766ddb14a5056", x"e5dbca31deb526ab", x"0be7088e585a5e02", x"66bc27e6daf02f96", x"f257cd8d47f5ab11", x"d197dacebd86c9e3", x"7f60784e9abb0d9d", x"32ba5e2b8c6a970d");
            when 2477503 => data <= (x"79dcac4b1996ae96", x"16324de8eecc40d4", x"14bf0adae9e73b23", x"fa04695694bee449", x"5fd78b37c9fa353f", x"9069a39ad1f83ada", x"ffe4f2e3f0817f1f", x"780d97de302175a8");
            when 13775751 => data <= (x"57b7abf584d02d97", x"931261266eed0f2e", x"230e0fd070727d3e", x"4a4cd154ea0f641f", x"cc5535c06c7f82d1", x"2ba93801a6253acc", x"e84188d8541709e8", x"ebb3d121d35d5519");
            when 30730193 => data <= (x"4d7ffbe5bd05395f", x"75f12c1966bb551a", x"0664fa3a8641b38f", x"d0b2cdc02c4e49b3", x"2e584163b073ab6d", x"462e74bf4eb78c68", x"878df7a4d9a957f9", x"f02150cc025e7496");
            when 23371459 => data <= (x"cbc9de03175f2857", x"f8279f7676e4eef5", x"608bc67ea001f7c5", x"2578a681058abf8f", x"5bb319fc6ba11d75", x"06ec825464628c7e", x"ad8a67c36ef0ea2c", x"02c64732d1e9c530");
            when 33004849 => data <= (x"f5efc9ff37fbceb3", x"8e656289c4e61283", x"96130216fb1e1c02", x"d266717669bdcd21", x"21e67e72e44b4680", x"dd778c73d5c9dce6", x"f55efcbbb8eca290", x"fc6c60c32c1498d9");
            when 29409441 => data <= (x"e0e6adfd704c8145", x"6c37552aa8275581", x"f9a669ba23c3b009", x"4b65e38eb9df8c55", x"f1dd4eebadc44ffa", x"ca8245b0ea6861b5", x"a5860ae3dae490f2", x"259fdc5e7305c60f");
            when 9870761 => data <= (x"a3fbb261be458ea6", x"9d83b0300bb2fcea", x"fdb4ec240de57114", x"562be078bbfe8d7d", x"64d229f0035a0d30", x"81fb5b7cce556250", x"4cd74c3a3db7c128", x"bededdb938566736");
            when 4580131 => data <= (x"75a0080731163f93", x"ba5ef84cdd602cf6", x"b0a64843b11d5b6d", x"99862608b81847a1", x"a43a8d0ac1d84e13", x"1e8866f866d9c4bc", x"13b98eaf414aadb6", x"bcb54f1530b5e18a");
            when 17847969 => data <= (x"9b598c5854f2c34f", x"f5dada57daad339b", x"56a738abd27edd80", x"22406eb35d7e31c7", x"5da7a8be36c2914d", x"298a26f465d10185", x"563872db83aea863", x"ef50e00159b6ea33");
            when 22601524 => data <= (x"f8a24252c89d47ff", x"54fc5f1aa6c03083", x"eafbb40ea529bd1a", x"44fe1101ccdad9ec", x"3b04037103067703", x"2a308b659445e974", x"255e6f31d7e0807d", x"eb52a20f30e80448");
            when 6626497 => data <= (x"4217754508adf92f", x"d7dc42f0de0ded3c", x"6ead0fddf05ccbb7", x"5d0ff1068340b4ed", x"efef819ded16d029", x"36ebf34fa976e263", x"4dae0a4756f761db", x"53f4098363ed387b");
            when 4952203 => data <= (x"d55610a39517923b", x"2be818aa347b7e8b", x"a72a5fd0483866bc", x"62daa9ffd4ed5bb4", x"80cd3fca052428ef", x"a040753152e320a4", x"d62f8cd774e0bbb8", x"7138b094871adda7");
            when 6783999 => data <= (x"e84173dd477ab856", x"37564af1579efe66", x"bc051d879b237636", x"c9e97aab1fcde9b6", x"608e7d08219f9505", x"81b217323e706a45", x"ee5ab8aa5b294cc1", x"d667e06d99d5fe4e");
            when 3305584 => data <= (x"3798c2f343678eca", x"2e09ab38f03df827", x"20bc313122490fe1", x"aef36b7fbb57a129", x"79d1fc26cc146bbc", x"48289466e30cca2a", x"0fa72f72feb3588e", x"80975de837461950");
            when 30708628 => data <= (x"a1eca90d10927f1c", x"fad223da5c125cc1", x"e7094740fc8e7826", x"731466b3db50813d", x"9b929b75d027eebc", x"349398886257d438", x"8251e61c31bcd2f3", x"e50e968e9880902b");
            when 23893176 => data <= (x"184617838ce4d6e7", x"e9386829ab490d27", x"99ab553dcd8a9d54", x"0cb91a06ce9f934f", x"daaeae49768f0a4e", x"51ae2d43a20e4099", x"4e01bb2a4609755f", x"b0562be5fa166898");
            when 5740517 => data <= (x"67be7ad8bb6f869e", x"b76486f115650373", x"2ff9467ebbdfc2e3", x"cdc4a6929495d910", x"eaa5795d6d72ebe4", x"5caa328594788a7c", x"a26e69005c082ab1", x"059080cb2f88b01b");
            when 14628031 => data <= (x"ef4e03041e251383", x"de6341359ccf7abd", x"07d878f365667c85", x"7963166e54c0ad2c", x"a534e3e1309b3ac3", x"d741ff6b736f85fa", x"d0cceeb0dd708abb", x"b834ebdc87b6d75f");
            when 21937689 => data <= (x"cfa50d7adc9218a4", x"416a88bcb143a6da", x"1ec40e4705c084f0", x"da94b1e25cbd8c94", x"0405c29e9acdc4e4", x"73539489ad17ddc6", x"30fc35f12d2f7148", x"317ce471bc83990f");
            when 6588525 => data <= (x"1ce24f2c4ee2555f", x"254ef0e472e9de3f", x"b46cf57fd75e8305", x"bf0cdda38bdfff85", x"0ab7dfcbeb681098", x"cdd7d7570b39bb69", x"a9ee58517e1f5d42", x"f8545f675174509b");
            when 769392 => data <= (x"49062cb5c3903b2c", x"6f253c295d41ea3c", x"70f3afb05b900fc8", x"db7d0a4ff7acda48", x"dc43348477c4a16f", x"044e9d136941e121", x"235a4e013c898c08", x"4fc81aebbc6e2649");
            when 14149123 => data <= (x"663d76fea46a1d36", x"cde984886816345a", x"f23d5e175f8b3e60", x"568b8aabddf1dd2f", x"b6a5bef9a6e6f69f", x"b047060c77c369fb", x"0c577fb5951b091f", x"8543e2a6a86c7450");
            when 13142777 => data <= (x"3cd7b76238bb39ee", x"3e252d2ce22df0ec", x"439a64a2a5760712", x"ec0b44a8900040f4", x"7a8e099f93d4373d", x"8bb81437258a5341", x"18d176dc245fe8d4", x"585df6b3e58ab0ae");
            when 32015885 => data <= (x"e838871fcd0b8fba", x"f3e295613900bcb2", x"1938c121707d4f2d", x"1d1294c49883743b", x"772e556cd588acd0", x"8fb7a57036fc823f", x"45003731a1e65596", x"8f9384304f409def");
            when 22150033 => data <= (x"5e2be619d1f4b612", x"58696aa11ac4fe1f", x"a3ec707ee8458c4c", x"4e7549ec3e8a8f35", x"cb35562282817e46", x"89ba6876ef6a029f", x"674ceec0935c2830", x"3234a9d7f69ac0ea");
            when 11047734 => data <= (x"ad4e42536edf1f3c", x"67c91517ef86248b", x"5758b333f1d95d15", x"72f932279c310d37", x"5237adc83a55f8e1", x"e15f7fbf73fc50e2", x"7fc1b2fe89e00f7d", x"8c9f3d3e6df52f58");
            when 27900593 => data <= (x"d1bebbccd7c5a8a4", x"b92c5f90987696cc", x"b71996f462eefcad", x"9e3a4fea33acd825", x"699cbfcf0c2e79e6", x"4f9e1fe6f70565e1", x"06203170d86180f4", x"227d56146e20276e");
            when 13217722 => data <= (x"4a7a98a6c773a8eb", x"e08261125a0c8305", x"ff0a10c14fff6271", x"df4d3bd9ea339ba1", x"9ea6a794b5f90b4f", x"8433bacb75a6cf2a", x"2f863b780342c04f", x"26efb8d6e46d5f01");
            when 19640449 => data <= (x"94e542d2e2a04a05", x"b72fc5d276a0f3c0", x"38f7bccb224c7bf8", x"fc520832ef5d0a05", x"6198ef0550f24108", x"f1059c0bff190a25", x"5936c9dc960579d1", x"33e09be381069b17");
            when 1874845 => data <= (x"f97940f844d64de6", x"afd823897028e765", x"1a7088e0bb999838", x"08d07de060291045", x"9d1f96292fe57bc7", x"bd0f7c8d5a4cd5c7", x"ca5a382037cc87db", x"4a21d84402521b7a");
            when 8751516 => data <= (x"2a0af52d051eb081", x"14d5e0900cb7e34e", x"852cf6df4426409e", x"03f08670021daae0", x"fc67d8d71ef84ef0", x"62fdee54e1354251", x"3e46c52a1d2affd5", x"39c13707c76613c8");
            when 21373137 => data <= (x"bdfca49680d67b2b", x"aecee7c706963cc2", x"28ba6b6f9dceb0bb", x"e2b763679103c001", x"001b5b5f2d3c63f9", x"7459230eb420d125", x"29f666a3a36c783c", x"f20cfe23e615d537");
            when 10062680 => data <= (x"1b80bce48e2007a7", x"c63bf3cda30bff35", x"d2c8200cf550adf3", x"781e1cc30d029c8e", x"03159066d23be4d4", x"67febd0a43e94ddf", x"e4898d24eafd125a", x"75f0bfd33c2b45dd");
            when 25029379 => data <= (x"0059237036b071db", x"b598f8cea5b61c2f", x"9262ea50eef0c119", x"2d0d87ab6fff0d12", x"8916610242dc44d3", x"31d9f2ca1c94d313", x"1d0386d897926ce6", x"d9e921b33ea576ac");
            when 26586489 => data <= (x"ac038c107b662ccb", x"15eb48912b4c8428", x"d3baa55ef6bf57b7", x"3dad72fe4dfc8cb6", x"ae8c302c357ceb33", x"bfae52daac3a1ad0", x"fd6a0fab4f14c450", x"ccd24a195062c8e7");
            when 14781750 => data <= (x"ba7c1cf7a6278a5d", x"b04d4e2686103166", x"80d3f96bfb79a437", x"1baa04a083c91693", x"91c1d7537de2ab95", x"d0892b4d5d6e3862", x"ff8dd76c22c24392", x"e45c99439ef3992d");
            when 11704790 => data <= (x"f17dd18c70919b05", x"a53ed5c32257b256", x"2157aa1364b91295", x"43b25211870ce1af", x"3eb8872d83928756", x"b025673d201154c8", x"72604eeab1f5d725", x"cb4c8142a4a831a9");
            when 5194993 => data <= (x"cbd4fa22045f394d", x"8da486860865c042", x"607e9ad86231eacc", x"527ebc4c7d3146c9", x"c34f3dcb44f513e0", x"b31885bc1625e947", x"356d0dbc074be3af", x"565d13bba0305a34");
            when 15898541 => data <= (x"2a5241da368daae8", x"e6a947431a274f04", x"9529ac821768558c", x"1bf16bf2071505a8", x"91aebcb735bd02b4", x"efedeb264cd7ba4a", x"dff61362a2eadd7a", x"596154c7341223ff");
            when 33666967 => data <= (x"133680a9788462b3", x"fbed5c24c9f8c1c3", x"190057251f30d2c3", x"00c8641afa5b4047", x"a0635a3760b82e4f", x"4ccbd2bf3fa36f94", x"a4da3ea105622487", x"646d13942ed2c684");
            when 18457202 => data <= (x"bc3f7853989fe063", x"59a723cc0a10add9", x"ee6798b9dfee583e", x"f317dd1cb2f4c07a", x"06882f3a3f686811", x"039d08f8386189e3", x"900c119a178a0b72", x"c96e940008035083");
            when 1904491 => data <= (x"1485637ad155872b", x"8c72b224cc5a18fb", x"7fd0e57a423cf6f8", x"e2a24d432853370f", x"51cb3fdba196a69e", x"e36edfe2834f4802", x"12ea80400a6b8a3b", x"66bbeb822b89e238");
            when 29372703 => data <= (x"5f537e07edda8805", x"737e27de3e0cde05", x"995121b0858567c1", x"2393f909f4f9f6ad", x"e1110936ecc43a3b", x"85e75843a0b728c1", x"0fac1ad69814e012", x"e4a675367d4a636e");
            when 19070117 => data <= (x"c9ae0fa99525d0f6", x"57722900337472ac", x"5b3c0f640ceee0ea", x"291c375dd8275c42", x"c6444e180aa80fea", x"e925fc3c2a3103c4", x"414b577610221c0f", x"49e6ede654406dc2");
            when 19103065 => data <= (x"e924da2522b999e7", x"e5d850966eb73288", x"c4639f9987028838", x"e8eb1f17fc38ee0c", x"134f64a08ea5fa37", x"4bbddbbf06d12f66", x"ad9d3510ac12c154", x"564f67adba002019");
            when 25284179 => data <= (x"d5e1eb13c187fd28", x"6a88cdf0e32df24c", x"51af37f832d350d8", x"bb88f1d0f49acb94", x"15960e2b2002f136", x"a59e32d02b17da55", x"68ce88cff0841e8b", x"102097b68635c474");
            when 2254049 => data <= (x"43e394d697291110", x"031f9200b0f63382", x"0e5574e99cbb8c41", x"2b6018b54287c33a", x"f2a00ddfe4d330e4", x"819c378def3020e6", x"8146e91cbc01730c", x"2c0e9dc9942cf6cc");
            when 18245159 => data <= (x"722d889805d5ef45", x"54500f7c8e763ec6", x"58c1c0575efefdf3", x"e90e63a6080e68fd", x"8de5e3b423db2e91", x"00611d293a0cf2c3", x"0a726f4e2deb2a30", x"3e2b973c157a14f3");
            when 9911312 => data <= (x"072de8d73f68a6b8", x"7c12e075bc3d17bf", x"5f03b66ea19ccd15", x"52d1eaba5d597648", x"a57495f2f7b33410", x"6153c5d6d1b0f0e9", x"849413ede102bca4", x"5e347191216bba53");
            when 9287764 => data <= (x"384bf2008b454cf6", x"c25307ae4cd98ca8", x"9c392f085adbae4c", x"261bbc36a9d790b1", x"4243a1ca7425cd7c", x"1c2b9d944ffb0afd", x"151732e3d136a9a3", x"557b0d883db9d4c2");
            when 28934472 => data <= (x"c5c83d08bac488d9", x"e0418c03dd172019", x"609c7f15cb97d198", x"1cafe90514a12cfd", x"8b618d9911d5e5cc", x"a541f9dc4c428ae2", x"54af6c48c8889363", x"d47c0060a0523213");
            when 18704359 => data <= (x"e5cac08f9ed2f88d", x"7379b5fe7bf93f28", x"09b44f1cb944582a", x"05b21f02f4dbe963", x"69d5c9cc176406d5", x"e94364de0f030641", x"2dafe1ab03a890e7", x"ac2957ab9b01e6c9");
            when 9952121 => data <= (x"72056b05fd6527a4", x"4b0dd0f89dd8ac59", x"6ae6746c4c9ec97d", x"6bd23978745c7b7b", x"4f6bb3e45026b70d", x"d908bab8b757915b", x"402b4346c253ad51", x"3b71ae01d7ed1f23");
            when 3326149 => data <= (x"56e3e2e69513a6d2", x"222eeb0ce68c4c0c", x"97315a8c876cb4c8", x"58c3f64d3bf422df", x"97263482dbc0698b", x"ccb58b9d5cff7add", x"4fec8d92f4c0236a", x"e4a587638e9b1e25");
            when 25970087 => data <= (x"0cd4d9c3aa830177", x"56180d7e12896f6b", x"fa8e05844b3c672e", x"7bcc46bf9a298d2f", x"0d47b0502072d6da", x"e340546c48381707", x"a33e100b66c93271", x"5a4a41d7c9aa4243");
            when 9906458 => data <= (x"88271276d6ee110e", x"31938f03daf8ab67", x"9d4648737ff7c6e0", x"acf0d58bc0d3cd79", x"033a455f479c02ee", x"042406ec163829be", x"08025b43488522f8", x"a0d8e30a3ab58efd");
            when 8612407 => data <= (x"26004a54788b2e6c", x"da3584832237725e", x"ac4df1380f626a29", x"21732ceaa578c087", x"c79f6f831bbb2711", x"5486082bdce33844", x"4ae70fef57efb964", x"fe8b9b0b5ad3fe12");
            when 1237107 => data <= (x"f142a464a7f9a7a7", x"7c080dc3b74636ef", x"81032a228f702610", x"8342db2e36cfb5f4", x"f43f92b10048127b", x"5dc60590e6de8096", x"245ede042d8ca809", x"80a9494a7d63b075");
            when 5671622 => data <= (x"074630e23ee8a526", x"64f97911655b997a", x"73e67dc67562e58e", x"818370a22e221c48", x"6629ded85291fd9d", x"ca8e619c9a90d839", x"93fd498f73501898", x"b17708d5a727346d");
            when 16261876 => data <= (x"dbc0fc0cd6bafad7", x"d29a3b363771ab83", x"1bee6f02164d9cd3", x"d91d445595212724", x"90df182294649e4b", x"40423b3a6a90e45e", x"8701ba2418f3274e", x"ff6776e8eb4dc923");
            when 1326275 => data <= (x"be24abf1d1909038", x"275440e92545d406", x"b663ccd7bece893b", x"53a0dd9a51f93bf8", x"ffd48c11ec662207", x"8cb91abe7243adb0", x"e69afdfdf226724a", x"43c2d62f63ce8f0a");
            when 19308402 => data <= (x"067966d1ebe43277", x"cfcf7ff61980c432", x"2634588f18f8858b", x"b89fff5feaf173e5", x"8960981471ad6601", x"6d3d2207649ef894", x"b9736bfe4e2953b3", x"61dbe2bca59bdc7e");
            when 8597791 => data <= (x"f4f556c5b0abefef", x"cdf6ae3616168271", x"d759e465fb88553d", x"5761e7699e63cd49", x"6ac0c3c424d6b65d", x"f905a2942f56e40f", x"d264807f5d920f4d", x"cb8d5699b12400b8");
            when 5328848 => data <= (x"261f2dd4b2bf349f", x"bed3ba46e1c52603", x"23fa4340afebbe91", x"8009436bc297b186", x"190a89875cf85303", x"173821602e352492", x"7d9419ce3c0491f7", x"8c89d6b1cfe7df23");
            when 23282087 => data <= (x"469a5ef1d3d9ad9d", x"4998e7505985980d", x"ffaa36a873389aea", x"5b0c50b5afc2e757", x"7400e916341c8a04", x"dd4904c72fc85d61", x"c8249294b159dfad", x"7639452de9ffa6af");
            when 3267329 => data <= (x"d4103897a496298d", x"b399810b2bd5dc34", x"a547e544f1ed053f", x"d078c62abca5e243", x"8fa3807581dc8aed", x"c930ec15f1db0057", x"977392ab95e92c84", x"7d6712be00908956");
            when 18325358 => data <= (x"f2efcae59b7131bc", x"315a49a3cb4b178a", x"e67e04a386fa7c10", x"85d550b44eae572f", x"21f0a1844bc7bbc5", x"22017f314209acfa", x"a1649eb7277e2f74", x"4d7a5e5759313ad2");
            when 8760141 => data <= (x"5bb3cccced31c031", x"17d2cac0c2cd984c", x"a2c70c0d795b9c0c", x"c8dc3f269522636c", x"883402e7532f7e7a", x"1551d9011b0e92d3", x"a044e7e2e56f5888", x"827b1742bc25ad8c");
            when 10957700 => data <= (x"2b0ad57e84e279f4", x"3833f8168cf3abc0", x"09e0c91c08e8962d", x"0dd8007c8ee56b33", x"00446a8cac2d0716", x"34ad004d22a48402", x"7d71b56012845993", x"c02dae1dca02bdb7");
            when 9162962 => data <= (x"e5d515d6e3effbaa", x"117e086802a44658", x"44f051daeffa0447", x"7c7afb062775a23d", x"f3e16727e581c640", x"2722c3306653c902", x"35c25bd5d7c08ff6", x"d4c0385f936754b2");
            when 26885318 => data <= (x"f2a442fd95d4cd9d", x"946c4c62a027c20f", x"8f03111955a19a43", x"e85796b22b41a0f3", x"35b4232d6e78f0a3", x"3f2cdbb7e4fbfd66", x"8899eea40ee7ebef", x"ab270e3130031afe");
            when 26385953 => data <= (x"27dbb8f9995a3e4c", x"ad451dc6a410e866", x"ccb8fc8a4eadf4b5", x"94e4128dbe3e901c", x"6d34bf0415b3ee42", x"25891efd45c11dae", x"3b36602309e38dfc", x"39134988757f53cd");
            when 6364266 => data <= (x"c1b35566450a5745", x"9fcdda8aa4bfab65", x"e805f7d0c9e0b001", x"3f9aaaefd04c48c9", x"5147aead4f11bc32", x"48513aa28232e83d", x"818c3327bdb0de62", x"a79c97568823091d");
            when 31474125 => data <= (x"ac51b23f3d0aecdc", x"6a512cce5351e8f0", x"9bfbe1cdab3ef935", x"c6fa2283cfd280d7", x"50ff21f0e043f417", x"b35e6f3a3fa840f6", x"1a8eb33084a37947", x"ae2d357c1f098ede");
            when 26233924 => data <= (x"9ec8cf0e429300de", x"b71250b33d5112a4", x"0dfb97aaf14d8013", x"68de6db346b71f6e", x"960ec59657030892", x"092f6bbecf7f948f", x"53a5e90512f82aaf", x"ee606534ae5c6d56");
            when 20502242 => data <= (x"9f929042e6763ff3", x"06f413565c11e787", x"103e1260164fe65e", x"bb259e96a465b26d", x"0beeb96a2d64aa66", x"dc22335c3ae92ef7", x"ef4222368490b344", x"4eacf6948b422c7c");
            when 9142229 => data <= (x"a4a6eedf1a68f2f8", x"22929f13f4ad8d8d", x"f5f016569982d7b1", x"1475dd3fa26eeb1d", x"f26ab23d0cffb76d", x"449ca796e8df3377", x"f9bf5e9aab51c555", x"9bec5b83c79dc699");
            when 25912831 => data <= (x"eeb229630f5affbf", x"aeba263a6f5c6779", x"87b3b48565bfcfa5", x"19ffe5b03853be21", x"4353955a45ef8d5d", x"561ad37ef3a234db", x"8428205627d76d1b", x"bc73d3c032232fe7");
            when 14797557 => data <= (x"aaca577964ff2c5a", x"ea73197d6011261b", x"15ed1052d648c8c6", x"02aa4932bba2eaff", x"bf567bbd914f5f31", x"9d1ca1dbbe487512", x"d89886fe2bc91317", x"b7ec76b9db10c163");
            when 22135392 => data <= (x"61ffc1350eddff78", x"c1018415e7a2f0a5", x"c2c6da14fdae7857", x"7d831b814ac6fe80", x"478e2d4c67778665", x"69bd6219b4b703d5", x"c4d0195e024d584a", x"d28e48fcf8c83da4");
            when 15408851 => data <= (x"e1ea6ddcceca2750", x"6da53a161f5de09c", x"d434abe62c9d5041", x"5b379ff5410d787e", x"ed1330dd3aa63600", x"8cad7ff99320300e", x"f19da0f240bb3564", x"839c51ad4b6766f0");
            when 30506977 => data <= (x"e89a78db1ce93355", x"733f1c69d7fba463", x"9660b2be615e6063", x"bf1e016a99e69726", x"e46b5e1585c67c90", x"ce27a1e2c450c812", x"f8270098776772ea", x"8d6b23a83e596210");
            when 2135051 => data <= (x"7bb4ad3d477880fe", x"e6a76392806f07b0", x"1c5abb1d22e6ccd0", x"e6692630a861fa3d", x"143d5130eacffa77", x"e5a98aff4c46b2e7", x"82b31c20df1b3878", x"128dafbaf6305031");
            when 20406402 => data <= (x"df6891fa27dab1f6", x"94f03905e30cdfb0", x"f44c9c0f0730252d", x"def11baedcd91938", x"b58abc9681a2f76b", x"43e28e4ea6aeaf09", x"42866d50938aee76", x"17e76f247855b58e");
            when 19155899 => data <= (x"902104504c0573da", x"84768528f59d2eb3", x"71c9a1ebc409f259", x"25a74bb8f636ed04", x"f929390573bd5fa3", x"f3afa376e7d8f23a", x"d55839a7b4089314", x"6c8a05bf0fed6603");
            when 13870660 => data <= (x"50a3f13484ab0496", x"5f52b255fd08eeff", x"5d4680231d8497f7", x"b735cc60aff0dc66", x"3be8b0e46d8bca82", x"c519a838708af30a", x"a8a2dce47831cb75", x"8197cd72879a206a");
            when 13807750 => data <= (x"41c32fbf8cbd74c5", x"3dafa9951f33cdeb", x"47e0a34f3c7d525b", x"0381ab4a212aba23", x"b0e2df8b0f7e558e", x"bd5d37bb3dff084d", x"6bb05097ed420a0b", x"bd3e7fefe1e40453");
            when 21663722 => data <= (x"55b0f087f60aad33", x"ada1b9670bbcdde7", x"2f31d75e017071fa", x"4d154390a5898278", x"16f5a802aed71249", x"c3f19ffef178e621", x"bfd64b89176c1d18", x"c3e1ae139c941821");
            when 16775137 => data <= (x"770779638bac3580", x"639ce96da800dd45", x"861094e1ce7815b0", x"1ed2f3cb5f658b35", x"06a50a5beb226975", x"da418778c94aec77", x"921fb569054278e6", x"57b03d0a130cdfed");
            when 30193320 => data <= (x"59df623851721b21", x"35ba42614b130d1b", x"6f0ced336c87a602", x"11982c84b7a77742", x"67ab9628c4481506", x"266cc0981954773b", x"be1bc2d70bd5c8ec", x"056cacd94277ef3c");
            when 6547559 => data <= (x"42d803b5755514dc", x"756f37dc56ee2327", x"adfa5b58b8cafe6a", x"2cd5a5ea02424101", x"2b2b7c18e1b9d51a", x"b4eebc5af30ecfbd", x"027488850e368e2e", x"1e0879ae2b181713");
            when 3075564 => data <= (x"e909fa23ba2c3162", x"1e5790a7e432f7a6", x"af187a0045f87c98", x"cba221ce781d1974", x"d0afd8e0a237067c", x"43dd4da557cb1641", x"0ed9781cdc4be571", x"de7f0ce5d26cde78");
            when 30896776 => data <= (x"dee4599e507b9e6b", x"a5848b0ec020ecfa", x"32e2abd39baaf7f2", x"8ffd980badc50da7", x"16b25183504217d1", x"12a9dc32c9fd30f4", x"cbee187e073b4821", x"5b8850ac0ad2b1b4");
            when 8797270 => data <= (x"6617aca1af650b7d", x"20c9efbd2b2422bf", x"b0aee7aa7961d67d", x"3305a8d52972f2e2", x"8056b5e77c4d7e43", x"82018a81c20046b8", x"daca36c8a8f7bb42", x"b723adeef4c81299");
            when 22737122 => data <= (x"6e52af4f971ff258", x"bbcbabe5d531d90c", x"d5d25ef4a912a83f", x"e6255842b05de005", x"af7329867afba7b1", x"136bd7bfd437adfe", x"8d06cdcc34bb8e35", x"ca5f8a50c524a5a6");
            when 24357401 => data <= (x"8104467a69f563f4", x"4d79a94b193e3a54", x"eba8a5b73a635d55", x"0620e71048794904", x"b546d6464fe7dc07", x"9cb86de514308708", x"f637cdfbecfa34e3", x"c45e57cec534d712");
            when 9586248 => data <= (x"503b53644d9844b5", x"9d8c34b689ff7d1e", x"fdb6635060d42aee", x"6334055fb1eecdbf", x"05c2247b4f927565", x"ee4c2486e54cd4d4", x"90d0c3f7af85ae25", x"2737bb665dc0cd79");
            when 25473529 => data <= (x"2a1083d261c507e4", x"ab541f8f21bdc2a3", x"bb9583001e512f87", x"d34173251442b52e", x"f9c11101d59fe5c2", x"7da020381b3a5d8c", x"375c86465fe876fa", x"716611b30703b95b");
            when 16834371 => data <= (x"b248c5e7be626401", x"4528b6bee499870c", x"994b700f8e86e4f4", x"4b3b322dd1df76f0", x"4cbe4f9fbcbf5e6e", x"cfccc4d2baffbca0", x"44d8590bff7a5602", x"4cd2e7c257f21928");
            when 6528157 => data <= (x"ecbe6ebdb8c75ec3", x"fe4bd611ec34c3bc", x"6918f3abd46d64c6", x"552b58b6b00d9dfb", x"9ac901002270580d", x"3ed730c52f27d16d", x"b1c8eef0aa07c310", x"13ebccf96b636f8c");
            when 21465217 => data <= (x"975d5197e7a8c37f", x"c5bb6131359c3608", x"3a421efff319321a", x"5933c3ae4b9f383c", x"aaf3e36d32c59064", x"f1f55515ca3861e1", x"d8730a117b166adc", x"efc9a0cd663862e5");
            when 13571069 => data <= (x"71a5ae4fffff9a3c", x"c35efd4c417e9047", x"e616d63f359c0bc5", x"940026d482aecb4d", x"aff5a3ef42ee35dd", x"a8a61259ad57f5af", x"6c3fdd5317e67902", x"c336353cc9f7d144");
            when 29652591 => data <= (x"d4b3fa05460851cc", x"d77d8e6800c1342e", x"3dabfb2da5fc1f42", x"76a8bd96d9d9c71e", x"8fc873a755ab83ea", x"cb4c1eb3affcf664", x"2faec4ae1921cec0", x"c444eb1db498999d");
            when 11736231 => data <= (x"11eba75d097c9789", x"6574ecf279394acb", x"92c82c3213b32371", x"e2e41523a9be99d0", x"d48c423a167a4dc2", x"2cdb4a01bd7d1bbd", x"bc93f228881e8eb9", x"2c7920debf5d1a4e");
            when 17801203 => data <= (x"431727c9b685f459", x"47a1790bb6f47d6e", x"78f94714eb20842c", x"c7edfc732e541ad7", x"7ac70bc0f2061216", x"cd1d57e73361cf09", x"b3f92fb8b050b382", x"ac75b644032678ea");
            when 21535885 => data <= (x"fd0104c7490f676f", x"b663bc868f4c60a9", x"17948314a0bee4b3", x"3ba456f02dc9d416", x"57436a8141c0abad", x"bdd189f1d6bf3378", x"83bc8394b2fe0605", x"31d4f1478af8c1b0");
            when 19729798 => data <= (x"5e528661869ffeb7", x"1b4c11f3baad64fb", x"7f0fc87fc5d49081", x"708cda9c405b2e04", x"beba91d8a9fb8a21", x"e671fb66b3a34b34", x"899e330a7222f07b", x"2de7e546372045d2");
            when 29650046 => data <= (x"0e68c6c8093f949e", x"8dcbcdab15963804", x"e898e19074861a3f", x"b37cb57a6a76ea60", x"abd432d924d86559", x"353053995a64d087", x"1543d3937716eba0", x"59042d9a6a218fa5");
            when 23673782 => data <= (x"fa14dda6a3efce28", x"b077e7cca73a6d86", x"cd697d9aa13db20b", x"c2cd6212a2fee12a", x"b620e2ca61174b88", x"83c37bd9ef010da6", x"7c508f8a077fc742", x"bfac4ef13467f281");
            when 22949420 => data <= (x"8e051c170a4a5db7", x"e3f941066679fe84", x"116346017420b7f4", x"aaa4e7e8cfd66758", x"6fa80690f9505211", x"5b6dfa8e4ec0724d", x"dd3dd0e817ce7ecc", x"8c7b43008d4c27eb");
            when 19864022 => data <= (x"ad084b67ee8bf2be", x"b3a7f1f384ad5e8c", x"a6745919229f3d5a", x"35d6cdd41a348a41", x"57b575c75e9aad73", x"54a7ffb2721373a5", x"b5deac84f031558b", x"669a907d44704c06");
            when 8887552 => data <= (x"92a66c72ef924d3e", x"a71290d87a9047ab", x"7ff6229a7b735c34", x"1b9875aea2943953", x"c0c35cf8639acbfc", x"07df442608ae22d8", x"3beecfe73e189020", x"e9bd53a56e69f200");
            when 1812261 => data <= (x"3a5fd0da53d39881", x"c54b3b52c00d49a9", x"154e975278b2befc", x"870fcc680af45100", x"10b341e2e0b5ff4d", x"28cdbd1781e934e9", x"34a47619bdc9c05c", x"9e303c0f60c4427e");
            when 16980633 => data <= (x"85f9fe71f0b204fb", x"f08ee55bc2ebfb45", x"0ca268554b640da9", x"6f6f0cba34916bd0", x"78ef7d3d3c882f87", x"b36e4d080c461d46", x"213a6035ea77029e", x"0d6402b9676f1164");
            when 27719491 => data <= (x"d54f001a9594ce4a", x"1e4b4c0ea8cd8ce2", x"243cd1a2bb2172f8", x"105569a4469a657f", x"1906b59f2b8e7e6b", x"4dd79c23b38b8a09", x"17c009892eaa3fbb", x"6208bdac802f3f3d");
            when 823043 => data <= (x"01d265934793c69f", x"4b1b45e2f2a449b2", x"439a9faee9daf3ce", x"98270eb98f4855e4", x"60d47d3149ee48a7", x"c4c21437fbde794a", x"12b664e5237048d9", x"f21a97f8831397a4");
            when 7394159 => data <= (x"570251f539f60e8b", x"094fd128593dfc8a", x"9a8b27cfacb4dfa4", x"b86d866057bd7e06", x"40cdae067b2f56d8", x"a176924c0ca9a759", x"fe6dc728505ec48c", x"bbc730a5dfc74ebc");
            when 19689977 => data <= (x"76f9c72ea6fbd5b0", x"b81d73a66649c442", x"a0401e5bc30cde3a", x"335a989cefa11f41", x"358d86b3f6a88261", x"4150abeb40581e60", x"a88dceb651db90de", x"2ed0b3add6168130");
            when 10692047 => data <= (x"91ef6ecdce390166", x"529ea63d8e177a9d", x"750475f3c52479c0", x"8ffbbb872ddc5690", x"e88cef45398b6e8a", x"ed966978425b2a0a", x"9da145d54c96fc37", x"07537582d1180693");
            when 13256067 => data <= (x"39b371ee0ab2a6cc", x"27900839502c5e0a", x"10bc214ff8fa3f85", x"b8e638d6dc5c592c", x"ce1c41e0a2a0fe55", x"a09195fa9021b167", x"8acb43a0cf803b70", x"6fd8d7a1511d756b");
            when 3739130 => data <= (x"6c9ea7a617cc7c2f", x"db9440df37ce74b0", x"57d97bd49013e760", x"3ba8cbbadbf2e740", x"33e81d5841c87679", x"acbb1dab2b7b5465", x"9ce37780c8b77efa", x"80be9bfa8aa294ac");
            when 18007184 => data <= (x"e4fd57cda7a98e0d", x"a1cd5a3754d8e455", x"3b2006e9035b25db", x"2e4a1f30eb28ec1c", x"609026fd69414eec", x"d55cc7b77bd10ae2", x"935c72801feee47c", x"5c3c724ca4d7dc72");
            when 26067418 => data <= (x"ba2c9181d3b555ae", x"7a3fd46cd65a02d4", x"820679adfa40fde4", x"eb588a0860d3a187", x"704a3f50ea5a96d1", x"0437bd1a5a115c92", x"010fc9974b8a7f96", x"ca6c68db18375dfe");
            when 24658267 => data <= (x"f731b670c0fd5a13", x"990cc3cbc82268a1", x"1155a675cea00dcd", x"9b542c968ab310d8", x"444bae12cfd7c756", x"898e3ef903a70827", x"cb462922387d6995", x"bfdb5d4dffdf3ca8");
            when 11675095 => data <= (x"92154d70ab5ab114", x"3122f3b753fb1379", x"0cb134e32ef930dc", x"3a997fc4cb363b0f", x"d050c65daf74fde4", x"d7d284f6ceb19c8d", x"83fd97aa98de3f45", x"b63e3abb5594e273");
            when 3596485 => data <= (x"3236d6972c1fa03c", x"0a4f2c1b4009ca1d", x"f91eba2f35e60f79", x"a6cb391a1f8cad1d", x"53988c08aaf50b53", x"b9567be5a084a0c5", x"ac090377dd2f1f6f", x"d0b81147e5e59bd7");
            when 27518397 => data <= (x"1f4d984cbb605462", x"c22ae5c77ea6739b", x"417f6099a103e6ea", x"8283bdd6449ab281", x"8f995606224939b3", x"6adee18ccde0d496", x"04b33f3faa1b1f59", x"74eb36373cae6f72");
            when 25727657 => data <= (x"4f51271141fbc228", x"70bca1d98db30afe", x"babfa0666464181d", x"32f983b4596657d2", x"2d1c671590cbe640", x"94912f5680856c86", x"5698f8c050d77314", x"7b8d6a7085c85dd5");
            when 2080871 => data <= (x"61364da274f2df42", x"f9b8124548521392", x"47f9c7790e74ae0e", x"3160f792d5951b50", x"cc3fda4e59c82beb", x"71c8a9a479edfc11", x"fd0a001577adefac", x"b0d472d9b5fbca44");
            when 11301034 => data <= (x"f602168f1d36f7b6", x"2e31ce010b38d3e4", x"9420d4a8cdf1f0c7", x"9f22c4a67902eb8f", x"fc048272bf979ae9", x"efaed76d6af5f38c", x"ef76c76a018682b6", x"677554736d5e83e2");
            when 32350577 => data <= (x"aa686731058bdebc", x"bb9bcf43f8848764", x"1f9e3745d2bbee75", x"b86fd03b401d848d", x"d22ebb95087e3b62", x"87078ec380054737", x"50bd4360acc09807", x"e23d0f04adfab756");
            when 31631374 => data <= (x"9f084c8b53bd9a6b", x"57e53bbec14d46ee", x"c00ce9260bac021d", x"9c40debe2e708502", x"5df9d6eb3f0490f3", x"03cac95b7dd4f86d", x"cdcac0a78d82ea73", x"e7197a54cd5b5b22");
            when 33460571 => data <= (x"899b705bc68f5086", x"811a18f3189f2adf", x"b9cc42ba7be65565", x"723ba180f9c3cca9", x"dd7c00386f5309ee", x"62638e725e4d19d6", x"5fb1718ee6fe74b4", x"540042df5e001cf3");
            when 23818986 => data <= (x"44e78e977ef99e99", x"a3896cbead5a0148", x"d908cf56eddb915b", x"3f036ba05ce5b6ae", x"c1a1152fe016a4bc", x"2910a04fd5da6a06", x"3b7e7e8e5cc64f0b", x"cfe94b6193fee62a");
            when 13852273 => data <= (x"bef3757b4fbd35a7", x"f13445875cd0b4fa", x"559d05823e6b4c22", x"8231d7bb2a0e260c", x"7d1da4f3cdf1f63a", x"fa0f26e2818dcc24", x"4a38500572d25f42", x"bc346954324b220b");
            when 15422229 => data <= (x"8feb5ecb7cb839b4", x"453d286285ff9340", x"d5c1ff3d25f11437", x"f5215b04c74c729d", x"be415c0b5c5e1177", x"539a4357077b3e47", x"e429cb4ecbc08129", x"42196ce868b9a3b4");
            when 17805087 => data <= (x"e378885e452a61db", x"43a8e28f6bc70f85", x"7049563b3c70fdaa", x"5048f29b44ed500a", x"df246e60f7371ff4", x"40ec7461403065e4", x"246b1a9e93f3f601", x"02da387a4897f87a");
            when 22767141 => data <= (x"2a740639b602491d", x"b8da1ac80802a51c", x"ab2cef6f7ebca7d6", x"ee805d64fb908415", x"8aa8e5664d31af71", x"30f6469fe7a3eb3e", x"1ed149f30363776e", x"e5780aacb4515163");
            when 32082877 => data <= (x"3d7e6bc411627fb1", x"8e3448ccdbb8da90", x"3f95e952fd785f58", x"c475d29328a62e14", x"6f131d67b22e4c91", x"9aec062bd79db8bc", x"aacfb83122320b35", x"bb6b304d01b0bd32");
            when 22291207 => data <= (x"919f15cdf26da15e", x"40cd2fd68fef9b31", x"a16a8721d6817fd5", x"8639701579f944f0", x"d0c15f46083e38d3", x"18ae248a70f856a3", x"1cb70cd17dce477e", x"b3b995647aad47a7");
            when 25644785 => data <= (x"d8c3d6c0d8efe28e", x"486569e4e3059447", x"0b01132c66b4bea6", x"5143fe12ce8a4cc3", x"cd7a586c870c6a63", x"ee3b7ae8d701ca59", x"36fccf41195bb918", x"f159d27a77fdab35");
            when 2671025 => data <= (x"0f35150b37d8b566", x"9fab0aa9af8e1c07", x"de625a8099857602", x"000c90bf3b3d4dcf", x"89fe7ddbb5a2866e", x"ec178a66ded1fe9c", x"d43951051014ed3a", x"3f24eb0a0ee5d058");
            when 31666849 => data <= (x"ed612eb16e5b4628", x"af860e93a953228c", x"6911758cd4e650c3", x"f1e6e1b6dd1ba9ad", x"2d301f848bf39419", x"b6b7b9dc864fed92", x"c7faf9f29936162e", x"140b372310608b03");
            when 2860640 => data <= (x"bbb5129b55ee7e91", x"0ccab1664b81ae25", x"f8f22ff6f9f08428", x"a987e5d1f7313899", x"14ceb2e7aa6ad7f4", x"da8c58fd8db3f3cb", x"b0b445052694f0cf", x"4a5d803bf1335cf8");
            when 31629110 => data <= (x"154355b53c2c7833", x"47806b4ff2c67e22", x"8a5b0a85cecaad9c", x"7d28fe73d832dcd9", x"8ff73300bb11de22", x"92494545bd180b07", x"fdbb6fc127dc7e51", x"363834e881626790");
            when 25722661 => data <= (x"081fdce7777ddd55", x"5891717b46406c92", x"badd72c9673b3420", x"4647444615a59227", x"86eda4d71cb67252", x"4ee81728f1d46009", x"9ae251adecb2c50d", x"0eeb29fd3e23bcb2");
            when 18502239 => data <= (x"af6577eb0966dfcd", x"e0fe0cfa5e403b12", x"e8deed0fa5ff0805", x"6eca33ed4f7ee727", x"f29b7d558f541b31", x"014e7d439fe0a4d8", x"e80b12ef0996ff1a", x"7b61580035da8b69");
            when 12313566 => data <= (x"ca431f166b0488fc", x"338c7ad2a80019a3", x"39dceb9bece38fd0", x"a3c17715de460746", x"6a6a17d9b7b74765", x"e031a6973611d73f", x"4a5e95753bf5ea83", x"8ad8bfdfe3a58e0a");
            when 25977948 => data <= (x"ae667a1391818a0b", x"a2befe36aab18df9", x"231b985afad8cc51", x"8f0767555b4fb4cb", x"572a361a844a9213", x"1951d141066f2b13", x"347bd9ff57d3e850", x"870f58922be1c08e");
            when 31315018 => data <= (x"d7941747c05e58ea", x"22f1917aeed412ae", x"6a87439807a1673f", x"35326929f0b602b8", x"10478b00324f45a2", x"14e189c78a0d8073", x"9c03065d5d672616", x"cec9bb3a1516b299");
            when 22108329 => data <= (x"af3479cb079c7af8", x"3f16f3fa4dc7387a", x"84ddea143c6cd9a6", x"0299eb0269eda9d3", x"ef62bb79412fa276", x"1d28f80dcada0dfb", x"e8acfb94977bbd2e", x"29692a6c8dab05e2");
            when 29100990 => data <= (x"a2cdb74d29683bbd", x"1e9dfb9abdc533dd", x"bd65c2a06d2b2056", x"3edb91782c879a21", x"a8b990a634df3069", x"faceaf83fda5f834", x"4a9cd24bbf5b7521", x"e573574696c0cf80");
            when 24125743 => data <= (x"bbca4d27bd58ee31", x"4b6382166e5ccf97", x"650358f376fa810d", x"dc73311c692bf262", x"155568b5818c42a7", x"bf35dc2cf48b8703", x"5da0b3f436bba98c", x"238305fb18dc98b0");
            when 22603205 => data <= (x"11f1b127f480d3af", x"2d201fcddbbd18d6", x"6eaff3aed8aac38e", x"bb1959505646aa6c", x"411c307fc768a556", x"240c4ff11111f955", x"86e3209fed2f073e", x"200a34faa8599c2e");
            when 10620587 => data <= (x"340962bc457d6c98", x"a9c7e2028987a3b6", x"9da07994eb1e5e5c", x"27b1870700ae31c2", x"20b8c459d8222582", x"5f7ace5540caccae", x"3a01a0fd243731f0", x"ce75d9c136a16c35");
            when 4449831 => data <= (x"cab2e986efdd54da", x"1de8053d2332ce39", x"eff98ec228cc6e9d", x"5b0687bd470dcf2d", x"ee66f9e9f14693f1", x"6e7aa1d6c84a8114", x"83ab434b4ab18ae6", x"97b156f5c5808c38");
            when 5236626 => data <= (x"333406b6aedd094a", x"51187b998b173eba", x"d75c7bf973c08d23", x"0fd1a6f070ea1568", x"4a3d977e827770ae", x"0cf68c3f26ed8f83", x"3d4a9d059ccf563b", x"aa02fda5d6db7281");
            when 7740215 => data <= (x"dc76d2ef6cab73c7", x"dc195ca2ec7aee67", x"56e903c678b75872", x"f0b32eef2e5ccfaf", x"23b5af20f2a06341", x"7c242767778bc401", x"275a855163e61eb3", x"b08364a85f6380c6");
            when 17230867 => data <= (x"bd8fd7e853cb224c", x"8b960cfbcb668865", x"ebaf47b4b2df1fd5", x"809c2035497a5c81", x"1e139730b7b67c35", x"bfa0223d63edc1bb", x"eb0e3eba90540719", x"cc25ac11b92b350b");
            when 3865120 => data <= (x"caeb3b907dfcc78c", x"bf7578d8cb95f2ca", x"395570a24e2d8f47", x"facca57bf075a0db", x"4b668a2bb207a862", x"50c37e4f084446e2", x"002091885348c159", x"0f37958c87daf8c8");
            when 14024851 => data <= (x"8e50759d0ba8b23c", x"dbfc5f2dc6b2f4f7", x"e94b5e63a25c2b8b", x"034b89ae4898fb32", x"3a737bac231abfc0", x"4d12d81befac39ee", x"806901ec85b24147", x"20440a52a55b2de4");
            when 22894336 => data <= (x"a34d21aabfad15ad", x"41c961de38499083", x"b3ebb55b27268356", x"51a0f2ecfea4921d", x"e113c330d9272acd", x"bf0f84e5b6d0e2c1", x"59ebe64fef3ad817", x"d4db207c4d6104b8");
            when 23142836 => data <= (x"fad41cdb8a2f5b69", x"71dc215ef61c139a", x"94f9ed2eb5261458", x"6fa96f0205d5c66a", x"c51914be8cd3e4a0", x"55550342a6d249e3", x"6e8d007c162d4a72", x"2a168dbea8e5a216");
            when 6025937 => data <= (x"d93ffde50106928a", x"a893ec0f88f79fe5", x"41d0a70e453c9881", x"253d5795be49d064", x"74bbd9eb756982f3", x"7ccc2417f1f0d885", x"2085c6358011eb91", x"575e20360dd10190");
            when 29480314 => data <= (x"3b3b689fef3c4f4f", x"e3197d351bbe2baf", x"cba8d99ea4887106", x"0a8ad878d4670ed8", x"cb066497141b2ab6", x"d3b744860484bf23", x"23154e84478193a7", x"5e1fedc4e671986d");
            when 16088658 => data <= (x"8189d9b4278086dd", x"282efc8ef2b55dae", x"bd3fe29af09f82cf", x"a810758faf3e10ad", x"d87f406359842ba2", x"090af7bc3200b53c", x"3d23431b2012d69d", x"b7c893b13c21e87d");
            when 14465549 => data <= (x"e1039d7d4fb35445", x"85187b55f72fe27c", x"9478754913d45190", x"74ed310d4d67bb34", x"3735d0a5ee189c66", x"d71aff32c90fc0de", x"8c223b06efd5f66d", x"d57fb09fff550b51");
            when 10516027 => data <= (x"f9b24da4388798ce", x"7bab0f73e2acd7e0", x"b9562b353140d1c4", x"2f508eb31692f6c9", x"01c4e03724f5f2b7", x"01abc944b5662d08", x"5d9a504c8aa124f5", x"448d660021a71823");
            when 23289864 => data <= (x"d82ecd881e49b38e", x"598bc867717d3e4c", x"a7cea5f601c6ee99", x"dd023631cbd94ff7", x"d29ea3c5977d7ae2", x"e489adac474502d6", x"fb69a16f366d131c", x"e724192a811da4f3");
            when 6614743 => data <= (x"507f70a25df371b7", x"00023054b932ecdb", x"de164978ede29470", x"d1ee0c4829985c34", x"08460d7634c13275", x"bf6d39b99796ad76", x"91481612c3524e5a", x"67c37c27039850a0");
            when 14115709 => data <= (x"f3ad2f8fa61919dc", x"2a8127eb943f59fd", x"98700e1a3de0ba2a", x"b3fd40f98ca64d5b", x"09ef2e0a0d68728e", x"7d8f471f5b0d74b9", x"a2e9bb24a56dcef0", x"1c2ec3b72bfaae8d");
            when 31575579 => data <= (x"273e71f44ac43ea5", x"b904daf6dbf3c012", x"4df5cd114afa54d8", x"aad18a2459ff8723", x"6274a881a81e1e65", x"13e17b1d02f661fc", x"48a919ae1d43b838", x"2e8556d432778525");
            when 6343820 => data <= (x"099f216179640f66", x"7325d3fc2b87f1d6", x"4884b1e30476dedc", x"c7cecd7b6931f08d", x"d67ad7bb1fd6b617", x"a2c392fcb0f50190", x"2e5ccd0e431dffa4", x"50e0741b92858aa5");
            when 25396802 => data <= (x"ff0b10eb805c53d7", x"eb649ba0c3798209", x"dad17780f6b00c96", x"bcd06051f74649c5", x"92705c0c1a31222c", x"9ab088e57985c6cb", x"ef12a44c7162981a", x"8cc1ae4901726f6d");
            when 6768252 => data <= (x"55e719b77625bfa9", x"1bc2031d20c3ab2f", x"ed487b6c92d590ea", x"14f08b7d365030de", x"8564d33b73390aef", x"20dd8e3249cf141f", x"24adffb9d9be3c0a", x"b48c6efd71e6c6d6");
            when 6009969 => data <= (x"969521af0833d2b2", x"2a2cfab3cb8e0e2d", x"783f08c87db4b791", x"3aa705419eb29222", x"156e64e51121ea73", x"41a3e1c6ce59b0ca", x"7a25c95e235b308e", x"595b4d19328809a4");
            when 1430990 => data <= (x"0b4d279dc3207a67", x"2de388bc408e0cc3", x"c8a99dd04ad6192b", x"4a803ee04ce29704", x"d58625c4bcd2f48d", x"5510e845ae2dd766", x"68e078f8ae78aa58", x"43d50b24862c2138");
            when 8454923 => data <= (x"d4ef31bbe103db94", x"11972ab2a81cb6ed", x"a63a2d707145bb43", x"fb4ae33cdb87ca0a", x"cd72edade1a04656", x"75a88ee7e9a40425", x"4261c0c82de6b672", x"288f2fda6b5f8a7d");
            when 14958716 => data <= (x"5f798551749eeb89", x"e43a64d2befb1fc1", x"9fb796d2eea5f841", x"178bfb45bb2b6ca6", x"9628919f623c90d4", x"69e37a75b0569b32", x"bf61b4bca4757a0e", x"4b092cac342bcd35");
            when 4147145 => data <= (x"dc5f46deb21012b9", x"9ddb579a16ff9562", x"afc931d757cc8266", x"16792c01b179959c", x"0e20b558b04e08c3", x"6103f57662968774", x"80c0588d8ca3a144", x"d3a47dd5bca96927");
            when 23177752 => data <= (x"4f06fd0d1262bfdb", x"8fa4e60a21e59477", x"519cfe1fa5c9f2d5", x"13ba80c650ebc31a", x"04beb89e9b4e2eca", x"bf9b391858ed08b6", x"9c7a533382a725e2", x"0a71af46f055d025");
            when 2694001 => data <= (x"64ededb2c972b6e3", x"ccf04ccf66c64363", x"58471d1f47bbd644", x"cb29021047cbd017", x"a435302f9f0c713f", x"b98e06a24df84726", x"9c92412d2522d554", x"1dc97a21f1122ba6");
            when 33008801 => data <= (x"cd4172591a6f7063", x"9e05b6fab533659e", x"66c9b2f9df7fc43a", x"079a666d0c0825e9", x"c889cbf3d8e7a074", x"70ebef8e888ae151", x"8385e9f914b51562", x"65382fd8c1c8b228");
            when 13813017 => data <= (x"2565587049cb8d1e", x"424ac03d7207141a", x"6e1b65816a5ac260", x"b28bf06adada285e", x"c58ecd8de525d7d6", x"6d47948b11dc7129", x"2d88ac5021235d05", x"c4bdc475294dea5d");
            when 4808535 => data <= (x"e78bcb3d04969b92", x"8fddb26950be9314", x"906d434d5d326bb5", x"a55026281f9a96ba", x"55562ae6f073710b", x"192c30614774faf7", x"6257b3a5da7645a1", x"427e88326b108ee1");
            when 21871401 => data <= (x"b21de19e31d5d81c", x"82fe3f938c3ecc27", x"275df62ffcbd5b71", x"3e8c695a6548103d", x"c98725b1069edea1", x"a22acb398c886aa6", x"86f4e65a60ff9410", x"4c62972b15694ca1");
            when 6701336 => data <= (x"159098090a77f568", x"54da1db8c23ca08d", x"bf94b19a7819fed1", x"9db7494b1c2614d9", x"35bb50cbc0a298fc", x"ef1162cecac6e505", x"8ace69400e4cc699", x"584d352182b54c2a");
            when 21534856 => data <= (x"44ff14f669302330", x"1462fa92ebba06d7", x"778cc4aabccd3205", x"9115d8890a46abda", x"dcd0362ea1201fcd", x"34512cd1db3e8afe", x"3cb6cca4790e0a99", x"02dc3a16c9205cd6");
            when 6047868 => data <= (x"740fb257a79cb90c", x"12df2831441e81af", x"edc3c8e78d37895f", x"3750ac66209a169b", x"12920c62cde3e4ef", x"c9c628d94b695a33", x"dfa3d1e18bc6a886", x"56b8ecd0973bd44b");
            when 21910766 => data <= (x"dd2d4abc5f782df8", x"526558d60c703f0e", x"72d95abd8c8bb59b", x"4b2e264a4fe23b4b", x"cd3fde0d4af2c032", x"549a63b0511bedce", x"ee923a0f06bc2ac9", x"967797e62df59b4c");
            when 13518800 => data <= (x"52cdf25217f69465", x"1a11829ca7abd251", x"eb9d4bd18c7cab4a", x"bea99b588e429d69", x"36baf4ae5075bec5", x"d8c0ba03a862218a", x"6c37deb9ebe38fb7", x"3fdccb9b6835541b");
            when 4521030 => data <= (x"cb98583783d46a87", x"453943c74654fc7e", x"6fc0c452d7878d2d", x"7bc4310a6aa53742", x"c2a476c5c7b83a8d", x"c5621aa3d59d94a0", x"c3c1fb107e47384c", x"92cebcb3b44ac822");
            when 31783135 => data <= (x"50566a2bdee63f06", x"4a8b627853bfd143", x"77c4bc75a7f86ed0", x"6083b7e9e099ab29", x"915938e5e53f2dea", x"95cf0dd7da941674", x"471125e4be86c663", x"20d6f39f83a7df63");
            when 32409966 => data <= (x"21314904edd12e3a", x"347482c33e44d2d3", x"bbf7b245588557d3", x"79e3fb9b1fdaae31", x"7a30d3164f1171db", x"04532513f0cbe9b3", x"711081e5e847e6b0", x"6e2cde42aa7de43c");
            when 18542569 => data <= (x"b572f59fdea58ac0", x"f06304299b13984f", x"86c5d8928e3c83e1", x"79582e86e88f0d94", x"f844aa798c6271ff", x"5693c59c4bddda97", x"6e604423efc3eff5", x"fdfb2c94f3d341b7");
            when 4317808 => data <= (x"8b1a6fdf30ae8943", x"9ff3c6a9a62745ba", x"111559e61e686e10", x"761162523f74995c", x"028d35c679a78d07", x"7aeabc70abfc6f06", x"0897eb957903cdf7", x"fc664392b8fd5440");
            when 6281804 => data <= (x"d3d01ef4b0b6195d", x"30af6f5af81b7d45", x"8cc673bf6e1da159", x"ec90f4d8e2905829", x"71ff4fb7eaad8789", x"c9702c1572b1d7fa", x"d03a07b20da3f525", x"b0a2511b1ddb38ee");
            when 30106644 => data <= (x"dec28a5af2b63986", x"f28431ae83a028bf", x"b16dc7ea8e0b709d", x"12c48293cdb4c797", x"2b0760923f7bfb9a", x"10100a456ac593d2", x"e90eca05fa7c0814", x"e1126a09d12ea04f");
            when 25900901 => data <= (x"917d023003a5e73c", x"2c0ccf6684fec749", x"f754c1873290f0b5", x"51b2478b54b01c8d", x"1267c1954fb5e969", x"286f5a21f89166df", x"7aa72d56058ee91b", x"a252716f96afadb0");
            when 18916454 => data <= (x"14ac2f253751d47a", x"c93f830592bee808", x"12240b10f315c4ad", x"af3c41f22961c28f", x"3b81016df4f90abf", x"57d07f83bb10f433", x"4e16ddb09d13bab3", x"2811656c60fa50ce");
            when 5129434 => data <= (x"12de0dee778f9fb0", x"8f5c72571ed639da", x"aa2d528d6c50b153", x"7c8ed9f5e0a9489b", x"45230f77e4a2fb74", x"0fecff5fc6738643", x"0827cecc80a98fd2", x"a07cdec9000af296");
            when 23532000 => data <= (x"57125631cf72da0b", x"ababd5f1d95a591e", x"ed6a52d4e883b6b2", x"ff61ebd771b9b1a6", x"51daf95c2688c053", x"9afe5bafa2408559", x"a70588f1cf38bced", x"a9f4493518c22caa");
            when 13509616 => data <= (x"3d55e0690f14eca9", x"f6b9888bf2a4b40a", x"ab192e0b34601c66", x"74121bd853dbe137", x"1ac9687e760a3826", x"1ea33059316501ef", x"81768ae5e664829e", x"b2389912d35f6e7e");
            when 19730351 => data <= (x"0d54ec86cf37ac12", x"fcc4d5dcfe25e02d", x"3c629fcc4946c67b", x"2a45d9aa77388e12", x"35bdc72d1368a964", x"a0504de7f3e34ec6", x"18505ea5ac8c4407", x"4bfa54d60515ea29");
            when 7663862 => data <= (x"cbc961388ca8dcc2", x"2f3ad222da359045", x"78a52a9493e90f52", x"d2d0e06fe8ab8268", x"d1ead2cb57ac4229", x"47110cf660014c96", x"a727def2769d4121", x"ced4311e58bcb217");
            when 1964539 => data <= (x"f5077660bc083272", x"7d18cab66dbbf4a7", x"54ade431721b4d76", x"86b6f4e1a0e798f2", x"f1437b315351501b", x"0517848df8183557", x"c2bc56da6c2d2daa", x"5f1770db393621c4");
            when 19065142 => data <= (x"2116fe12e6ebfc55", x"bec4f342fd6f9281", x"1b2720fa14f9128b", x"5100b04755ec324c", x"f23ed9113e452f60", x"e576a613448d895f", x"54b2d9098d3fddd4", x"dbc8c5805dc4e993");
            when 19962469 => data <= (x"2994595fff8ded7b", x"7e65414d9dbbcbdc", x"7ad6a7691c35fcd2", x"6742ef44b1be5d65", x"f9ce11364da51a8d", x"41ca259b83550cb3", x"09bfc6fd8fca2614", x"8e2107ab7e291252");
            when 18562352 => data <= (x"aef55727c54b06cc", x"daf7988dc81af589", x"646f957f0d33c66a", x"2401fb53f6c55330", x"e1d99cd7dfca327e", x"699f3b8c0b964d59", x"31c727332139d358", x"5696630e34b988eb");
            when 28871776 => data <= (x"9fccc0ba75d5a603", x"12fe9f2a68b518aa", x"ff627f2cc52183b0", x"44e73d4bcb7d41f3", x"857fd92ad6967924", x"2ca110e7625a151d", x"d192e9565be5bc66", x"31cd6decc9b4dfa5");
            when 14476568 => data <= (x"aaa19bc40a013314", x"e84bff47db93114e", x"caf8e7b566739353", x"29e9285cd375e70a", x"3fa0fc8153a08a1c", x"b102920d3108ba93", x"3518eb7106a68499", x"daaafdf567ef6855");
            when 23680274 => data <= (x"0b2ee2330e0a0fbf", x"edcfdcd77175128f", x"d61c1d9cf19fbe05", x"0b3879361c33caee", x"62365b9662a8896b", x"d1c66bec0755671a", x"e1a072470efd1300", x"7797eb8f4c50f43f");
            when 23514172 => data <= (x"9cc637390fcee7c9", x"a70a126836c20b79", x"947d15bf24ecd41f", x"2ca866bf9dc9e177", x"77f53295e8a2a55e", x"b7a28c68f528b25f", x"52bdfcaf5a0057b4", x"c83d7d89c6e7947a");
            when 2062810 => data <= (x"a8e1fb3e6dccceb5", x"740218d201a6b2f9", x"ea02158a9f10960a", x"9b4abbd4a70c7413", x"360f9c671fbf806c", x"84b65a62bb33011a", x"932bdc475b4b926a", x"92b4a2658e6a5729");
            when 21859952 => data <= (x"fad4c5aa46b7e50f", x"76a56c23da6c84db", x"08ee1430d100b6b1", x"886d1ff0edca4c9f", x"56f6f2c68888e4a9", x"922befee4b9b3098", x"aa1458e1adec6031", x"5d143a3f29ac94f4");
            when 19977072 => data <= (x"88a2d2288dd8be4c", x"4481a1b70047576f", x"1ff9a8f985d6a032", x"187c411d9458834c", x"79b3e0eca68f6b06", x"05e4fb84802e860a", x"577b42c67e5966b3", x"50940565dd843e66");
            when 5327258 => data <= (x"3e36ba583d3c918d", x"8895e3350ab46079", x"14e62513ee9152c1", x"5264368242b2fb76", x"74e97edf46bdb473", x"323dc9b1becdc2b4", x"82a7592d68b649a3", x"b06ba434a32936c9");
            when 10248416 => data <= (x"a34d525ad466863b", x"2272baba907526c6", x"21fe0e9f07847b35", x"83acb20b36470734", x"2fc26c3485865d16", x"ec2c089abd01c8da", x"0929d45071a683b4", x"b35ba2e55e29e9f1");
            when 7819028 => data <= (x"e7f8737643087781", x"1f87a92a6e95253f", x"52847aaea24635bf", x"217df6164515d836", x"e14837913b61023d", x"b5acbf0a4aac14e5", x"8108a16e85f2dbaf", x"d3619c2275af8ae7");
            when 5054198 => data <= (x"6ec175ef67a70cf2", x"e821621e8c6c9618", x"d17b6ae416369bb7", x"2c9c3607efcac9bc", x"2ad2eed55c215cf8", x"c80de6a616bc64fa", x"36d4cea770e2cf0f", x"a76b1b083b9c2917");
            when 20303871 => data <= (x"5c07e4fda1ddb9a8", x"9de84de4bf7c5e40", x"24ca116ec23ba0c6", x"53897c88dd0bb21b", x"213cb60b662c264c", x"a738d6b58e04d49b", x"215c5fe079cfe676", x"4603defe9d0d0f08");
            when 5124195 => data <= (x"5ae9808db2a823d9", x"ca2039e327250b15", x"b01badc0e525c45c", x"ff1ea009309a1787", x"7da799fcb0c0aa37", x"fdd71cc0cd12eab6", x"da12b4db8c24ff8a", x"2f066ae24ae0f9ef");
            when 11548014 => data <= (x"03c654e86b3030af", x"88f8474d34430066", x"716849749678fa6e", x"a827f35a5cd46301", x"4daa6757df3a32f0", x"bfd6781da42e5bd2", x"8072ea6ea36eb803", x"25ca1c3bb6a699d9");
            when 7952731 => data <= (x"6f847a6baef68f6e", x"75c3d8376ec13a38", x"5c1cfddffc740eb6", x"447c0ac529b49f70", x"c5ef7b4f92e60963", x"0630b56f92bc4a6a", x"eb9fac24513a8a59", x"d51a68bf70c9714b");
            when 28482781 => data <= (x"d233ae0040096579", x"d63a8a7cdbe45c8d", x"56887865e40d80ee", x"9f72378a0fa28ddf", x"6e07bc84241fea64", x"27719399c5fcd46c", x"ebbb36897b79271e", x"8a550dbb3c8b6d86");
            when 13020731 => data <= (x"62ad3a5208dbb299", x"41067a16220ba2ea", x"400b7fccedfe3f55", x"d869e343f66aae0f", x"ef89dd0273bf7a18", x"5a0143f5c31de4b7", x"7135289f1d68b086", x"88841b987aeffad8");
            when 5963723 => data <= (x"460efca1a2f5851e", x"9f1441902f5b3a19", x"4d287a5e68703fd8", x"4dfd3f29a04f515a", x"697ac4b9b6054a75", x"89eccf36983656d2", x"fb6f81d24f67673c", x"a9948a7b7365c4af");
            when 25731279 => data <= (x"004fae69595b0ac2", x"3a87059a18bbf228", x"00e2d1f3aac7c707", x"e0f47a75f50525b5", x"44f209e435e36e40", x"dd3b71438e3959aa", x"7a34cd4d6a2f2cd1", x"b478c51597e56154");
            when 31038131 => data <= (x"563db96892aa06ed", x"0a4be50c88f70754", x"35784dcfe49e0cc6", x"995e9c09cfd21c00", x"bbbd8cbfb5c3a652", x"e803242ecaa8e4fd", x"dd89fb6a0170d582", x"1a85f82397b01a15");
            when 3039448 => data <= (x"0c8c1f4184c9a2cc", x"b81e43c723adf290", x"25b2450f0e2c9aec", x"f8763e854ea206ac", x"b83c05b8300a9272", x"2f1006357b8e2dff", x"8c93bfb38ef685b9", x"450351aa48492e63");
            when 18617458 => data <= (x"0854357801843b9d", x"a33f3fd957f7e8a9", x"bd83b5a6f0a86317", x"d1fc1f12febb062c", x"ee964bcf5eea6ffc", x"0a6d4831c4bc646d", x"eb74bf29395f06f8", x"cd332586ab933736");
            when 23629482 => data <= (x"a02acb75e4cf0636", x"a7cf4062029a0f82", x"7689013259391a66", x"7f561269e06ee4f1", x"eddcb2c65e4fa350", x"f032aa7978f38fe9", x"5f08d5464e1836a7", x"acc130c35a388e4d");
            when 27176266 => data <= (x"dab5824869b9a3f6", x"ec083196e9658a39", x"5e28c7318e843db3", x"9d6bf34778b309b7", x"2b35b659eff812e4", x"501a5636fac16b9f", x"37fa33921cdfe5e7", x"b30fccba214e28d7");
            when 27297033 => data <= (x"5e106cb73f3460c3", x"a5d7225694cebee8", x"45ae2e753a5fcd9a", x"97491aeebd1af98e", x"b77dd29f0c9031cd", x"0034ccdfbdc14093", x"05506f941a3a9e17", x"e8ab0dab0093f52c");
            when 33771738 => data <= (x"b9d83d54e029ecb5", x"d10dfd1c563a30c4", x"685b3fb0b0eacf04", x"85b0ffa584f8292b", x"3f6304912bea2091", x"56a67292abc97d48", x"af2da5fc8ca7101a", x"637554c27965ff9c");
            when 28163352 => data <= (x"e7ec7161f1871fc7", x"cb7bfaef737a659c", x"99fceaf75cf0e955", x"28d6a59897e5e396", x"3cbf36ab6ef2f533", x"9c7273cc91085da0", x"f7cabd53a6097548", x"a2d878079c84e086");
            when 4990803 => data <= (x"10f5f3b2419bac7c", x"fffa441c192c11ad", x"713b7ad7be0e151c", x"ed839256360bfb29", x"641f71251923b64b", x"e71fba23ed4913f8", x"eaaff2e988d3ccf8", x"4e56a5df5ed4b817");
            when 885252 => data <= (x"5da7d3de3ad55c90", x"59588ed2daf01529", x"37680b003acfd8e0", x"0a0f3dedd731f382", x"bc6aecc973495790", x"cd4583905f0f42b6", x"bfacb7df33aba39e", x"3ada7f519018bd92");
            when 8900548 => data <= (x"d3ce890a4ddfaaf2", x"a35ce13d14d92ac9", x"2dcd078177405454", x"0c22899f005901dd", x"d56531f2104b3152", x"2828fc2238d0cbbf", x"21fcc4f94019516b", x"45fca18ae9a1a95c");
            when 15181554 => data <= (x"f04f768a1fa5f51f", x"2a24b6cbbd695e6c", x"1984ce8de313e41d", x"9e0903486135101c", x"4f12c99fca0a3c03", x"c4bfc0bf4fe57410", x"2f941a57a4607b75", x"0b86aa40c32d5c3a");
            when 27226885 => data <= (x"535f1cc2f9339f86", x"6640edc3e6cfaee2", x"91f66e972549e3b0", x"aa08069d55054921", x"4efe3c5ebfb9a73d", x"0c886c94b0cca85c", x"37b89122fc6d76e3", x"0fdae3bcfad5ce39");
            when 29836677 => data <= (x"2e428005ec529c79", x"71d815c666c2558e", x"2aed3ceacebf86f6", x"73ae64b9b34acdd3", x"5dbf3654ce431dba", x"fcdc9634c0473845", x"81ea853fe548cf2f", x"1460f8d9ae030db8");
            when 3993546 => data <= (x"6c3397fb1e97a2cb", x"6e0fb1f7cb04cbd7", x"71f434a6fcb21a6e", x"1164d91a2fc94f40", x"9e4cdcf4932165cd", x"83078e5111b26df4", x"038659fd0a8d0241", x"e9adbe2f01a17578");
            when 15033385 => data <= (x"7e1bf7becdf851e5", x"3eb2aeaf4e91faeb", x"cdb7891327577dbc", x"141c706f1e1930db", x"24ea935b60ce9d75", x"abd1d6ac273f5bae", x"69454c03b87262fd", x"98747a12b4f9b69e");
            when 9869578 => data <= (x"4e9a05fcd2f84e83", x"2bca6ab233332d21", x"3d87fe86122f6897", x"e30ddc3bf0eca996", x"5427bfa99699a3dd", x"4c850f7565cc0df1", x"03c1512adb98ecfc", x"5fce9ddd59780c77");
            when 33238523 => data <= (x"60ec582cdf57d16c", x"c0d87d8e9c780d19", x"58086270b65ed0bb", x"6a91f0962b2f3c75", x"d41badafdd10ff1d", x"f4405d48b1c58c9f", x"25abf612fc848edb", x"315760d512fe4cd9");
            when 23565969 => data <= (x"bffbf322c96babfe", x"42ffe9dc9d219ccd", x"f3777649e4593dc9", x"8bc5766645a3d103", x"ae466162aa1d45b2", x"83bc7921982c3d5f", x"6a816d5c89d57f75", x"9ecc3e0e507a1ba5");
            when 27811495 => data <= (x"4e0ecd77034a9ba2", x"eb41f4381a9c1141", x"cd9fd78ec71c7de5", x"e2cca00009d2e20e", x"96d354a246eb2ccc", x"086cbb49c8fed97c", x"7d30356293a16eff", x"915c8019a4574844");
            when 31058339 => data <= (x"456d8917ce96c1d7", x"319708c84dd9a1f7", x"1e49b2c9aaad74d8", x"1496418d0caf8a8a", x"996abb4bd8d07dc7", x"92bcdce9300b3aca", x"07667283ea2300a6", x"9220b09adc56c708");
            when 33151437 => data <= (x"45fb4ab37dc45f52", x"631d301fd30e452e", x"018367a08eb8a2d1", x"162a5e2ca630db36", x"3a560b9c5f4df699", x"9e8ec31adf067ceb", x"9fdb4a86386a4de7", x"1122505cf5292df9");
            when 10174323 => data <= (x"9636f76095140ebd", x"558335df279b8198", x"41e80b8987fe3ac2", x"3fc830cdf371cc98", x"85af498d7da2ee5c", x"f1f764e36578a6af", x"6d430bd92e880b59", x"0ebe41a63a2433c0");
            when 18870990 => data <= (x"f581405c7586c917", x"0108fc5efdf1e62b", x"90e25a16ce47cca0", x"fa9fb7e947172432", x"fbf462bd05aaea38", x"ec879f2c5ee7197c", x"1bf63339599b9308", x"a43bcc79201b463c");
            when 16581663 => data <= (x"40312b90466eb99e", x"928789ba930f8561", x"ce54bdca13fdf633", x"aa6481e9b5d429a6", x"b2b4175433d9da73", x"b1b009754803cd3c", x"50e25fd6f6331a0c", x"7346deb3edab4deb");
            when 11085982 => data <= (x"5971a6a47d197e7b", x"3f90ffc8e199ae22", x"6da398506dba7f95", x"b0bcad47f39a65f3", x"a94143e848bd08b4", x"142c4c7eace3eb94", x"4a6beef86a9daf99", x"e19633b7cc4f09b3");
            when 10648212 => data <= (x"c7fe705f0973d3b2", x"a921e4ef2ac1da5d", x"157ae99d0d69cdb0", x"7267234463781969", x"24ba0b7cf4638d76", x"90e13d79a1100457", x"f976603cc60c625c", x"904d62d4a7996f8d");
            when 10652729 => data <= (x"f3b8f62d5153bb38", x"2e5b49dc3630474e", x"b99eaf0f74532589", x"6c335d4108a95955", x"f5de58457ebe8e09", x"b7c8c7595f10eaf5", x"5abb00a006259304", x"dff450fcff7d80c4");
            when 33005128 => data <= (x"d869a534be4e105d", x"a258d52e3d5918ce", x"ae33256bbfcbf620", x"15761f6732d233ac", x"d0f1aeb6d287e7b7", x"17ac940afd9b740a", x"61cf2ed0d7bf3bb9", x"b2316448038a31dd");
            when 25000971 => data <= (x"cdfbdad1e4de47b5", x"ce05e7522c202aee", x"7f4832ecb2cfdbc2", x"854c9abb12be0f99", x"457ffffac4460841", x"2ba656bff324e9e1", x"056513620b3550ec", x"150df7c2d9811250");
            when 12442405 => data <= (x"f8d6d2a44054d099", x"2a8c79df64927d03", x"e5b6a4771769abfd", x"81a37f498792f27f", x"b3fa6f81680efe78", x"a780258572283885", x"e7c11c0f33b39958", x"23c3c96a267c301c");
            when 6331124 => data <= (x"6fb55cce96e41c68", x"d7c1da29564af516", x"e2d1c04e90196194", x"c6e2dc0da735de60", x"6f914cfda629ee5a", x"569d4de9a53acff1", x"82ce5865ae58272b", x"32a305ebb749ea05");
            when 4552735 => data <= (x"695ba6584b1e8ce9", x"6db2d52aae0c0f1b", x"4970e9c4e013795b", x"7cd7387cbccdea81", x"d50669ef61432c47", x"5c379f31758cf44f", x"fb5c42235fe46ab2", x"35c5b38751c8f99e");
            when 17804068 => data <= (x"6fc24bfa1139fd4e", x"f3a6ff995c80dcf5", x"61776fc64aa12d36", x"b24bde792d87a0c6", x"aa414f48cee083f6", x"da2c5b2b48e9b44f", x"b3293d912aab4996", x"05ce4f54e541c99e");
            when 27320990 => data <= (x"eb1e9386eef6a786", x"59fd0e1897f2378f", x"3e201d59cb67f23d", x"0642989af3aab1db", x"df55930acff6f477", x"a8f4bb8a45c6f840", x"09c6bd25c243e11e", x"5169a9bf8e558770");
            when 6232619 => data <= (x"2178f57385f1a5c7", x"219ea2880df25c71", x"84dc9a065307b830", x"ba5bb7e9a969102d", x"e0707ef7ffb6db50", x"6abb2a42c4dc5cde", x"10a669d5c1b8a1c6", x"13f0ed16c48117e6");
            when 27243717 => data <= (x"dfacb64b6ebda65d", x"7b41c19a99bd51c4", x"d58f4e89d065979e", x"389c9839db1b66c4", x"4348517334d7729f", x"e5b5de3623c76750", x"8a7e2ae4260b9a5a", x"104801489dcea28f");
            when 21102347 => data <= (x"bfe540be06953738", x"4d62f5471152c016", x"12ac559183954fcd", x"9d3d244307dfe0bb", x"c67e0f3235d9b6f4", x"82ce07112480cfd3", x"be6d3ac4379eae36", x"ca9e7a2dabe98283");
            when 18768185 => data <= (x"d7e8f646b5c7238b", x"d109c370ec63e851", x"ec92c64cdcf284e7", x"9916b5025383e564", x"a9aec3100b2bf0ab", x"729760090942fd76", x"10b306413da69a5a", x"ccb10be746fccf5b");
            when 16366310 => data <= (x"facfc2728a745b2f", x"51dae99465f208d1", x"8f53bacac460ff33", x"dfb3d554267ff267", x"deccf6a1f52a2509", x"b23f3c6ff19492ac", x"a92ee7a187cf7d40", x"61dbacc2cc795575");
            when 33638825 => data <= (x"fb3f0e91f2704ab2", x"79e1293773a08bb7", x"0b6c1657dcc84c37", x"32662f1b82ded343", x"c82c8144436847a6", x"cc8f4ed09d42ea37", x"89a4844cc0f80b8a", x"732eea3749e9be4a");
            when 29678778 => data <= (x"4f5c3db5ad404015", x"6bd7bd1fae2b3c32", x"f0cd3145646aa50d", x"b00f55f17c787ed0", x"fd92b011dd2b667c", x"f912f0b6057a68be", x"83d6c22a23ae6853", x"65208b3f0dc45585");
            when 24711796 => data <= (x"46dd847b4a930105", x"90bd684f9b8b6a53", x"002b5a431c12a592", x"b61409c4215e0e25", x"381f0a0091ebcbc0", x"a79024e32e9df706", x"79086d37946f650f", x"e939e3d681751b8b");
            when 21513227 => data <= (x"9b50b165b8c9194f", x"1700883bb453cd0d", x"b7c48bc48759e95c", x"e1c71741dcac36a4", x"d34b078262ef82ea", x"42e988e8540b01de", x"f35897b89e4541af", x"ac908a13e889eed5");
            when 3187338 => data <= (x"db678ad1486258a8", x"18bdbe1c151c9755", x"10e8f9a86921fe78", x"8f2422fceb848b36", x"09ddceefab09dadf", x"c8ee3d21e8be7d15", x"aed8c6aa1877bfce", x"391ffa8b716aa415");
            when 22695593 => data <= (x"a2e4ecff9e2381c1", x"fc33c0e365ad286a", x"b180b52ec3aa2177", x"bc76306241f9baaa", x"1b8c1bf973a2cce2", x"c0b3cc875bc12098", x"92110166ad72b91f", x"b0333f2e455b1269");
            when 15975399 => data <= (x"6be3d7dec1578caa", x"874c5de4fdd70141", x"f4b3e91089fd6f58", x"2942ca2f07f45079", x"3324eb34102974ba", x"99f3b958473c03fa", x"91d7400657b2bf2c", x"986622d3362cf2cd");
            when 27847008 => data <= (x"9164b4d235a4b9ff", x"26ed1a1dc79c5b99", x"6023c821b316cb75", x"144a2bc9f0ca215a", x"d31884eb7f7764b1", x"591bc5c04471d208", x"f77da2ea31003c5d", x"4fc63a102a3b3dce");
            when 14025779 => data <= (x"4bce59c268e1c846", x"4a6382317b20fda2", x"0cf02fdff5734c61", x"8ab1540a6257de6b", x"7ac72249411464f0", x"ffef522c130340fb", x"66a8cc1af1f2935e", x"daa3aee6fc733402");
            when 20432364 => data <= (x"56a537b36fc062f2", x"239118944938e10d", x"d64c3c1cbb846e37", x"c714628647e57d5f", x"2cdcaeb033feda29", x"44ce514a30f94fec", x"3eb7e1f26958a47b", x"c51197552f7a0378");
            when 21692046 => data <= (x"616703c68124c559", x"8f9f4fe6f19d2dd6", x"328f89fdbd057f53", x"846b29f5f257b977", x"44e2ff4257cbbaf9", x"dd16bb9cfb50442e", x"03285891f5871069", x"d5393746fbabb2b7");
            when 21058686 => data <= (x"2f1d57f67470ab25", x"fc63a0ab9eb338f7", x"d9a68e1732873dbb", x"e900c224f46b97c1", x"477f6d06dcd99b57", x"530b1c3af211c8d3", x"d304dff9518473c7", x"52384e7075eec278");
            when 33146274 => data <= (x"2499e3b68ddcdaa9", x"4260d617e52f1f5e", x"476873a6bc468a84", x"b9237a45f21bfd62", x"558f444a95630845", x"036be57be43be7ac", x"fb0427c4a8869935", x"8e8a335beeb07e3e");
            when 16396238 => data <= (x"7f56d1e834b940d1", x"4de750f6fa53a522", x"74d1eed4a1a69599", x"030e26f59ba8e084", x"ce4fb21abb0193f4", x"d1a34c78ebaef5d1", x"b53719866e12673e", x"afb1fdcbcc90bf00");
            when 24170988 => data <= (x"17dbe16249472f65", x"956fc708c57254ef", x"261d773ed299b188", x"50e2f06f63d3cb19", x"9587009ed9468ccc", x"fd06ff688c4b1366", x"2a6e1680c209c173", x"55e53024944f5f47");
            when 9456268 => data <= (x"5a74888558e73bb8", x"11ffe6c8f353f9c6", x"6aba9a4ddcbe2c15", x"2f8a0fb2f80d46c7", x"fb159e9b8fa4396e", x"4cbd5616e525f35b", x"5e439ac2e09fc3e3", x"69fd30df89071e16");
            when 29855836 => data <= (x"d2bce5fbd2f64c52", x"94661e4d31674cb7", x"9d799db583689259", x"0c28cc8d91301030", x"d496fbc0e695a591", x"16a2408711bde646", x"9e6707347dc75968", x"7399050807fae770");
            when 11592113 => data <= (x"c496531fc8a4c8e8", x"d926c65e9ac693cc", x"cef15c2d8396b219", x"539f8c7a1e2fcd2d", x"4ea4561be61a52a9", x"21622d3dfd9a7ea7", x"d1277dc7180bc6e9", x"b7e8788b19f7ad98");
            when 18726289 => data <= (x"1f2c20bd5c6a1a2b", x"bf074654186a2b79", x"16edf1db05520293", x"42e34d6c53f00390", x"738b195f2ffcf8e8", x"42c6b4248c943a14", x"bd810eb11a9c8abe", x"0cb3ae0b2e03b264");
            when 31535160 => data <= (x"d7750adad7b22db3", x"6ad116dca448977e", x"80a9d8fe8d7798f3", x"0abfabfe0fb818d4", x"5919b12cef2f6f71", x"88b76fe153b1be75", x"a078861167e0a8f8", x"5aeb419af616fbd7");
            when 23286534 => data <= (x"5177eb6520ee5cf0", x"73d4ca40a5457b84", x"0d498ef3eadf04ff", x"6d03c37d118eec17", x"1f95c57de10be4af", x"9fb24538da6f4298", x"8bb8c8f1a949aa78", x"4591a9401ef93e8b");
            when 13730449 => data <= (x"255d91fa9c4ba2fb", x"303a2100f275e482", x"a340327d3868790e", x"5c9f97ce2fa28051", x"b92c6056dbc206b3", x"770b3497fc454e1f", x"513563c0a4e507c6", x"6d07e7ebe3669bac");
            when 8552310 => data <= (x"f5a9691071627999", x"0ac562b197174267", x"938cbe646c728f3a", x"040eb23501f32d66", x"6578a398ae827190", x"4eb0a699cf1d5b1f", x"7e65a19bcaf66bde", x"3ff6327715b99546");
            when 17146902 => data <= (x"c9c52d0b2d0e6842", x"e32dcb14db0bbb80", x"dae321016500d407", x"3ac95adbb7913c0a", x"a2c1a56c992ef744", x"6ee17bb87d8b5b52", x"f692b568362d42e7", x"6743f0d919758026");
            when 13442957 => data <= (x"e880062f04f756f2", x"c92a4b526900d6c1", x"7fdd5d7a42255c2a", x"161c1f9a78ef2bb7", x"b874edaa6ebd1f30", x"4d987f9eb7cfe5be", x"a9f97cde31fe65cb", x"a7418d7a6d9e2171");
            when 29044408 => data <= (x"8028fef5436a7812", x"8911b575fb686ceb", x"bdec5307f4a390fe", x"03d1f318bc733a75", x"842c45397b337728", x"6fd8b780c86cdb8f", x"2060151a7fd7dc32", x"afd0c4580bda07af");
            when 528626 => data <= (x"57fbd9f0f60e0df7", x"8b7d0db5dc274393", x"1154f1c58fe3f823", x"f417157d89394983", x"a9efd1fa0bd40920", x"9a87792b0f6002d3", x"27fa4f28e767fbf0", x"548f6a618015261d");
            when 19129837 => data <= (x"6ee3571ca521091f", x"19ea5ac44cd6691d", x"b4477bd5602178f6", x"325f2779d514ee59", x"1f1cd0ffe3169320", x"1b718ce4d89ea20b", x"6571be485fdcad69", x"0f04e9e1f71ec2e5");
            when 16767280 => data <= (x"bbb6bfedf44df764", x"17fe48d781fb58be", x"336630ac8f2814b5", x"0a004bc87d55f141", x"e6eefacb33c22b24", x"03956e5d84877750", x"02d7518d45d2d507", x"7bb7f0400ab23d78");
            when 7687955 => data <= (x"871ac5ba7545c83a", x"e0651bd35949222b", x"481b687436dd929a", x"a8d4fb397d3c3320", x"f00708fd2fe297e4", x"a88bf698f1022f77", x"ef03da5bbdeafee4", x"ca4e446e836df6ac");
            when 1691311 => data <= (x"59dbbb7a32210dd5", x"fbcd9c76a0d98bf4", x"4ef0fbf342ecdde6", x"aebd5d782d53a215", x"030014d6a745e6d1", x"e123ec1cdf2f2839", x"95a9223ca089a221", x"e900209eb266b655");
            when 16156470 => data <= (x"2466c8d98a646a98", x"39e6ebf934157a69", x"8894a0af7e7cbc6a", x"a09e9cdf13dcf656", x"43e097a9a9d769b2", x"a9d388d5a5658e1b", x"943896216db42944", x"c623f989a6d1169c");
            when 25998335 => data <= (x"349a56afe8f95c07", x"2c90d9320c335f4f", x"3fb70c8e6304792d", x"f00d9a59b9245413", x"635b35adeda5d31a", x"9bd2dc5fa07edace", x"892e0d90b8acd0fd", x"c5a6dfe9beeae333");
            when 28934245 => data <= (x"230e97b7244f5051", x"5e97e0ab4bbeaf18", x"3eaf35354f7f6006", x"e6653a1c936f4220", x"18b1ef7912b405a5", x"a92aca00f17558ee", x"e9f35e06f0297552", x"ad4a3ed0dbe3547b");
            when 3034245 => data <= (x"c53774904feab753", x"ddec6ad7f02ecccc", x"7340eda818307356", x"bc5d79dbe7c56189", x"216dc71d9ea0b63f", x"8163781fad294ade", x"19e45fe994951af9", x"7b5b095c2a2fa597");
            when 31639458 => data <= (x"ae55943a182c24d8", x"7f2950f8d75caf20", x"fc28b24c4048ae87", x"8ca4a3fdfdecc57a", x"6a5c0730e7560d91", x"86eda2258758d2ab", x"59803580590c9f57", x"3b5c8f1f109a5ccc");
            when 6674099 => data <= (x"c3be211d226b95bc", x"fce5dde0ef389fb6", x"5baee03497a32544", x"985cc8d945ba40b2", x"82a8ecf69cdcc9de", x"c3f34e6a82fe8d98", x"a464771ca709da10", x"2c891aceb455f23a");
            when 18580574 => data <= (x"db848f2519bf0695", x"a6e81ef675d7286a", x"2af9cf39899a4c9f", x"e67eb13abd4015e4", x"e0aaf70bf208824a", x"63539b3b74b42cce", x"911051162d5eb990", x"00678838a438b856");
            when 11695361 => data <= (x"9c95eed37be07d95", x"6ef7053cdfffa7bd", x"aa5711d73c4cf32e", x"ac9cc879a87b1797", x"e1a6308c3a64473c", x"3ce13b46bafbe1a8", x"64fb956ad4f2d3f9", x"09c74a74ab655b57");
            when 8401386 => data <= (x"1011d08a91eb753e", x"0454f2f8204d1567", x"16cc1c42b8e76760", x"8b600c6d056b8b88", x"496dd0af0cd418a0", x"aee0f59e792c5ba4", x"38350f89ad6ddf26", x"1c47189be3f2df75");
            when 33639595 => data <= (x"bef882f2f4865db4", x"b2cf573b14ecec63", x"72d9faa282e028c9", x"92498c99704fef6f", x"c0d8c5dd9c4a9522", x"d305cf84817af2ab", x"4c91d9269b1f3f40", x"036685de51310c36");
            when 24319677 => data <= (x"34f42d2c0b38bc02", x"53f9fbdadf173918", x"e9870e0583709bde", x"347777725551f4cb", x"12098c7225d7706e", x"efc0a5f2b727e740", x"2ceab828439dc0ba", x"074376e9f276b686");
            when 23566856 => data <= (x"21dd5ed866e213bf", x"6d9db17645e7edc7", x"8931d10c46f20199", x"e31478b51e4b1a0f", x"93d0365591367e4a", x"db624e52669f03ac", x"eb0dfaa518eea649", x"aa36c2c45e0414aa");
            when 20677035 => data <= (x"fac4a033472b1581", x"c8be021cd31f83e7", x"27c1f3e5d60998e2", x"1c3fa483630158ee", x"aaa68d72d794eb42", x"de1c58a111c0e0c9", x"11886a32d90f8b98", x"c20376d9dcc83e66");
            when 20738343 => data <= (x"fc3eaf5f190b4bd3", x"ff98f19c77a30048", x"cc67704ae3d1f5a5", x"35545222ca09ffe5", x"8a8c7762cefa6a6b", x"540cf0924e637e39", x"491d6d004606cf81", x"fbb6d4312b5ad0f8");
            when 2248283 => data <= (x"ceb30bb2d84aa135", x"062b5231567097f2", x"c77beb7dce35c319", x"d7445c22d47f7a43", x"b5570025e85eb727", x"3d10e042bcd70fac", x"016bda3bea98cade", x"2aa2501b8ccd1190");
            when 10740106 => data <= (x"ed38fd52078d82b7", x"3fee0863fdeb8d11", x"99e2510f928e8ea1", x"70dc3e3084f4fe57", x"a233b18918be3733", x"6e04eddb91b39cc2", x"d6242baf99006030", x"31d5b80468a31313");
            when 21221111 => data <= (x"1ec127383080068d", x"f40561f4f6e3241a", x"8144aa5c53efbbb8", x"c48edb3bec9874a1", x"d454766e38132bcf", x"8482504cc4941da7", x"1552d4e131078ae2", x"491e7c897dfc6c87");
            when 9697626 => data <= (x"bc80f4d32b3f83ac", x"2163f3b6bb412de2", x"21e99044f5e9b30f", x"f55ff19e59904a93", x"df547775fe85c6a5", x"9fb72512c61413e7", x"553ff8391075aca4", x"93ae312a80687de1");
            when 7193282 => data <= (x"bafd5da59c67a699", x"bce2df0fde46a0d1", x"19b3cbf7c02f540d", x"112dd965d1990e94", x"99a131205f140b02", x"dd4b236ed3509aaa", x"b58e1a5186d0ceb3", x"6d5e203b739b9dc0");
            when 658133 => data <= (x"bd1d9b781c0494bd", x"7f6f6938050deea4", x"b161aad3fdb32a87", x"697444ea081c6529", x"54d83679a56eb6df", x"e92d2cce30fd1d11", x"76d56ea314dad4c6", x"904b01c4290de66b");
            when 14626540 => data <= (x"d0dd194dad97243c", x"e64fc04d1eb0a754", x"8c76cdea82c863c6", x"10dd9f399158fade", x"da3ce6f2b8aed6a6", x"ea104c434368be34", x"01e1cd413ca6b6e5", x"0b864d67c576e608");
            when 4775768 => data <= (x"917f6c3b12a09144", x"6b0352d9ab3d5fc1", x"1d138ff8b0b11aac", x"f49dcbe0e5c1539c", x"8ac5e50809bd40f8", x"592f8267b37aa714", x"2da8c6af982ff884", x"205fd95cb7070c78");
            when 2522409 => data <= (x"4dc0a1a2a437b10f", x"0773271749aa67d2", x"5ed4de6455113b6a", x"c837a398cfe62cd6", x"540d1add6ba30430", x"00782ff90cc4e86c", x"1094485f0ff17856", x"ebc34a991a13028c");
            when 18616165 => data <= (x"30aef6c12003dba0", x"0b73fffea718d949", x"8aff50eb685f9e9f", x"55b0193c6f2ff8f7", x"4ad54c56a6d0ba1c", x"dd99ef0cb0c34475", x"ee2107dbf43592b3", x"1ce35ae833dcbf60");
            when 10942959 => data <= (x"796bf7e4125b22cc", x"3acfa8a1e87b78f6", x"ea91c888abc679fa", x"c8d4d347c9b8231e", x"4a87fc01f3d3c3f7", x"b67a3f716d12ab96", x"78cbae6604c27601", x"3280114c3a8935a2");
            when 29262718 => data <= (x"4ab83e9e623f9017", x"baeda56ab14ddac3", x"a3ce18e973a0672b", x"bc73350da829f4e9", x"2fbdf5b39ee16585", x"789087584428c5f4", x"00ac7bfbfe85dfa7", x"29b0a9f0f5915365");
            when 16701361 => data <= (x"8439a80d481732c8", x"2465380317719627", x"4027e429456e48b7", x"360a272314d44af2", x"8f84a872ab15523b", x"4357afdd0500796a", x"b4621d66b8fa26c2", x"3fb7e17d12fd2baf");
            when 30054894 => data <= (x"11de2db434a04a5c", x"dfe16c1a38da3a5e", x"f31e7aa7dc31b3ac", x"a1a526ddcf99e150", x"47cf0cc76db8f15b", x"ac1a3ac869029bcb", x"a65f6bb456f13afb", x"6e74e7fa3f247767");
            when 7313493 => data <= (x"bd28b4a6fc1d435b", x"78aca5670d2dbdc4", x"c4371fb114c154e9", x"61ee4df9f7c9cf3d", x"bedc0404438c330d", x"56279c98fbcd6d38", x"4455ff5e2743ebe7", x"fe5dcb3a3a1fc06a");
            when 22013184 => data <= (x"ebb47a0b94ec6118", x"fa927f941ea054e6", x"fbc3e6e1ddfddc90", x"ba9301fc611dbc77", x"ab5bb91b2c4d3a97", x"93145b844c777099", x"27525490eb6517c0", x"ba756564090cf4d9");
            when 7825974 => data <= (x"3aaabf693db47bdf", x"50d5bb6bbb142a51", x"51e21e807b3102b3", x"1c2cc1727eebcb8e", x"faf6a0c9c83f1bd5", x"6354fbda46b03127", x"552aa7e30886b564", x"d367a11534e5777b");
            when 26713398 => data <= (x"11516054a93906c5", x"b40d42db74a4815e", x"647548053bc6b560", x"5b9beb055ef61e64", x"5851fdcaffdd56e8", x"29b366db8c34d2ea", x"5ec02bc119702e8f", x"7e3266de9a8f3638");
            when 781019 => data <= (x"5adb0165f1fce32e", x"2f591eb1bb3bf07e", x"91e66b6173ecaa78", x"42a51d3c45fbd142", x"356ec93a2e5e2b9b", x"2a07e602d0492f12", x"840a5aabcc180211", x"ce169b9370df26a3");
            when 31590520 => data <= (x"584bf8aa4808e429", x"4577a7c00a7c9239", x"4d3e86fb3a476d34", x"086cf6a579dfe870", x"592603fe76412410", x"ac04b739533f04d6", x"567bf0200fea7624", x"e5a7a62746267656");
            when 3379410 => data <= (x"83628909820f8aa0", x"5c45d377d52b46b9", x"3cb7f46d3156d221", x"ed045e9635622f2c", x"cb75d4831586deb6", x"05be236cc90a6305", x"6cbf1b7b10d93deb", x"635f0da9bf6ba7c0");
            when 17233007 => data <= (x"b008db30a6e01023", x"ca4030c72d3bdf67", x"6c8bcb6ff5a38f9c", x"6d175fddd1681747", x"192d1a00b0fc64f9", x"ed56317734f8c094", x"6007f6fb01abdb94", x"83c87955ad0987f2");
            when 10185285 => data <= (x"b3ec86e9f33dcf29", x"327f7d203e0ac12b", x"a6a78de1883e235e", x"56a678f93de0b3d3", x"b4d898e0d919237b", x"1180eaa0c5a1b3f3", x"4195f14ac979113f", x"2c6ced41f0fa544c");
            when 22835641 => data <= (x"b716a4375d909c85", x"0beaafcbbc51befa", x"9384c1aeff707222", x"c102a195d2f4d1f3", x"15070ad07e97da19", x"6950dd891426724f", x"78bae92ed6933851", x"39779e151d1e6b77");
            when 6273079 => data <= (x"e2ba99be25c97550", x"60c20782c386c310", x"4fcf39a57a7a3953", x"0631988561301f83", x"087c1a46fb3907ec", x"a80e29e58ba50d00", x"6716235286e3c1ed", x"7c1050cd5cf76a85");
            when 3974557 => data <= (x"3e260e83b1d9c756", x"2f5e8e408c18ea50", x"a8b2956dbf2b429e", x"1f0603d4ca542d13", x"ec2a2d982e175ddc", x"e9a36b3353638fc8", x"8e8f6b893ee52118", x"be8763c88c253888");
            when 5210458 => data <= (x"fb6f5b4540375a0e", x"409b69e1142d0328", x"a5fbc55f9baef63e", x"81610b728defcd0c", x"71af205687054159", x"18b86d70e2e5cf59", x"5b05f078ec7ffa39", x"803f7b50e27f81f3");
            when 32342328 => data <= (x"eef44ee0bd762b6f", x"214aedff464aa453", x"0d13eea9a74e80fb", x"a5911bc15283c5fb", x"0e08170015a2dd71", x"56238f5c18aa93bf", x"36c17e4c6cb22e69", x"20c2f5de2ebea60b");
            when 32350674 => data <= (x"b405514a08e0b688", x"98b7c90234913fc2", x"07d73fa4d006b0d1", x"8500b802446f512f", x"76b92a53ec0d2b21", x"7f875a7e905aa6f6", x"6589f7ef5a74ebc6", x"8b208e0218003103");
            when 18768235 => data <= (x"6700170368f778bc", x"a04afa1fe01be67c", x"7ccc989b0d8ab8d3", x"38382394c5c24509", x"580d28b2aeb45961", x"547b1ce9c75d345f", x"fae337d36364c2e1", x"77d336a4ad628001");
            when 9355766 => data <= (x"c6c8dc8095fe5f14", x"88044d4b89e06fbb", x"35f9d90a58dcf97b", x"470aaab4605cb381", x"f1d86587fd3987b4", x"5885b63df2c22131", x"d87e0791d48436c9", x"bff9e45e8fb79367");
            when 25653561 => data <= (x"a8ed77913df97430", x"fe7df553739917dc", x"901c64b7198c148c", x"5533172fdf48c609", x"1e2f55a41f89183a", x"9ab0868038659cb3", x"4457dfcabcef7be5", x"6a5839fcf162ef23");
            when 23609097 => data <= (x"ee41810fdd508c34", x"f9d5d4ca611b62d7", x"2ef1d1173da50e06", x"9a63ad39b08ac586", x"ed6be09f97ea3ddf", x"3682d4408da144e7", x"a5879596b8e30dea", x"1f7ff2bdd0fc4769");
            when 17237343 => data <= (x"dc74e2a75e068acc", x"bba43a9fe5449ac1", x"f0c545eba8dd7bba", x"c7a6ea0514b5fb90", x"ef2673dc8a940574", x"ec47f33c72e04ab5", x"0427f9ff6cf179d0", x"a171042cd5f58d68");
            when 22726403 => data <= (x"1a79da3403ab30b2", x"89582e3e746ed9bd", x"f5ca2ae22fdcab77", x"6d85610620fec6f8", x"7c430c8518ed2030", x"3ed172830a60c847", x"c16b53f1402524c1", x"5a59cb6d0329ea5f");
            when 18747572 => data <= (x"f1c60050ea7bee59", x"93a97fbbbf3dd155", x"b8fe6e0a073db1e2", x"b4791ece111bf975", x"3273e45e8d0c9d11", x"fd55811b09d33515", x"2e84abc41f52c1ad", x"31cdf8a57e82091b");
            when 4467452 => data <= (x"8d4ed67680cd6789", x"a2176b6fad7a90c0", x"9eb564b707aac2b7", x"5386b6da618a9d4e", x"645ad067c26cfe3c", x"85a9a5f14b099192", x"ba1356e16eadddab", x"07e152b362b2f398");
            when 25914001 => data <= (x"1e06d29459825345", x"a707763de5a4a416", x"3bc2fe22db97b353", x"a5d8abc271e0362f", x"015c5470a7f9d0cb", x"427f59e5dfa8ac58", x"6d4220cf09fa97f3", x"faa1dae27454baec");
            when 33080377 => data <= (x"dd50242420424a6b", x"6c5645c8db3756f2", x"049ac8b98a1204e9", x"fdb3b22591e625b0", x"8960be774c03002c", x"521f7bec17a49ac8", x"d45fad94350e74ff", x"2c44495068d9def6");
            when 27693478 => data <= (x"6ad807bb8cb8a3e9", x"95c7e8f31ed5a9f7", x"98713419a059a691", x"d202d54bbe78afb3", x"c775f1d703d95b01", x"a1cffe4962a548f5", x"84fbd994c6a7071f", x"ec9eac0ec4837d4d");
            when 24406465 => data <= (x"75dc8d6fdf637d16", x"775bbdc6e1d047b5", x"229c9b4e88d266e9", x"952a40fcb94949d2", x"f11abac44a73e3c5", x"85fac50102af5a74", x"ac56f5033f5bc328", x"d40434d2014eb61c");
            when 7074899 => data <= (x"d6fca47691f1c2d4", x"20d38daf1d179160", x"05a6d89c182155a0", x"0dbd6982ac4bff92", x"bb305e5537357f9f", x"99b0e37aa335727d", x"f3506d13fe27fbfe", x"dae728906e5c875b");
            when 21160732 => data <= (x"1ca7f5b28edde42f", x"c5e96a64916e2c70", x"1d7bb504e31c1c30", x"6f05a191f42783b2", x"f3124ae20e8c7d54", x"ccaab430bf19541e", x"7d05d484521f731b", x"2fefa4931d065116");
            when 10750863 => data <= (x"c76156554fc54150", x"f5cf2e1970f9fb9f", x"22141bfc715c1b75", x"0a7274eeccd3d692", x"42c026207bc7d115", x"f49825c30b7bd9f6", x"8f1a27f632c93ffd", x"a667a8e73ab7d6b3");
            when 29834148 => data <= (x"e40fe0fc5deb99dd", x"5c0b5c56a3df068c", x"9bd344f32af100e8", x"7ef55d6cbe94bffe", x"6d827abd6d3b8da5", x"2b9fb65e532c25d9", x"ff0fd540408dbcbf", x"cb107b40d2be199c");
            when 25910108 => data <= (x"630afdc1b0e48ce5", x"987d536e89bd9dc0", x"b8b748b5a2c8b777", x"350596d51d1ae8b0", x"f9ba5d01656b4cab", x"f0a87b6a604aaa64", x"f9f4249acde7a541", x"258c4341bde82724");
            when 23816950 => data <= (x"b2946af68d2abe15", x"35f506e10cd4c8a2", x"dd053ba20c564629", x"4663df435380a018", x"883d8d856d7d349a", x"2d0d3194481fd8d7", x"d8d14c82ca34ee48", x"f7988e46148e6f62");
            when 26870133 => data <= (x"de3f7da92a4d0d5d", x"1eb7f6b4bcb8ae9a", x"f1cd198e0569f602", x"37f598da1a4af0e4", x"f491b8412660c241", x"84010419dbc514d6", x"8da413df8b0d8691", x"864c1cf8c062e4b7");
            when 9471801 => data <= (x"54959ad315431070", x"131a0c59344c2e14", x"726cb574cb6a6327", x"ef536d66d86d39f7", x"c16f6d9c79b29660", x"a363ab0b66c0e607", x"c9e5501e93e2cac3", x"9e1088d066477b1c");
            when 7898327 => data <= (x"6d306d7d675c6108", x"c8fb95ae1f1b6f20", x"c54f00d525567d16", x"1f4f2eebb123cc56", x"93d4fa52e9de13fa", x"6e488d83f7d51fca", x"a2dec274a4527fbc", x"483366b547bffd73");
            when 32889145 => data <= (x"a0fd96250e98e817", x"4a1268c655d54e9f", x"798b50febb489d31", x"6451e8f15de8297e", x"7218ade278fa7c10", x"f4d2abb3d1d0859f", x"6294b98721bf4b99", x"48b8fe24eb236d0d");
            when 5989323 => data <= (x"0ebe0162037faf25", x"55716a1648c8031e", x"1d03de23d1b92895", x"c455e2ec18b49887", x"5d52123ac0a41823", x"fa7b77cace8780cd", x"d852961a9c1a1d88", x"0b3dae810a0a17ca");
            when 21955595 => data <= (x"228d05b51a976860", x"e698b617e3a0e4df", x"56a7215679d14a85", x"70bbe293b2dde416", x"c41049e618b42c1f", x"20cd9e5de0433a1e", x"b2ccd2a67a468195", x"50de1dbdebb4c7fb");
            when 18782091 => data <= (x"3c06f7026096a3fd", x"6473abc7404c44ec", x"9a501dd4736a89a9", x"f3e16ed942a61c23", x"24284572357fc0bd", x"efbe38299e73ea72", x"32600e413533ee4d", x"2933e67a8a43d6ba");
            when 2672502 => data <= (x"6d41f85e194ede99", x"1c09d2b87fa51a15", x"fd0e2408b621c248", x"0d183686d0795f88", x"8d8d99dc101c4567", x"28e538916cd3a38c", x"8f9321eb97543b62", x"cf5d0704983469aa");
            when 15239035 => data <= (x"3747a8cedc05a319", x"f7ce8505c9478a80", x"c4fe5ebf7f676145", x"e275aadd4b226333", x"74b6660911018478", x"237145998b092d3a", x"400d9457368a322a", x"f3a1dfe1068c215e");
            when 30864643 => data <= (x"89250ad75349d3ef", x"193c9d135f724e7c", x"06202fec9cc85c5e", x"b1d51ed77f4c0c9c", x"7d30712f4b888e05", x"2fc16a2655bf0820", x"62f4b76e886879ff", x"2713b5805ffbe3cc");
            when 21150076 => data <= (x"426ca27bfb860315", x"c5e92ebfeacfdb31", x"0d2c95b8b224633b", x"9e3c9c0f9ead1b79", x"2043aeddf73a5b8f", x"f153d186fad244c3", x"1e3884ee4517c636", x"535342c3f5e3a2c3");
            when 1618892 => data <= (x"d34f8ddb663cac3a", x"5d7263c2a1cd1154", x"2ad5a44d1933f3e1", x"945a86f7ad355f18", x"f0fbf994c4383264", x"1a9b23a19ab28f3e", x"e2631fccee9655f6", x"2d4b56b52567ac41");
            when 15336861 => data <= (x"552c10c4d5a7fcc5", x"11f4c41bb1b3785b", x"9da66203c6a306db", x"153e8af353ec5a69", x"91e3d132ec0ff94d", x"37bddf7a53cafcce", x"4616a535fbf0da7a", x"ab9bfec512b2a1db");
            when 29874315 => data <= (x"60e0814e89269b92", x"952a3b049f0b3daa", x"678cca26773caa73", x"e0d62ba766998b09", x"308eb52d3ee3aa2f", x"bd1f3e4dffd5482b", x"e87e41f3b05e5268", x"b3effd9cd4b695db");
            when 26349504 => data <= (x"2b1e4c87375dbfb6", x"5637244bd483fd36", x"e80ce2d66de3eebf", x"aa025c31babbd0f3", x"0a62b4e3dc12f1bc", x"8c8f94d2c6d368fd", x"3da59adfa40bbb0f", x"0a053a6e21b86955");
            when 24453130 => data <= (x"bc4b6f6f0b80152b", x"e8f936b9845ae438", x"cc2d9416510334a4", x"904ea4a8f9e5a722", x"91f1e47aaba6f75e", x"ef7daf42ae5a0018", x"3049556b09d97d64", x"2d906f267cf3ae71");
            when 27505867 => data <= (x"4ca312a07be421bd", x"dffffb86b0b0936e", x"cc6de19e1ddaf155", x"9b52fa8120dfeb33", x"a46c8761a541be7c", x"da9bb5eda832b804", x"70571279509a2727", x"deb8ee4c8c6fc592");
            when 13310529 => data <= (x"e6135ccbcc3e0c04", x"1662508c45e9f00b", x"695b505d74a0835c", x"21e45a71080557d5", x"3ead7b77afafbcda", x"3051c4957da67ffb", x"317616bf9d3ec236", x"34882a5305badb9c");
            when 4567963 => data <= (x"7aaefcd3852a1952", x"fbc8e892c2a7873e", x"b890b2a6c1b11b8c", x"fa869aa99be523e3", x"82e4ffc21f3a427e", x"e8a6081372d76605", x"c83c190e81f8b185", x"14567cfa1bd6de96");
            when 7432253 => data <= (x"b82881cd8aa47603", x"3eeac7e4f4e4f546", x"30d145e41293b1bd", x"12aa9afd34939123", x"591b12a0b51f9080", x"5bca2fe6a22a7c02", x"e973cc7e48996d63", x"e2a20080b3fa4d93");
            when 24054082 => data <= (x"4b59e6f092d679ef", x"d11f241b9882d9e4", x"af50a03beeb22173", x"636ed1923e653bc9", x"f3aaf152d9002052", x"37badeba9b2a4d1c", x"4a80eab6c5f185ef", x"ff0f72c2fb422fa5");
            when 11823085 => data <= (x"0918dde3fd32503a", x"9ab7c30835223f0c", x"14bb17f13efc10b2", x"9716b78efb04a156", x"d28d7fabff3b77c1", x"c5ea5479b37c8f27", x"2d84f61296517484", x"0d1613757bfa46ca");
            when 1148726 => data <= (x"12e9354c87b53978", x"d3bb659a47a8c932", x"1ed7895684ac1290", x"b5f3f1aa8c17e4bb", x"858e342cf7993558", x"bb3554eae8b4bbb4", x"ed01c08d85e5a3e2", x"589b9886662e6b1c");
            when 22952813 => data <= (x"aa9de8fc1bd879ee", x"4c4a3351e75d6adc", x"0d20bb44e7320de9", x"aa14036720b455e2", x"6f8fca77fd5107b4", x"0ab4d78c6b547706", x"0c211e4526634ac9", x"086e30618208c603");
            when 24236128 => data <= (x"fb3f8aa4d72f0e7f", x"15366fbfc3e83659", x"34f42fba970559e8", x"e800d24a073ca407", x"ff7576537f60d3a7", x"bc6b0c5f696ae14c", x"bd0740803d3d1fc4", x"04b830afc7b305db");
            when 33778134 => data <= (x"5ce330ab6a3a2ec6", x"7c9cfc596a91b6c2", x"e7864e9b6537a7bd", x"ff0a0eb8e30073b3", x"8ffa4e6aa6829e22", x"573a668e5db2df23", x"9904af371af7de8a", x"708108818f0b4ec3");
            when 28166587 => data <= (x"f7b77420a828592c", x"0eba5fa718872e4d", x"3c05c61e444899c9", x"930eeb97f132840f", x"c1e91cd227ae7d68", x"5e3b649cbf16d4d0", x"5fed7f9359cf67c0", x"8ee2837ca132a5ae");
            when 20112506 => data <= (x"049778cefacd7554", x"d3c1a5034287bd48", x"c1218797700ffc34", x"cd7f7f451318c247", x"e29adc048433409c", x"0e84d94d068920b7", x"ce99197869a5a86d", x"4e831cc7c7288040");
            when 2374766 => data <= (x"46cfcdc67853773d", x"15e6aad0bdb06682", x"97c6366593ecd1f9", x"e1939954fa06610c", x"92f41054049ab030", x"ae3378c79f4a469d", x"e7bcfdee82342ab7", x"cff649e4dd8b2827");
            when 32111617 => data <= (x"dc39e8c07076c28c", x"0ff2be63799a6004", x"4eb3e4b06f147599", x"29f0ece19aeb3587", x"990fc6f4228f88c1", x"ece53cfa149518ba", x"e6ae02ea97f528e7", x"a8f0e0d2fe5b837d");
            when 15095551 => data <= (x"d72141517da466f5", x"deff54b192778619", x"767abd3402138531", x"1c89e4bc0563663e", x"b908dc68f6ff6fa8", x"f2897e482302cff9", x"ab4058540b311cec", x"c6af5e9a262f33df");
            when 20509280 => data <= (x"615616dac6a1e97e", x"02f43a319491de9e", x"64141a3051883cdf", x"18aec1bf92424cda", x"ddfbbdbc65e491e7", x"b99a442d4ced36f5", x"588e704dd9258719", x"f683ed911f2a39f6");
            when 1900315 => data <= (x"7da72076b65eefec", x"7d6091b3d7671be0", x"4e0c6b3d7336834f", x"9e9176ec548baad9", x"ab117f8cbb3a6903", x"9c7ab697caf41f18", x"a5c5807c00a02828", x"dbe6fce87c4a3bd8");
            when 10171813 => data <= (x"35f61e4f4b8730b5", x"b876d43a4a55596f", x"5285e8393a2cdbcd", x"f90dabcd263568c5", x"5f6ecc32fa5056f0", x"e17906602340c35a", x"c0cbf260a5796939", x"3682fbe7e26bfcd2");
            when 32576131 => data <= (x"91715254759a1d9f", x"a45ad9398d7fe7bf", x"3c833a055fe9a936", x"595e7fb69eef6532", x"bf460acd9b1fe706", x"7a6e8c7feec2ccad", x"98a131ca5b33c367", x"9a8239fe2ef4eafd");
            when 21293876 => data <= (x"a0af4e8a35e9f4ed", x"bc0c6834d911ee2a", x"84cafb04a28e71a4", x"af5a89862e3e51af", x"f89e25250588ad0f", x"0a25d842922408fb", x"2aa065049acfbce6", x"bbaeebe3eb957aae");
            when 23134554 => data <= (x"15be3e79b10859af", x"0a2b65abaa57a4a3", x"91dc95c6bbdc12dc", x"9af8f53edea2f342", x"aa8f930709123b89", x"b3d4b00e6c3c27f0", x"b98f68caa5222ecb", x"42a95c1864fcb63a");
            when 6389937 => data <= (x"e448814bef4c6dd9", x"175d6f46919d222d", x"29c9499166ac7715", x"c430d8b30b58c5d6", x"b9c251aa127f8648", x"eafb739ad91e62b0", x"7a09cfb959a4a2e0", x"aae6a9d6adde4954");
            when 31554546 => data <= (x"e9c55aebe89baa74", x"345b1e656651d20a", x"1d9a04714589bf82", x"30ca5fa7852889a9", x"92233a0cd7e31229", x"4b68282077ea7b5c", x"d6c27589f0451ec6", x"c33b081221e2a234");
            when 17940683 => data <= (x"222a0caeff4ad029", x"95e821dee35e94da", x"87a637b9078085cd", x"b6598ca298640e93", x"383620a994d02b76", x"c2cae988c8a850f3", x"9403e9a1475e3a78", x"90e1fde0d0d63581");
            when 24550957 => data <= (x"10512efaf3d22f96", x"fb6b21f23ffc703d", x"723b8b8b79d2df7a", x"195e3065931dc77d", x"2299ea4bfb2bfead", x"da4e426b10c05377", x"0256e835e954c172", x"d3e91d0009cad90f");
            when 29698922 => data <= (x"853a0581f6dd55ea", x"8d85ae8ae82c95bb", x"fbd4319e06e0ec2b", x"353a79d1eaa133f4", x"c319551c070913c8", x"86584d0dcf93acc9", x"72432006ffe91d4d", x"535585a7c92e5805");
            when 9698102 => data <= (x"a155730240ad15e3", x"9815a81e081a3de2", x"0d9a93387a947ca0", x"d9799c9fc5663d13", x"85122178ab0df057", x"17c0e780d9e47d71", x"ee8e1426128dfaf1", x"0a43ea14a63b58e3");
            when 26497942 => data <= (x"2e30c19110a50cc0", x"4383041dd4d5cc9b", x"8998c1965323c401", x"ab64e5656636ffcd", x"9bf2d70869d02755", x"d36a62067cd4e700", x"b6e4bed7dc0c4958", x"bb508c3d61cad798");
            when 25649986 => data <= (x"959230b955c1c970", x"c3665f2c9bf1623e", x"b853c57f1b9816ef", x"55c5cdfa1682d026", x"0f60db564e0f0c62", x"6e7a9bfc8ce3a92d", x"e694327c1ce7bd23", x"6b2c28fa274c9c0d");
            when 24869713 => data <= (x"0ffdb8d6b4d149e3", x"6b276aa653bf5a69", x"4960c0b89c38b673", x"8921aeaf027f59fd", x"e4c2b00c162815f5", x"486ac4071a4ec0bc", x"96d23887d19714f3", x"49106174874a228d");
            when 8690772 => data <= (x"e293bc35d45d9deb", x"bd1d7c34010fe05d", x"636b8b3fb2aca0ba", x"b3713df66c0fc6d0", x"87353108067ae7ec", x"26f321ff53621c7c", x"fadf0b3dedcf027a", x"8de7ea2ac8186df0");
            when 9158037 => data <= (x"887e9b8c21b97335", x"cfae23b9fc135540", x"773fde64ee52f959", x"fa02d740e2d9ce28", x"e91dafa544635b8a", x"c2729d8212e4ea64", x"16c618b7b9d3ad47", x"523667e47e74d0a9");
            when 6310524 => data <= (x"4e4655775d2287dd", x"31a8286956bdabe3", x"c49606752aac1365", x"a5f2606cfb5ee390", x"94c9d4604e2e7889", x"3a3d011beb7465f4", x"f463e9b2b04fad2b", x"22a201585a96abea");
            when 17154427 => data <= (x"93cc95f632fe243f", x"41e8e44351df433c", x"449191c7a8bddc0c", x"6958254312c0c8ad", x"022e2672f2416fd0", x"d5fc1e80d4f3b242", x"6eb8e2d038d45502", x"87b907ddf072519e");
            when 19830263 => data <= (x"2d486f2c3e4215c9", x"4454ba299d2c4dfe", x"99efe35e26b1b781", x"42e6a530c3d6672c", x"4c6c23a61956226b", x"d76b73012cebaaaf", x"9cd6491ab0a25ef0", x"c2d22f8de6193921");
            when 30393586 => data <= (x"9bedc3a6248a39c2", x"cc37fa98fbec3101", x"f529000f996474fa", x"e63b418c200c66b7", x"3c76a1fe691d25ea", x"5e7a1a269a62f857", x"4e1d49db4b188290", x"6d28f729fe6b8b53");
            when 10464280 => data <= (x"dfd693e763efb302", x"ce53627ecba97cb8", x"efbc58ce72c25b24", x"d20e229d8d9c23a3", x"436f4dbc8817f52a", x"1ea8f4a87d595efc", x"ab102cdeb9fcfe55", x"98c199476e70a62a");
            when 22545947 => data <= (x"424de105d351d11b", x"c0641c6a57172859", x"939593044f747589", x"0ab8d4545a597dda", x"96165a961ca8ccd2", x"30295d7d37dae578", x"02e9a04c1fd45911", x"7dd1965366d200f8");
            when 30400835 => data <= (x"009b9de0d5d79b00", x"31cbf2668e731851", x"b5728f25955f85ed", x"2927dde59111d28c", x"0fd88e379fd92e3f", x"269af285d85319b0", x"f723272075d396d7", x"1898dd8d952f7a38");
            when 24376222 => data <= (x"eec106e9ee7f336c", x"dc0f4747292b0e34", x"d9deae97f3d82a52", x"d5651535864d7ec4", x"4dc43ba32080a4b3", x"1ec5c7357e1cae97", x"bb94b29befaa7134", x"c0309fc982dc3a32");
            when 3500538 => data <= (x"be8b9e0405947e23", x"f7daecf14abda4f4", x"2de5e4fc9f66dbb1", x"75e4b83494f9847b", x"ac42fc36da678a6a", x"52df2583467ce7fe", x"9f974d5b9a4e6378", x"9faf684149d809b3");
            when 21734890 => data <= (x"640ebb700ca6cb36", x"74784bb20d54c5d3", x"b8155d7c9a96ddea", x"84090b4b411e34d1", x"1829262664a3ffdf", x"5a8fed62787b33ea", x"c72a0ec5ddc0331c", x"372b6541c4d2a064");
            when 5545408 => data <= (x"ccfae5aa498f7be2", x"6b8483c7dfeaaf05", x"e7459da6cb47d0fe", x"d88914d0a42b17c5", x"82349fb4c7014b18", x"bdfb810656c93993", x"b37b78f6dfd185c8", x"400fe145f9d832d4");
            when 31596988 => data <= (x"bfc94ab1e29d3a05", x"c387fdd8a5ca04bc", x"93ea3c738973f566", x"fd692e7a0f7b035e", x"a291744598926694", x"b7ce54a48c484521", x"ced76f8c13bb993c", x"a6c57c641fdabd79");
            when 29864003 => data <= (x"5c5ddaced34780cf", x"109ba75798e4f33d", x"a8e04f0efa1cfce4", x"888c31c9db4c2bec", x"0400f4012671fde0", x"b98b17ebf4bb6265", x"d039167e719e9c69", x"59e015be64964a55");
            when 18521975 => data <= (x"b08586f5f93cb5b4", x"a28215a689ebd5c1", x"e625e8a0f6cc561e", x"2ec2444aac0548fb", x"7a62d1fd5247a03f", x"5b1a685a30e12fb8", x"d4d600a0775f2d64", x"63d6022086c17ab8");
            when 31531197 => data <= (x"a6667de5544a6d74", x"38c0e90346b0589d", x"f77eff2a7a6df1c1", x"580d22f2c816dddd", x"6dfd07bbd04395bb", x"2d58451f5fbd7657", x"e7f8365622a14f62", x"87d376ee2fa7ea89");
            when 4327479 => data <= (x"23287d40a8504cfc", x"0bca9af7f7f2353f", x"9251a5e461deedd0", x"56e92d9236ea66cb", x"d656874890c46573", x"0f5121065f0b4054", x"fceb0728abb82fd2", x"572de6290c6700be");
            when 31737817 => data <= (x"8ead6ea6754e5a3c", x"633e7ee492d22ff0", x"7e61edc7234d8880", x"c146ee74d8a01971", x"087b29b0da4fe536", x"597e6edb831dfa38", x"cac9240885d51474", x"4f9144fb3e76f100");
            when 12242129 => data <= (x"2ccd0bf3fba065d3", x"90a5acc6f56e45ca", x"707854a18e0eabea", x"9b35ac552fcee1c2", x"ca9993949dcfedd0", x"acfd7b0df474c075", x"a252b03df511ab50", x"05b7e6ee56dc7701");
            when 31330502 => data <= (x"29e7b79379bc33fe", x"c577c5da1e9cd106", x"2a0c1ae438d7cd52", x"9d6c3d72ba9fe536", x"d04c2059fb2e1e8e", x"8c02407eceab83b7", x"43d99ddd3d9265e7", x"4d64fe4933759455");
            when 20358401 => data <= (x"a63fd754d16240de", x"fb5d0644790f30f7", x"f68baa1f864d5c8e", x"af24fcffc897e36d", x"b6ca50bc4b5cbb94", x"1f19f130225a3e3e", x"2fce3bee77b68ae6", x"0ae13a30719b1451");
            when 6926707 => data <= (x"ab2907490b1843a3", x"b3da2e897857a9fd", x"5f4746e8168b0622", x"b1c878a4da47f4ef", x"3333d3bad0d1a889", x"b9ed6a9700228bfd", x"fb7fd94dccca0a0f", x"ec09212863ec035f");
            when 4822041 => data <= (x"140d8b9360803b7b", x"a4fa00b3c0ea6a74", x"62e1ae6c4bf879d6", x"d6ca34e2596dba29", x"0effadaa5193b75a", x"0442b5d6b03bf3e4", x"94b74ba7754b499a", x"218e5953cf7e32f7");
            when 18742132 => data <= (x"d8d5857244f8c595", x"c3e8c7f259d52b88", x"0c7e6e5c77f90c7f", x"56195847014f1699", x"caa687881b57f7a7", x"b19c98c8d4428493", x"9b60a9109714869f", x"59400918a4a7b719");
            when 31933320 => data <= (x"b0d59cded71eb955", x"466f0a636dd52f03", x"70da0b82499407b1", x"b4aaf39feef4989d", x"a9b75edfd328e496", x"73831c1088872a5d", x"651cdaddad4cdfab", x"2ed8d9e4ae824393");
            when 19003804 => data <= (x"4559abc607e9528d", x"8c8135864c28538a", x"a6d3d6cd1d4e97cb", x"354d9fd7d9202d0c", x"81d4045e97d29541", x"86732462d2c136fc", x"14264b5f3ea01639", x"3747c0d6462dd20b");
            when 6946858 => data <= (x"eb6550f2c30d7088", x"1dda7498fbd9758e", x"38e4f2d306450f68", x"11a81962dc14247d", x"d97c1490812e2fd4", x"712e6edbc5509fcb", x"1c93ac8598c2ec89", x"1621e6c30cf1e62c");
            when 18025939 => data <= (x"e63475ee3dadfdbe", x"6a351735344ed34e", x"588aec31c4a76cb2", x"ca2c079309fecf4c", x"7d33ba599bc8373d", x"d9ec101efea7b8ad", x"6d351dff8792b86b", x"20ae5ff7e2f8232c");
            when 14038282 => data <= (x"95a195a2aac06526", x"8cac11e4122d6cad", x"bc8ecbd0cb3a9bd1", x"94426fa78785e382", x"7c55445310b206fb", x"767ac8c9c3957663", x"71d0665cefb08642", x"e91fc7f0ffe9c88c");
            when 20340855 => data <= (x"0262949b32b6f0ec", x"c59754d83dede9fa", x"1c06fb1500d65fb6", x"c0edc18163080c96", x"2cc9dd59a3be56c8", x"01705bb37e2321a8", x"923ec5b7cee09657", x"bc57321e6f402b2b");
            when 6224812 => data <= (x"6c6dbcd44cd2dcd5", x"d1deff7087fef7a1", x"bc7952875c231c54", x"a2ad18928785bb98", x"dde0ac05a13cde42", x"6f7023070a60bb07", x"99e19ae895a9610e", x"ce33ca8d39ca5d4a");
            when 29924849 => data <= (x"4f208037b9f83d4a", x"7999de5e19cc586d", x"5865e4c814d8cfe7", x"e725fdd34e8a68c5", x"42eb6c44d2e4c8ee", x"ee96bf646d3f129d", x"49a0ef86e4a5fcae", x"afd073cefdb9b4c4");
            when 8266547 => data <= (x"0d9aa262bc3fddba", x"4586839d049578a2", x"73184c0cdb23f9c3", x"a073c1efded8016f", x"04ce7a015cb0f13f", x"d97ae33320e07117", x"a2716ea4cb5d939c", x"4d9ceaca55c685e2");
            when 22648596 => data <= (x"4e576b0d09b4d22b", x"aad2bc2cc2539f71", x"5ce1ebc332bc5e58", x"d4673ac8eb19e9f4", x"3374dea5b0855182", x"a11d8a4d70b2c913", x"0409295692b94dbf", x"2719368f8c17821a");
            when 26294244 => data <= (x"620f584c2542ebe6", x"40f4eb829008cbd4", x"874533de54def1c0", x"88eba9d8b815e7dc", x"a11ca2a158765f2f", x"d09e31b2d14dbe6e", x"89ebd021107e696f", x"5a9ca50eb5a82ad8");
            when 17676992 => data <= (x"5c253c722e53faea", x"381ab344a87ddb93", x"80ad79e6c08e5428", x"4007fc4f662b8ea3", x"e2c21ec7495174a9", x"88f3face7edc2c61", x"613ed45856760594", x"5f4308de6af87b66");
            when 23496374 => data <= (x"4a113586657d18da", x"1b647966fea6df5b", x"8febc5a194b44193", x"5aadaea49cf395ff", x"d6a10649952a99ce", x"a60f447bdbc07d74", x"347b482d0bf8d53f", x"782a92889188e98b");
            when 7990466 => data <= (x"68e66c97805762fc", x"feada6114e1bff21", x"0e505a8b7504129a", x"2a023a923ccf57e2", x"6cf759fd0b511073", x"50c84b98ebe9a0ef", x"8cd96a077364642f", x"9fef204225ad1c79");
            when 23841468 => data <= (x"e630857484a8e4e0", x"eb74fe603cda1108", x"ec01c749cc4182f2", x"2d7938e3a7796d37", x"fbe4997dda37da1d", x"c47e6e4c5c48278b", x"b10b988bce4a2a14", x"c72b63df77c3f5fe");
            when 10699468 => data <= (x"266e69ffd231c750", x"db6c7fc289d6eee0", x"f74ea1e4f97a7e58", x"7ac6d60b92e4116e", x"a4cc8518cc837b6f", x"6317aab621e7eb69", x"a1c5d8389a77273f", x"bc9d17504473a3e1");
            when 13402084 => data <= (x"fa602b68d3421f80", x"9ef053805a55039b", x"96e7c62cd8bdde32", x"dd296789c26a161e", x"d4180747f1491e5c", x"abc57aa0e440d7cb", x"29993fb146bfb32b", x"18448dcda4238d7f");
            when 3718285 => data <= (x"29c34400dad90b72", x"3f6eddb2f34ee335", x"1491160fee8b7995", x"ee248606d2856eb7", x"dc00973846a38693", x"276801f1b1d7a268", x"7e519b9bfada86d8", x"7ed1aefe01e51129");
            when 16030365 => data <= (x"76c26aaf5a5c0c94", x"5886896cfab75a60", x"68cfd75a3dfd904a", x"65802c49cd9ea98b", x"889dc304e82e5e7e", x"2b5c5a074117ba05", x"b10881588909d8a1", x"c9e8506f55029d0b");
            when 33890236 => data <= (x"051beee40e38a1bb", x"e7e53fb93f9f3702", x"043bbfc401bea9df", x"256c71c8da7af504", x"8d9aed420fbc9182", x"aad2a27a2671b448", x"df3b54041d5d7350", x"8ed246c904da5eab");
            when 20290277 => data <= (x"0034773377a206fa", x"8e2038fc157a16c1", x"3cdf40ed6db80622", x"276157a7bca02665", x"6e7e4bedad39a85f", x"08dc3bdbde4ddfaa", x"5dc79fe838629c64", x"1be02fad120ff943");
            when 31086640 => data <= (x"c0fd4669342f8b06", x"e0a72f67501a2c8c", x"fa346815967e2f87", x"043d721530594e1e", x"08db74e173663f9a", x"7affe359eb45afc9", x"0a8c9889b5476cdf", x"41ea46e7858ca150");
            when 32436034 => data <= (x"352b3340ce5a633a", x"e91dd3b9762a6d7e", x"ce70007d322751d0", x"e5f978d0829bef8e", x"ae0c5c70024d1055", x"1d105e6c377c631d", x"660f35d671025cee", x"a2eec220101115ce");
            when 19051138 => data <= (x"f765f6d2e0df57fa", x"9ce3d9ea6966b2e4", x"8139aaf789f6ea70", x"eaa6e1be3d96253a", x"a0d8552242266cea", x"35944bacb23c7057", x"1f7747b6686daa4b", x"631c6d7d8d69e259");
            when 27162483 => data <= (x"9dcea7165863168d", x"65150ecfff7f5e22", x"42f3a1f8a6c6f8bb", x"b6e91858a7ac173e", x"8525b55b06437abe", x"4ca286825e5b6220", x"1a3163be2c818a84", x"9611d3179fcf3e0e");
            when 17329013 => data <= (x"d80cdf6e1ebc2019", x"d91c8f61aa59af7c", x"4f22d54c209f0d0f", x"e104f1c490f6135a", x"ea988b34fe41e17f", x"03950fe1fd725cfe", x"bcf65ed8021e88b7", x"3c068713a1ca4d42");
            when 32752396 => data <= (x"0add576852b6e90f", x"e9e0c171b49e4cfd", x"e5d5cdd8ca6baef6", x"102fe1a5dc6cfab5", x"9ac58057d7c70620", x"99057410ab5e6806", x"e2d3285ed9655e9a", x"4bd82f3c7147d017");
            when 25981544 => data <= (x"ebfac1ed44d0848d", x"f8b441b7ed20eca4", x"be90aba648bf3a3c", x"9c3e699bb6b5dd85", x"be056e3419b0bae4", x"20ae254a40a0b564", x"e50a3811b5eba789", x"eb3f6e99be64eaef");
            when 1093898 => data <= (x"65231224ca020754", x"b7241147da6b1af3", x"4b3c6637a2a1c486", x"8e8f876ddbca5227", x"9554b47956e968f8", x"ec255d08f6233639", x"ceea3a69e1000277", x"744acb179b94f185");
            when 20098527 => data <= (x"86b2b27959024e09", x"b60499484e55ecaf", x"76f319262ad5ffbf", x"6be21d65b7c9e3c4", x"0ea6930c80fbabf8", x"cf66a28f52df4d1f", x"eaa7d52c35e34a3f", x"d52d82012b9a3a94");
            when 1665092 => data <= (x"2775bcb1cab087e1", x"3fa57e52217b24f9", x"9c069961437e52b9", x"8eb6ff11cb2add52", x"59401e9c38debacc", x"2fa45964079e8ed8", x"08434ebb1f8d6df0", x"1e8dd60e587614a4");
            when 18099957 => data <= (x"fabdcd062c24b8e8", x"5acb1cbf45068607", x"703c1da8c4ecfb07", x"7595cde333724c66", x"1962baada0fc125e", x"1d5d3021e970b5e6", x"8f0570216f410cc8", x"e96000d081d195f7");
            when 7848663 => data <= (x"302b3fdb5f268dab", x"05e6f98f5ad50da9", x"04908c70d5418d8e", x"39ffcd92e064e1e4", x"0361260dcbe12747", x"90476164687f4f4e", x"5478cc207b76bea5", x"3e81f0a6666065ca");
            when 27230961 => data <= (x"e99b065d7bdee825", x"ba3d69bb126b1b77", x"65c6e6c5ec942d3a", x"7139164ff58f9dc4", x"42a94f66fe033286", x"6a7c82041a29ea81", x"041a7bcdb36213fe", x"2064ca5f61d49df7");
            when 28388916 => data <= (x"0d088038420c5efa", x"e3dc9e7aa56c468b", x"d57e15356ae4660b", x"da303a3aa785d426", x"460ae58724cbd445", x"9e363ce54f454120", x"0d13618032e34b74", x"116c67b503922d89");
            when 5757303 => data <= (x"4ba6ccffb4c1a2cf", x"8f92e2a34a01eb1f", x"5506c838cafd77d8", x"ba7716a736e254ef", x"c402f7f63df299dc", x"b64d8cd2dc5c3cd8", x"3514e2d705a4040e", x"f479f971bf740df3");
            when 25268829 => data <= (x"d90aeb76579ec326", x"b9a1d9f880a56a6f", x"1dee5fca56b59b26", x"d115d5f008eb045c", x"35c04f3acabef047", x"0725f3517ba17dce", x"968c31a49e247479", x"ea0797c5f15f03f1");
            when 32806213 => data <= (x"d1da6a13f685cded", x"e9633e242500a2da", x"afbad752e753676f", x"92367d0944595201", x"9c104c4335dc1524", x"dc9948ad6d617a8c", x"4941ae4cff37d1c2", x"367f79f1401e0e45");
            when 26330815 => data <= (x"780ee1f71afb967e", x"26cd050ca528c6ec", x"616ded1ed1348564", x"bc0654248038e1ce", x"f4866435e08356b8", x"1c226b2438c99ee4", x"25c905a8bbb5b2d8", x"b49fb2cbf7cdc5ca");
            when 19652640 => data <= (x"c0bf6715b5a0808a", x"40f05c716e537392", x"b1f40974e1f93990", x"f103a484e36e893a", x"3ef0cb8fdb3f08cd", x"3839ea2c549fbf8c", x"74b28a3e20dd0caa", x"8bba18784a0163a1");
            when 24246031 => data <= (x"5be2f5cd58bf7be5", x"679a0714d3e8f852", x"ead1f65df169f81c", x"cdd2aa2e2ad84de5", x"3fd007312fdb51c2", x"683e6578426c88c2", x"4364fc9ee7ee7c65", x"657e33264ee02f2a");
            when 22782020 => data <= (x"93f4a8f484ea1719", x"83f5a4331836466c", x"c4d6ca9c9b500d95", x"da7a9d1b47c06ad4", x"48832677daa573bd", x"f76a6fd21a2cddb9", x"31399690c4b14193", x"c16a6fdd8bea2c1a");
            when 9000434 => data <= (x"f9d123a23909cdc8", x"8927ad569bcbd587", x"a1c13582962bb7c8", x"bca4bff729c01637", x"475559972aeda970", x"8a54cf06502f48f0", x"a021346173be6993", x"0640a7174cf831b4");
            when 12789955 => data <= (x"4403e9be8d51c453", x"97aa69727f03b59c", x"dc7162d9c93b3350", x"c69d9b72ac2eff11", x"7d7561db5b7a1124", x"b9412d6082546a78", x"ea0e3cafb34ad56e", x"120dd7ac5775483d");
            when 19925772 => data <= (x"18dceb85e0b10115", x"b84cce8a8bbc6aa8", x"b952282429eca30c", x"80572d5ed025ccd4", x"ddb784882560e8f0", x"e506274ad137bbb8", x"d8a9a416798ef0c4", x"306fbd67fc64fa03");
            when 7246179 => data <= (x"efd40ae1f0e2b099", x"82d85cde1a6e6a54", x"6ce233b8a3c8d738", x"79a169d314e84815", x"d921fd3ab06580dc", x"423e328e07582126", x"7bd262bb8fcd2154", x"639e6884f5e98857");
            when 22651984 => data <= (x"f7ed33b8883cf767", x"3586d2d75b100891", x"d00c83624781b048", x"9c0716d7fa94e3d5", x"766909a2b282533f", x"c76cd711820c2a2f", x"ca75919dd639bee2", x"ff3706eda5b2ba48");
            when 33343930 => data <= (x"5b1cf562d1dcb873", x"02f39d1c6ea6414c", x"2a4ca008b203d322", x"e199a496593cc650", x"34479a8800d93d3e", x"6337d6bead539bf7", x"54ac3f23de95ff4b", x"88d8f8135093f4ab");
            when 29074455 => data <= (x"1c6fa63f515be2d0", x"c15574b5e37f6668", x"b58203f8b181adf3", x"b0702b78e8f467d0", x"dc961c8d86f1c735", x"0cb3346cdbb3e26b", x"2172f0d9877353bf", x"38f6bf24717ce985");
            when 15102849 => data <= (x"f07d9d53a8c041cf", x"6ed4d7ac41ca987c", x"0260f68c644fa458", x"635d0e75119d7d9e", x"b28704d6d628ba49", x"0e85eddddd494dc8", x"76fdbb9a2f5db0f8", x"0f959abfe8dc9723");
            when 2257139 => data <= (x"8e611e7209c7a9f7", x"3d816f9b232fe078", x"54319777341653e8", x"7c49816da303d19f", x"0fb152104c636fa7", x"40531df8408faeb9", x"6b834542b4eefa82", x"b2ebf7949d80b121");
            when 22026780 => data <= (x"c04b83dd598e8ac2", x"fb9dddbfb11443d6", x"ce7a4b10680bfa31", x"515f7b29ba13a80d", x"853b487e2297ef0e", x"f343dd539999d6ab", x"5d6857ef5ca66c2b", x"8c45a13e83bda460");
            when 24481829 => data <= (x"6685bf599af25623", x"af151a33cdcfac58", x"d723fe97736902d3", x"a38d42fee6692334", x"7d4203031b997090", x"1b4ee6175d0e5ab7", x"289b53f3711b0777", x"9c54ca3e652e1c62");
            when 18631267 => data <= (x"a52cba2283963b66", x"0015be3992beb4b2", x"0fabcaf6f8e88c3d", x"660f3dfd7eca9389", x"8c7dd2f503ac873d", x"edb067db5a721139", x"08c71dfa7fdff5dc", x"8472785aac6d74bb");
            when 2575779 => data <= (x"0bcb4cba81da94ae", x"1d9eb70db5f07b14", x"c90a5d792fa65a93", x"d04e6b3f31eafec7", x"ffb0c5164411b08e", x"38896549b1bcb734", x"e51cd59dc443d1b7", x"d3bfb3ccee21ad0b");
            when 19852001 => data <= (x"67d36d36fc8e26d5", x"c51939aceff9617e", x"ce6e1833b86ebc39", x"0194da9f1339668c", x"ae07568e7b1538df", x"cefa7168c2cf5de8", x"25106cc595209e85", x"04436cdbe95a4b4d");
            when 5696606 => data <= (x"74729ac86562b9b8", x"a2fbc1f43044a496", x"a4d1308a65b75b01", x"656fd671ab0cee5c", x"183feec3b83dd17d", x"5abc8ab49abd2947", x"b36d66fb82beff77", x"517e915dda982046");
            when 28550651 => data <= (x"430b109c3b2cecb0", x"f95eb06dc545662d", x"5dd293b9594689bc", x"c654f44bc01d3267", x"bac62d27d289c680", x"8a5d4774e3f212cd", x"5e62d258bb701679", x"4a2eede51231cab3");
            when 2220761 => data <= (x"78e27820fd89d1f7", x"75eec4053e221bbb", x"792550ac05c4a923", x"7cfb87dc36590cb3", x"3e5343a4d438338a", x"3a4b2924fbb521ec", x"f2a46197598bb7fd", x"5898f75826d05fad");
            when 1506560 => data <= (x"d19db87203348b20", x"8b328dff09e60812", x"8030b282779e1116", x"affb6a833947a565", x"01844cf8b9fbea64", x"d4de29adcdd44ea2", x"c0b373991dd72d9c", x"e8ce4f0dbc600f49");
            when 1377505 => data <= (x"8de15359e1721156", x"83c1bfe0289ca9f4", x"a587a1722044a968", x"d583b5b7c0490d98", x"2f4bea0c5aeb5d01", x"b802e1482a98d744", x"8d11d99691360b60", x"2c8c98f54e59fcb0");
            when 12852845 => data <= (x"af2b35dca77d86b4", x"71a09a9971bb2ce2", x"d2e3791034639023", x"9115c8555f35f0e0", x"23bd5de5d150baaf", x"0d560696c8d27ddd", x"ff97c525131bdd54", x"b5966e8c8bedc559");
            when 14166438 => data <= (x"40c228cc54971738", x"90c79290e8197e06", x"f1be8aaa13ba5a84", x"171d5029aa419393", x"b4fe5a17b18724db", x"a671a248de65b250", x"6c385d9d4a895f84", x"4886a23580d861d1");
            when 27969268 => data <= (x"fbae1d61fb51d5c5", x"9bb7fe758b632e31", x"718328fcfc96b746", x"ed70d11184e429ae", x"79f0003832066a3d", x"b959afb86bcad15d", x"c0a263b40337e5ab", x"b639c7bb57e48f4d");
            when 13905310 => data <= (x"47231120426afd27", x"d912ce9a38080036", x"d6461cd8818afec4", x"394b3edcfaea47c3", x"0c49c6a45ba9f1f3", x"61b6b23084131438", x"ba4aeb3218f310aa", x"b1586a9ed5751519");
            when 28526328 => data <= (x"91c155855be31569", x"70de8b8d1f846146", x"2256a0f50ed22570", x"a9dcabb9baaf8614", x"15bd12f54087cc5b", x"c7648387fdb82976", x"319c1b6d5cd1eb3a", x"22313ece8d2051ac");
            when 26378294 => data <= (x"59ebab293983c91e", x"dea408560059d370", x"0a2c662d70d57ece", x"5b7cb2de53f3c667", x"3d2eed2e73d18be1", x"d7e47857a0509754", x"0b6034bf7036b562", x"a6a78e472bdb59e7");
            when 19828013 => data <= (x"8af9cf9d573c7d02", x"a0574dc4fa0c486f", x"4a6f9543d89de2ed", x"993ac793d5784127", x"daf4893a5143a2b4", x"cff3e4577e3ae9d7", x"9415ff93e516e16f", x"c44ab9d90387a3ce");
            when 20359583 => data <= (x"44ed9509c71cc296", x"88974e7a7eb7bf45", x"4663fce7262932a0", x"74cdc438323a208c", x"00847c4481e6f7b4", x"95699d21aaf7fbdc", x"9c9da0da32e756d7", x"e6e2f4136a35fe27");
            when 33402894 => data <= (x"120a7b51c8cb1bbb", x"b7f9e2c05eee3a14", x"958ceac6cbb29c6b", x"d108969efe4b7fcc", x"39110ae82ee54456", x"d05d96c5f6222f76", x"1dc872f5415be0bd", x"04e74a37d1069316");
            when 18656002 => data <= (x"589cd4136c44a4f7", x"1775b2c98b044e2f", x"7e2998d67822c546", x"5180242edd546747", x"00f3e72c01ff58a3", x"55ec7fd15acbb7ba", x"035560dd5d16f2ea", x"1e68e0101526be7a");
            when 2127954 => data <= (x"4051939f1c7a3b82", x"e6fa22f91cfbfb3f", x"ed635b852d231484", x"ffb5133c150d6539", x"792b76c06cb18353", x"592faecec53735f0", x"7c0368527cf109ed", x"095d098bcb438979");
            when 4639284 => data <= (x"8c118ee3794b98af", x"0e38459c3243cffb", x"5465349cb7178a7c", x"64ba2b6c5e9c8049", x"0ba69da3ad627e22", x"d22766825905bdb9", x"f122aa3612f40ac1", x"093063b834a15f2d");
            when 5131536 => data <= (x"4f0093b90783c9e4", x"e244a417beb7a1b1", x"0214f34c746e5746", x"94e946c48101973a", x"b745eccf5aa07a53", x"f2aebf9282814fec", x"cd95e62d99e89c11", x"fd952426bfaba2d7");
            when 21559443 => data <= (x"8725828c402bf526", x"5ef956e5ef7d2b3d", x"412045e1cc23f33c", x"200d96beaecbbd6b", x"521b817d04c15f39", x"63caa7143ed13ddc", x"96e3ebe76cf2641d", x"ec7b95f1aa55c94f");
            when 15622362 => data <= (x"60a21525c0c5d2f1", x"d0eb8acc190bd84b", x"4d0d568ad669b21d", x"1956c63c89db93d1", x"0b90bb6c40539d23", x"3b008818cf4cddfd", x"6e7230ca1ffd9fcb", x"008cb87940af4ba2");
            when 29445706 => data <= (x"825f86b2d7239431", x"cb5aa2c93cf1acbd", x"586fcb33a59ef60d", x"109693535f4d8535", x"4b0baff777ae44da", x"a759b4dee4731e9a", x"9cd09ec0739383f2", x"89445ee8f49f08aa");
            when 17279890 => data <= (x"9d426b3f7666cd63", x"ed18ff79b92c7d9d", x"83335a5c0d266248", x"e0f40e097c207a16", x"7cb0458557d687ee", x"354c4e617b7fea51", x"1b096e34a67360b3", x"c97ceaec9b657cad");
            when 14035701 => data <= (x"e79aeecebc834a39", x"79a571da13e2abaf", x"d8d9943c35125285", x"382c395c548b24ed", x"c6fd4743da34b32e", x"7873168114262d24", x"2279224b61d813f0", x"c2a9bd562081b4af");
            when 32241735 => data <= (x"045449c14de08b60", x"34080de9553e9463", x"a393034b1c0dfb83", x"a474c6ea596ea471", x"94bd33dae7d4d2e0", x"d72ea05ceb8ea67e", x"504ed4fb099336e5", x"c6fe58bdf72599e7");
            when 5604280 => data <= (x"08bd2589bcf0e123", x"bf51780f079d068e", x"809e6505f49a2502", x"c490323b0af6c375", x"47901630f375e7fe", x"ff810e4d4d9a2d1d", x"66acb6361a44d513", x"1a2c324974cdb1d9");
            when 28834450 => data <= (x"4fbcfdec170ec21b", x"32a93cdc692aaf4c", x"498edfee901933d8", x"f678d432520c316d", x"4e2ea4ec1e999ea1", x"7b01d42e5c692206", x"78df604354964b5d", x"a434e7726ce70353");
            when 2034554 => data <= (x"89a7ac26329bae91", x"3fce5541acfd9724", x"67b7bb7d9796782e", x"71bb281338129dc3", x"bb6667335c62bd4c", x"3cd73a341fb86d3c", x"ff22d0059404f56b", x"a85d6eafa7da6c7d");
            when 10300748 => data <= (x"32ad2c5b76743b7b", x"ff7b924c9910311f", x"d438ab74deb4e784", x"a76c73f141a6c424", x"8da9df7c8e4f43d7", x"5536fc144ef831ba", x"3dfe2df3c107ad59", x"2341563e8b0f0a83");
            when 25869658 => data <= (x"317d0ca843fec5da", x"cb2bac08a94a90f8", x"59459e61eef42fc3", x"ba4cf0b92d12247f", x"73fcb7514fdfdc64", x"ccd78feee2603e62", x"b522e6e62f2c980c", x"cf6dca035cef168e");
            when 13019413 => data <= (x"28d34525a402f95d", x"4cdc9787df6ce0b5", x"8d0f3672464ee461", x"cdeed1c1670915c7", x"8351f174c2a201e1", x"93e0432cd5a01b93", x"b0579ae51abad9b8", x"d4caf1880b1dccde");
            when 15154026 => data <= (x"3d15ee48ff719d49", x"87ed6ca97960d313", x"b39e4b6c764b3ba3", x"f083a6e0380daedd", x"4c251667ba2669a5", x"cb7bf7e70b2bc2ab", x"bde5bd06d6e3bde3", x"c3c3f1b2c5ff5d95");
            when 16207209 => data <= (x"33cece05349fb666", x"6bb9fcb8a98c4bff", x"10ed19454e4b21ea", x"061026e81a046af5", x"9bd64d3949e5b3b2", x"0639bea25cb48670", x"f9e06d4b2aeb7c87", x"ac686ee9f7abde3c");
            when 33876481 => data <= (x"1e9c92bbbc83071d", x"6e1fa77e970a5d16", x"bae60991d354d5e3", x"402fd9981926d4ef", x"7ab4fb203c605810", x"dbb89829eb92ae08", x"ef37f54bc515e808", x"9d1846100bea99ff");
            when 9137442 => data <= (x"d394d975a40ed12d", x"8247dfb1ec23e46e", x"10caa078c247664c", x"e7e70629c137b7d3", x"b47b9e24402fa541", x"735b99e5134fa2cf", x"274c04ac92e26c2b", x"12217409d1ddd2be");
            when 3760146 => data <= (x"b49906becce9d8b4", x"6e8b23f540971e73", x"a4960adc8d4561e4", x"f94832cb6a5efb69", x"685dd254d18cff82", x"63303452a35a53f0", x"b2df23c4e2e21c98", x"6d59ed79b327fe1d");
            when 19106581 => data <= (x"42676dc6a334b7df", x"ea0f6401b5042767", x"15f952af7c3712bb", x"b634c58bec4b4edc", x"e71fe9ddeb173bfb", x"0d95cf21378a113d", x"eaae9467761aca28", x"168c02ef46f3114c");
            when 13351660 => data <= (x"fa23ab68e86a3a05", x"de9b567db9d924fc", x"1afedd7d67dc6ed7", x"2d8162c3cc2b9ef4", x"35173e09681d3b76", x"94bd7848d0f6450d", x"0a766ce7b625fef4", x"b56f0e87ebf8e3fe");
            when 22676785 => data <= (x"ec02ee41e1e10f75", x"a4710f744a27a12d", x"6fd03f72ffbc8874", x"6d968de54c87b4b8", x"4da65188d06104eb", x"edd76b01a24ac396", x"4dbd07c73d18131e", x"64e1dbf44335f3aa");
            when 30951580 => data <= (x"85345a299b9db438", x"67f76be1bd46be69", x"8d126586a8e347d6", x"5291dbab5b561916", x"bd64f48fd5e22f3f", x"916c5b41171fa794", x"de3753b642089794", x"d3842ff71248c342");
            when 21938331 => data <= (x"4e349a8e086670f8", x"878586f4b5262e75", x"80b56ee091532056", x"cc21b87003d9fdf1", x"798510528fefe105", x"e68174b7e8dbe572", x"2a1c47a15e15d3f7", x"8bab71254830489a");
            when 33060685 => data <= (x"63d3342fc3ba1e7a", x"96ac8646ea93c38c", x"b99982f0c0a8b48e", x"6ca2d7557f7e293d", x"297152c4137bafb7", x"c2aab6457fb91bea", x"b5ce5168cd4171e3", x"8c919f50b4b7ea0e");
            when 28866382 => data <= (x"f6a6bb1910c91a63", x"78196625297497be", x"e450123105759a31", x"97fc4babe5e9598f", x"c3922d7be570735f", x"baea93bfe9f49f40", x"a4b7e4218a0f9314", x"a9d3c7efb7dde697");
            when 12453949 => data <= (x"d2aee814d26b6b81", x"b290a0fa57b0834d", x"bfb8484810e4c9bb", x"4fed1cbbd40774b9", x"ae872af0d83e010d", x"48aeda237c3d2d51", x"f30cefa031d77c9c", x"d28bb8cbc8738ee1");
            when 20026140 => data <= (x"2f72842890328e7e", x"7616126826c44777", x"83e08e8954abe3e3", x"39a7714f3ad24620", x"56c920ff632404cc", x"1020028e69eb6c62", x"ab49a4168435a596", x"f9c16d000cef2b43");
            when 14296131 => data <= (x"5428754618c8a11a", x"881ad67a72069553", x"cdb6f19c7597992f", x"dd558613cdbca093", x"4676988e01fe7ed1", x"8660ddcf323d3aea", x"35f12b34dd67b714", x"7ff51b8405c0260f");
            when 26422261 => data <= (x"afceb4d069222634", x"15c4800387b94715", x"187311e6dcaa0843", x"b44d1cb09f0e4cf1", x"1cc8178ec6baf632", x"efee564a53b08e59", x"b479b51a4d3deab9", x"793923878d21ef4d");
            when 23147593 => data <= (x"1f25193e381fdf5a", x"645eab35bc3b345a", x"21e17eb2dc41b025", x"3dbd8ee1d3b3e178", x"3cc8e390e2092e98", x"5725a887341e4cc1", x"6b7dd157a4280936", x"f1dcab4d020cd85a");
            when 27948221 => data <= (x"13ebb7b2139dc514", x"254b773eb475ef50", x"8f3d4db819241829", x"8580cf2c7504c19f", x"b56fc58f2cd79475", x"460140ec562ca661", x"de2c0f6f1f7e190e", x"2298e827ae025478");
            when 32222166 => data <= (x"f168fc9d3f8f24bd", x"8a0564cca5043636", x"4264dbbf58e3178f", x"803df5de4617c9b5", x"dd778b86caa84f0d", x"cd6af68a0e7892cf", x"d724eed88321b4a3", x"fb7b01a33e8ba3c8");
            when 27165554 => data <= (x"1e89e2cf4c41ace2", x"e48e01318be6b34d", x"bf4571879fa06621", x"101941e94450208d", x"774f1c5f376b3325", x"252d41dd9859ef63", x"cad18b396a4232f6", x"eb332fb42fbe05b6");
            when 3407701 => data <= (x"b74b6d8d19a73b9d", x"9172219f2bcf5bdd", x"94c091953819b1be", x"fbab08cacbdc5668", x"3f5f76b2f9d7e19f", x"90ab60ea2e2082a3", x"b8efa0b9e32d5569", x"9df840e189bd4cd6");
            when 32607930 => data <= (x"d5379caeaf79ddf8", x"60f093a4745e88b4", x"ab417684733586d6", x"99cc9b492ad9fd9b", x"7a042aa78f5e53b1", x"e7deb43637451188", x"d273391f48339155", x"aeba124821c48f00");
            when 24486391 => data <= (x"8d68885df14fb9c6", x"0a4430f1ce3a31c5", x"17d4e135d2e7d40d", x"bcc640d48bf441e2", x"b59b0fa4fdd74718", x"e8d5f1441398be7c", x"5fb75b0dfd0b51fa", x"dffb6d9c404568d8");
            when 6091643 => data <= (x"4c48d562c230cb8d", x"463369dcefb3d9bb", x"2b2cef200873b6f9", x"5254b97160285c76", x"957563046c459f42", x"8fd85fd6c364433d", x"e28b1c53e3809203", x"2ec70a416b77fbaf");
            when 28491881 => data <= (x"a6604629f69ea664", x"5ed1cab10c3f3a3e", x"9040cc525a80cf34", x"a87704e5ef7cb3d5", x"1b6f1040b8080bba", x"e20f82ff40e5f5f6", x"2374338af2a9d014", x"a413222077ce3b7a");
            when 23249109 => data <= (x"0d2c321ff7c83074", x"6c565bf95dadc730", x"4e012796b6bcf6b7", x"8aab0da1aa39cb30", x"e807b5c9a493f129", x"29fd9ecdf3e2703b", x"9e170dfb583aa6d0", x"dc3bf61ccdcaa66e");
            when 22359800 => data <= (x"2feb6164f9e0709c", x"5e45c231f480abe5", x"5c9b6df2567989e0", x"50ef1ed51e916ae5", x"04a5ea260389a506", x"c78337bb1442ca53", x"dd7e60388cf2e64c", x"efa1ba3360fab4b6");
            when 427207 => data <= (x"43ba8ed3e7918b59", x"b7f1437b10f31a35", x"5300399d8f749176", x"a96b7a58b9fe9727", x"b966eaea895ef152", x"6c3d78f11c5fcd46", x"d8125f608379e000", x"3c9858b91acf7c79");
            when 24646164 => data <= (x"7c64bf78e549238e", x"dffed8bd7c1e8dfc", x"1e1ccd742a854cbd", x"3b4bb46f6519b71a", x"6dd8dbaeca6e29c8", x"74671ae0986a12fa", x"60ad6726fbc20b69", x"baf95c27a341761e");
            when 30471723 => data <= (x"1c230032c361e511", x"a1c5d11407f6b9c7", x"96d0d6817a25993a", x"104d8d1b2e9743d7", x"19a08a7f4d2c0fb3", x"5f2fc5ec712d8a61", x"8b3c10acfc460a91", x"1bc88bc59a3c1fe7");
            when 33168933 => data <= (x"d247a2bcff5f0449", x"05a232aca112249d", x"97f9ecf30f46d14b", x"a93da6ec0b087191", x"827179b466a88780", x"aecc61e8dc0afe27", x"d28d9479bf28d9ce", x"1616d70b86cde716");
            when 4213374 => data <= (x"fe09da17b7099bf9", x"fe924244f530b359", x"d2c5710bbaf3d1ef", x"2b9766328e2bfde4", x"5568e38619d9511f", x"e6418734af3e97de", x"d9c17c6513b302f7", x"6b1af38f5d7354ce");
            when 6900180 => data <= (x"2d5adfa75ea145f0", x"7ccc02df37a1ca5d", x"2fe1b884f0a9927e", x"5c225851fb1c9341", x"837f6138067802e4", x"90c26f0256e1f3b6", x"f544c50b437e7fde", x"174c92f532ad668f");
            when 2804262 => data <= (x"f48fcf2dbcb85f4c", x"26f91ce10d765d04", x"43fb7b0682f511fa", x"c49973bbb49515b5", x"e5416d66169c8e2c", x"828b570321e31b47", x"a27a8a6abf77482e", x"0ff7602c517e7b39");
            when 10461586 => data <= (x"1701d841bcfded6c", x"87342c3f6058315b", x"d5d61058708f982b", x"fdf395df6685347c", x"cd435e1e7dd9a2ea", x"8a95b2753ad618d5", x"e6543ef4fc5bd74f", x"c7cb1d3f1d009fa5");
            when 3683254 => data <= (x"387eac4f4331b47f", x"30fe35031e75bbd4", x"3c7795c69e88edf9", x"1861acf5958e2b5c", x"2a690fe46d5ef4e8", x"24a332d8056625a5", x"5b2eb93cd20f7a28", x"dad305da1cac520d");
            when 8210489 => data <= (x"1a82b8b0e365d859", x"f9608cf78862be37", x"4f9d6ed7cd218420", x"069819c45fb0a055", x"4faad8a5de548973", x"c75e0ecf01fc23ef", x"da7ed96adea98144", x"afac162fcd83f74b");
            when 32199241 => data <= (x"9f629839520fd388", x"e499e99776351c9f", x"8aab4d7c351ea063", x"cd04c95ea7ac0363", x"f58c2908b4884760", x"eb79b5d8c1c09f9e", x"1f95879d8c52ca7e", x"e92fee52140d5762");
            when 3686571 => data <= (x"ee4bf33a026a08e8", x"cbd35ace0f6de1cb", x"effe95e708977e25", x"d2d16f569d7e353c", x"7d080aaee7a1f5a6", x"0d8b485fb67787f3", x"2886e2cd67ef80f3", x"a891603d67fe7f6d");
            when 21374191 => data <= (x"f8f7313834db9e47", x"7cb1238f0b6dc355", x"d2a9b617521c5ab6", x"d80dd3e3dbe86cf0", x"b7af185e25fa2423", x"012221316b868551", x"5881597ad94d7a3f", x"ef28f99626f9d6d7");
            when 856277 => data <= (x"c9b6b670a2fe77d9", x"a7990efd85eef836", x"fd1fe45c0fff7ede", x"9bc850554238f1e0", x"9c157f688ba2a835", x"40eab52726d40912", x"4bb7a777125b586a", x"4e903876b5fe8bd2");
            when 15921660 => data <= (x"31bad780471e9a37", x"47fadd0b64d1a558", x"d88d6ad9cb0b9299", x"33be694ee22096a8", x"f5addc0ad11ea71d", x"0fada1f7ec6ee91a", x"b371f14409a107e8", x"cdb06758c8134f7e");
            when 7738914 => data <= (x"ff6171ce2a9bf7aa", x"6807fe3974df44c6", x"3d2e4597b84c5a9a", x"708cba1304e065ee", x"dd12c7b8e77d549c", x"ff94961ad0357391", x"b42a7746fa44bc68", x"e27928f47da4ef5e");
            when 15796840 => data <= (x"0298cb1ff3293403", x"4e5e01c2f2b2dec9", x"0e3deda6084abb44", x"20bd106a9c2363f0", x"3b72db03a785ae23", x"4383cbd7bd8de5a6", x"825226c19c264c64", x"42860882e3d5d8d5");
            when 15885604 => data <= (x"f5b45ad0227f020e", x"2d42bcde722fbd1d", x"7149038897f2073d", x"27534e5570727bb7", x"96c6de48528f8e9f", x"6a9be64bce542e55", x"56129cc552e5f637", x"ccbb230c0325004c");
            when 14354136 => data <= (x"079fab61fd58c4f0", x"d66114377f2704ec", x"205c64c6a9dc55fc", x"4f584f910c76c32c", x"8758b7b8cdde4e78", x"d296bcfa43d3724e", x"90dec65c18710fec", x"5404957fd8f52ce7");
            when 12369314 => data <= (x"956b708149419f73", x"4d6341a4c923c023", x"19744273568b675a", x"6cd31a3f67f19004", x"e68f2a52b6d1258c", x"521e0e957d610433", x"908228325168be2f", x"93b042f8c8a9eddf");
            when 4284423 => data <= (x"a6d3ce4d1761bf21", x"0839f3707209859c", x"d40f8f54898ac69d", x"0a0145cabad5a67c", x"1ddcf49e132fa506", x"47bbf4e5ba733653", x"eeb80f8262ba3501", x"445cafebdb4c861e");
            when 18370268 => data <= (x"da3a9ccb057b370b", x"f5f0483316bdc409", x"ed18701aebe06931", x"86ecfc86ebd4026e", x"2d0c0b2e90d087a0", x"bf64f1784e4c7b97", x"ed9a5d1a8f569490", x"4e092519ee1db623");
            when 33137254 => data <= (x"a92252ae4c9c5514", x"ee20f5815cd29ddb", x"bdbf245d4094fc9b", x"95660dd1b4c55bf2", x"1bcb62873ea15088", x"cca9b5e77bb385da", x"27e002ba9c074442", x"5000f1c6597fb6a0");
            when 30565319 => data <= (x"772822935ba194c9", x"3410f4d788070ff7", x"8e38789efc3a6534", x"229ce091cdc8fd43", x"8c17defa09e3b936", x"67175faa91249aa1", x"6e0969f2f199da0e", x"18d8fce7bb1a10b8");
            when 15996422 => data <= (x"0f28a96280348d76", x"49893c9a8d1c8f82", x"c7814bbb3c7e0459", x"7ff73146292d1614", x"070f93aa0b53b4f3", x"d7bd5c628c8ccdb3", x"30a016790d8b57b9", x"565a1948242eb15a");
            when 15416222 => data <= (x"ef4bbc007ac1fe18", x"4138ac3eb6bbf150", x"b1d7d1dab0de3acb", x"2eacc7de706506aa", x"a4d9b4e96b71890e", x"3f93d2ddebf21b22", x"7ba2f9a5ebf472bb", x"525e120b88b3cd38");
            when 14524785 => data <= (x"25178ddb0f5ac0b7", x"097e6743a0b0e68f", x"212c00bc090a5a1e", x"5c1257732b1aeb3e", x"135ec206003014c0", x"35e4bd379b42b38c", x"2f246c194711b7ae", x"1fd8607b0f5b41e5");
            when 31617015 => data <= (x"0ef929cb034f2ef7", x"5d8a9fc3ebecbda9", x"10a7d6eb844f11c2", x"c4dd3e11022126d9", x"06a10bbc3c6a6c6e", x"ff2a0e6984675778", x"ce7277e93b204a2c", x"2fd39007169d75a3");
            when 6477338 => data <= (x"0830d2e3a7bc23b7", x"8d5fc1f590f19265", x"9edbf2250a9b814d", x"50786490cd51a714", x"d46df65ac78b644a", x"55cf5815980940ed", x"6201fb3728e7a81c", x"c159f970daeeabc5");
            when 13960741 => data <= (x"044d7e753029ac04", x"9ee3ff6a85926956", x"ca8e68f3b1050949", x"0807cd700e6f2cf9", x"1a4c1a19b8ab54ec", x"0bb221f74bec3a91", x"6b4c42e42214cfaa", x"c36daedc08d6f582");
            when 22006140 => data <= (x"ea816def50d3790f", x"5f872a2fdf0c3773", x"997196ecd356f5b1", x"06a7d5d4c92d6a16", x"72c23e40df8bd906", x"77124e7867b7d37e", x"8f2d0a876b708808", x"edc32e8b97e546f8");
            when 29491440 => data <= (x"9e8287628f5d270d", x"3a82c307c1828cd2", x"d055a9bd05632db1", x"34f4d575fb4cf843", x"f6c81771557d3e0d", x"e5d216300446a57c", x"407cf2cadc16b872", x"55e715fa2662fef3");
            when 21102385 => data <= (x"dc148d4009989271", x"60706c1d22f67a40", x"4a48d66eb69350a5", x"792523bbe1dccc58", x"b089d879ce46edc6", x"9c5de6b0b6301e72", x"028e6389065a013b", x"d589d6588c542892");
            when 4747923 => data <= (x"e37f00dad44d8db4", x"6a19ff9d70b71f34", x"1950175e13fe3cdb", x"5907d1bb74d4951f", x"3e9f0eb8f914ae0c", x"645fcb90b877bd9f", x"f83d6c003c63a892", x"f24f467f11527be0");
            when 5379072 => data <= (x"3991e538d9beac92", x"ff9a61c3a69e92f7", x"b762d233271cc086", x"d0d46698aa691a66", x"1edf5d99b94317c5", x"5f92a488780c6294", x"e2efbadda0419c17", x"a102fd2930f089d7");
            when 7217794 => data <= (x"63fa5245775a75b1", x"28aa49294cc457c6", x"df05a21e705e298a", x"745b45cdc18be236", x"a13791fa888239ae", x"6859892b076a32d8", x"7a9677c22bf4c5a2", x"bdedc85548b5fe1e");
            when 15044920 => data <= (x"73527e7858f7b8ea", x"5c8312e859a90c7a", x"80650f9486a4839f", x"2c31b1705c960357", x"53b1f0b6e61ea42c", x"5464f2127b6a4bf0", x"3e2b3724b559c76d", x"d78ebdb1a882fe7b");
            when 30843533 => data <= (x"fd6e731b1d8d7766", x"c51eb6440a2a6198", x"6e36cc282ec37d44", x"e836b5bcef63a014", x"c2f68a447957e39c", x"1aae117090184ec3", x"766a8c4114e10114", x"2411e4802b5d17b4");
            when 25438133 => data <= (x"1427a7b49937e330", x"bc66fb368fbddd23", x"3a1367ce97ab53b8", x"a06ef629486449a5", x"13d543bcee1ceb1d", x"e75837a8121202bf", x"0f8a1ee7f28dd28b", x"57ae0015efffea2a");
            when 2083763 => data <= (x"c2e5cfe38060c35e", x"9aa2de63d7340816", x"283aa36ff29c3c0e", x"28f0838de0c3ce7e", x"37d1f55a194c20db", x"71bae0dbc8efb6e6", x"e1b7f61e260de09b", x"1436589b04c89a76");
            when 9579138 => data <= (x"ddc59c6d69295bc7", x"4909827630d7f4cb", x"20b8a9c3f475f453", x"321a88eb90167c35", x"28f3f6bed2758ba6", x"0fbc1dd1056769f6", x"898be21dd2d2b589", x"45f94921db6780a0");
            when 33908611 => data <= (x"e5fcd6921166eaa2", x"4cca86e1dac7ccd2", x"b70303eedc1bc0d0", x"94932f250567906b", x"e4ac2d06de15a40d", x"9b3b01c9615ff4bd", x"9211b5a1efb1fb45", x"5437bf156f120494");
            when 23197761 => data <= (x"afa02be15eebabe7", x"75dd19ef98165b34", x"7efa5cb0b1218c95", x"acae5d752a9abe01", x"b1d5d763f1f9f501", x"e92fa03bda66c298", x"752187c377dd17c4", x"1993904e5f27c11f");
            when 28305007 => data <= (x"abb47bac3fcec161", x"e64982e38c246171", x"2b2bae1ad232bf00", x"166975e255d30166", x"2f5a982a84325395", x"732aacc01ed7ed16", x"3b3a75237c3f25e4", x"8a1e21c88ded5b27");
            when 8616479 => data <= (x"72596ca869a99e1f", x"a6361056a9731a8f", x"1d17f7652a098a9a", x"219a664ef10cfd9a", x"615b20662785d6f4", x"ee12ee401d2e1167", x"b99b99a865daf574", x"c9577a036e88d544");
            when 33193299 => data <= (x"d4c0a92ee569c27f", x"1137fe5bf17f4614", x"303a89b0c9eff2bd", x"19254edd24288cff", x"2ba0c76ec0d0ec25", x"73407a97cfaefba8", x"88c42b67c6c1be6b", x"e4d52f3232155f5d");
            when 10422327 => data <= (x"188c92f7783bd380", x"c0e21aa360d6f048", x"bfaefbc92d75b43f", x"4663a7bc2796e702", x"8ca7cae8626af4e9", x"726e646991263801", x"e40e8d688f591d59", x"08360355750513b1");
            when 19559936 => data <= (x"847be7c068a42840", x"8a799566ee292da0", x"9a24c7db8bb17116", x"b4fc6c8cc5d66e69", x"11ed58028a479666", x"545b4d4104d3520c", x"59b563ad91994891", x"164eb60f4403e461");
            when 14268568 => data <= (x"50de4206efc14cee", x"7727b82ff34f2f77", x"aa95c7c4d06ee4fa", x"e45a3d32c8243617", x"463ee22e0534ee50", x"6646dda9ae092ac9", x"240a0aa370813d50", x"f7cd20872fb221e0");
            when 403418 => data <= (x"842a5b41f9cd3c4a", x"9d306e1c3b2769a7", x"f2fd74152333a12f", x"04a46bce3253f873", x"42f9ace8e637c38c", x"aa04276c1637aed5", x"2e49619fe7f9d467", x"5690902f2dc6962e");
            when 28031892 => data <= (x"550272c0743ead80", x"625bb9a9ce23f8ba", x"6bf7d54b2e45c246", x"351c2ae2e7229b0d", x"65b8ffc0e50c43d7", x"6490f5f4449d167b", x"03daf1bdfb8d4bd0", x"f92b0edff57d9d93");
            when 23339563 => data <= (x"c3191294865f043f", x"1fbdda64ea822ab6", x"c66b47908031fa97", x"0695683d4be52da4", x"e8a82eef19d7d7d5", x"6d75725a98639787", x"e411a6d5f71c0e94", x"d822434a855a3ecf");
            when 16608932 => data <= (x"ff10c769299776dc", x"20cf3b76fded74a4", x"f924edf14e524e89", x"26bfa65af9440898", x"f8559a1bf8b2b385", x"85aa3c119a3420a2", x"5c15e4e6a8859c22", x"389cdeead5b7a65d");
            when 14214588 => data <= (x"71f384f4fd510ae9", x"932184192875a769", x"64bf47b97c227f81", x"82709b7c82f75575", x"2b6706389744e232", x"596f1a3d5239906c", x"9d17b1c1db4695a8", x"2f7cb3e1782d3121");
            when 29585894 => data <= (x"ba9948e6d19b9d0b", x"ff1fb3a3445e9adf", x"6f4c731782fd1706", x"d63d908780077609", x"504bd8acbafc1705", x"7951b50dbb941c2d", x"90507ce1e845f8a1", x"11696a946100af12");
            when 25941441 => data <= (x"88efb143c14928a7", x"53e18b3830dc9f2d", x"70966801fc5d13b8", x"206371e871c32177", x"469b2ac4ee802ecd", x"54c859b57a9377c8", x"1d833daaea6a6e0c", x"5d4ab76478ce07bf");
            when 24035505 => data <= (x"da345ad5251bef31", x"f0af8fe7cf0eb702", x"b6a9a8edee03d8e5", x"a3b9a26d5b27f420", x"3dccdbb17ea086e1", x"3ed6b272461f8364", x"83bd753ea9231d3a", x"4cde58d942772fbf");
            when 16776893 => data <= (x"34b72c06fb38740f", x"a4d452ec1e3bf92c", x"1f8a218331415f83", x"9f96928dedfeb4d4", x"dd587594ab5381c7", x"b74b1bad78dcb139", x"5a5e286da102df58", x"5c00e266256d6104");
            when 11359851 => data <= (x"9e5bb86fe4899917", x"2488f2eadd592cf1", x"8a55bf960fe17329", x"222046bb754b5167", x"2715e85518e88191", x"0c781cf4560778c5", x"e510292199f5dec2", x"d6ef03dd04d05688");
            when 18510747 => data <= (x"25abaa5279f3c105", x"6c3573649a573329", x"2cd0f7cb9c2ac69a", x"8bbcee02f513ff6c", x"e0de0fd7c525b2e8", x"a0817ccce2a68b5a", x"6e4593b735d5bd24", x"ac465700f563ba7c");
            when 29444926 => data <= (x"1958b924ae2f3871", x"b16189181e510bf8", x"85c29000ab2bb021", x"7197d7edfefa3ba3", x"b31169680195ed1b", x"20decfeb6424444f", x"eda473efd4fb4a6e", x"2b38db5a1f17b82f");
            when 24739840 => data <= (x"4ac8f91fb1ed2389", x"5db4cec0017c328c", x"49644dfd2e7d8cdc", x"6d2fece94e37041d", x"c08f1d8ad1b8e7e2", x"27ef3552f410f3ed", x"cb4c66f2552ae012", x"e3b88dd06276628e");
            when 3106303 => data <= (x"1e15aa32995d6ea1", x"6afbc686aa186f28", x"0e85cac0483e2355", x"29987ef5e8023669", x"f71766809a1ae0c7", x"0c1debdfefc666b0", x"f0825ca7b3848fd8", x"b2a187fa1f8d20bc");
            when 23084873 => data <= (x"6359b82061e8a731", x"3f6889ef488994cd", x"85abf65f1af43617", x"69c7052d9b1dacda", x"a85e0f073688bb6a", x"da00616a58d3fa68", x"1d35440257890198", x"65451d9cc7b75cf5");
            when 9436228 => data <= (x"6771899499b7907c", x"d8b6aae0870aa4f0", x"dad7c1b347a5a960", x"95c63e2c3e9e318b", x"4dc2d75f55ac8609", x"6ec01d83e25a74dd", x"0305bb8bba486304", x"1a94a478e974946a");
            when 15448393 => data <= (x"5b99749f16199eea", x"50e7a1175a900f5c", x"81763a9ee6da1ddb", x"b5ef0d076fec6856", x"d846b5e71d040882", x"5dadbe393b321d4b", x"993e99683e6008cb", x"056d0b6333bad3fb");
            when 8051551 => data <= (x"18db125fabc2d402", x"b67f6f8ecdd790f4", x"793fb9a0f118bb89", x"c72e3b135bb1b72c", x"ff289e0da60c93c7", x"381f86b08f320905", x"df70ca5bf508fa3c", x"f1a535448b732425");
            when 4813881 => data <= (x"956bd8fdde4418ad", x"fb86087185904125", x"2df29494908e4543", x"6c1bda1eb2003138", x"de9b2768807d778b", x"c66ced4bddae9076", x"0f6c3f6d83d2e506", x"d8f4bee854111aac");
            when 32711261 => data <= (x"c7483ee3b109b10e", x"56616774f04bfed4", x"797f6955fe0e5419", x"b0622d376282fade", x"a48b1690cc1fb8f2", x"85b155ad73795a4e", x"1b133eed99523b15", x"b6bc51f0545cdf96");
            when 23799661 => data <= (x"8f2aa3c709f0844d", x"43caafd678324f83", x"dfc3e0666fbbe752", x"567e61078bf156a5", x"6aba57a83c9c5249", x"574968cff6ee2763", x"800a3c860eed24a0", x"7f94c46edc80ce2c");
            when 18546416 => data <= (x"34fe0a043248fc07", x"f9fc8a175606f9ea", x"8af97c4d94c402fe", x"eec59bbdeab49668", x"d982bed659ff3f27", x"90a6ed5f45d6eeb3", x"23bd43ea4611394f", x"aee149ec8a813f49");
            when 28030272 => data <= (x"d08db9e123f0bf60", x"46329ff12749e177", x"46b5602398a890c4", x"cb3abd99b111f10d", x"e51fe70e1e24354f", x"3763054425c4438f", x"352f8c046d8b9b08", x"2b856e85b647ad12");
            when 3884689 => data <= (x"27ddb608a09c3985", x"f5f662b8128d2dba", x"6326f525d093979e", x"173bb627463e2535", x"360e630bd8d28b9a", x"e09728628f39c921", x"d6d8c4143efc73dd", x"e8bb1f9179619d94");
            when 14268580 => data <= (x"ed8fca7f361de401", x"fcc1f7c02fe3794d", x"b0266f50921cc43a", x"8264473cbd0c2721", x"7b7d0c02536bbc6e", x"9f69a8e32946412f", x"36450c70d163af11", x"94a83bbda69adbb9");
            when 8163844 => data <= (x"597e8f87e05467d1", x"64fa667a391a0c04", x"64097a665636e2d3", x"ecbef2984c357af3", x"f3134b8ff9161706", x"516b04884473df34", x"66fbc63958e2f5d5", x"773ee951559c42c4");
            when 24823008 => data <= (x"f1c58a36db96b521", x"4a27a0ce714f46dd", x"7a8ba454445e7ccf", x"21296a17db930347", x"aee74930b30f53f8", x"af1f9dd32b9e9b2e", x"fccd1de79a89e2bf", x"91f8c6cd8445278d");
            when 24712064 => data <= (x"960bca5f169fddf1", x"f391f91f42116889", x"bf42199c11fa8364", x"93c4ba994fa9d190", x"25ca266866d0b1af", x"8b3d3a79c93884fb", x"0881c78e429f0e6b", x"14567364331649e5");
            when 33578284 => data <= (x"c868820fdc42a33c", x"6eff959041484b3f", x"bf26455293f52cea", x"b73f47a71237724a", x"e57c72f566f0808c", x"1d730eda64938c87", x"4ad135b5ee40e198", x"a9ec7af2032c69cc");
            when 32028532 => data <= (x"1967f29ec43e5125", x"1d84c84f3a9906d0", x"ef20306c562da798", x"faef8329f1c6df64", x"921f68be29693656", x"a994d5e16efb8997", x"6566131bd8db65c7", x"1791eefda40e09ff");
            when 7510278 => data <= (x"d97740832a0af138", x"987422f05b1c3e33", x"e8ddbff4205b5877", x"a076c7205f6ed397", x"a8a0b4716b6e8dc0", x"8b8a2bdd16ecad74", x"02bf590dc8a7c0b0", x"5c9184966f4664e8");
            when 18227337 => data <= (x"4d9eefe3f2e18992", x"f07ffee37d032ed2", x"1d2f7a6a28a1bbe3", x"dd468ed749a6ab22", x"d03b3ebe6a4567fc", x"3b00227320727ef3", x"cbd60574c1d82d0c", x"ccdba15db8a93897");
            when 18379520 => data <= (x"2b56d2e3eba9c0e9", x"3d350aafc6314a3d", x"4e4b551633a23ed5", x"114539a3dd82146b", x"54ceaf11941065e3", x"a5d49d09b14c7c81", x"411b5294ea9e45d5", x"2085098e880ed738");
            when 25366906 => data <= (x"0260a16bd559c040", x"25a34fb81c494bd0", x"2e1349ba95685347", x"d2dc1744390dffec", x"b96305a0acfdb30e", x"7dbffdf34c2e0045", x"63047813e3b63422", x"567fad525be81d75");
            when 19178238 => data <= (x"2bfab5b6406dfa54", x"e30f468175887a12", x"02dffe065ab7f8f3", x"575689ae23807ef7", x"605cd27a3cee82e6", x"ea67357fb36899b7", x"28f7cf46eb3c1340", x"1ef52cd043fc214d");
            when 27501726 => data <= (x"d8612a89d874eb4a", x"45382bd605144d57", x"0ffbd37169f90f9e", x"76a322bbf595591c", x"7b12e287c86db074", x"f0c6a2e41e63743d", x"99cedf61d7ef9e98", x"9f5a3c83b7d369f1");
            when 1549369 => data <= (x"a81d2a1579ad7b92", x"aab69cd8d58691d6", x"77a650993c12cb8b", x"cb9c46889653f9d4", x"95718710a26bb134", x"de6aa8383de8930f", x"f3b7e80c10a675de", x"f6ba56c646dde25a");
            when 32341712 => data <= (x"afe12d3d123a0a2f", x"3613d3ef72737fa1", x"25486cfaca917402", x"487221ec762b3302", x"e794bdcdd72f7561", x"6e3a3b4ad9fdd862", x"f4e5e1ec95032bb2", x"9727945266fb6853");
            when 30255893 => data <= (x"dda34ca22a018437", x"656ca8f0872e691b", x"2960b32792b498cf", x"5f8680d66b15533e", x"93e04cd6faa436d3", x"a62120ad7e7c7844", x"93bdb0360b31a6bf", x"eea3a9ac984a8aee");
            when 32330099 => data <= (x"8748c3b7b4b0ad0f", x"343fca1a1ace50cd", x"b2eadd5159ec934b", x"88038f4a6ad554da", x"8b5f85cee364d2d4", x"0e0ca08b2c6b7b93", x"a5922bd7740314e0", x"4ea9c6326520f30c");
            when 21047790 => data <= (x"eeeb2e625e26353d", x"31635ff7dfe79f06", x"35999da8c2115079", x"1d6b9b201b867e3d", x"efedf86a2e6b7b06", x"be2a0088bc9a9373", x"49ca1f1d2782306e", x"f196975d3ebaac42");
            when 3196679 => data <= (x"7e866a75cff27838", x"e081f261a74a8c97", x"a560a25fcea9104a", x"325526de49723f3d", x"d85a446455a480d0", x"25f9b4e0d4351bd0", x"6f28ea58faf3b076", x"f053c783e8c45dfa");
            when 12171286 => data <= (x"d575ea3ac9d3a05c", x"70eafe3a5f331415", x"15ebaef94b0a304b", x"0c96f67114d14003", x"c77721e97cae9f12", x"961f7955c677f84d", x"93b0c502cf03fa0d", x"3fb575db401b977d");
            when 29268300 => data <= (x"8edfd0490c53001a", x"c93a3e6beaf77236", x"48599537ef67363d", x"525f7540f6c73cd4", x"8570fb200c3a362a", x"45b0a4151325d7a6", x"97b6c323c041d03d", x"c73e1add11b6b538");
            when 18800699 => data <= (x"9b19bf32d33cdaa6", x"9e0150db28f8bc80", x"7504b8abe8c79b2d", x"2a4ec1d85840f142", x"70746680343a20ed", x"4e2677b0c9ddd4c7", x"476fb75c36117a2a", x"67922de351924c06");
            when 5293497 => data <= (x"1fa5a6504681ec74", x"69222cb463625752", x"5a5d79e5ac5d5ab7", x"3d0af2cbd20265ec", x"1782253a3e04e0d9", x"fae12755176cc321", x"6de7dd5fec702a5c", x"94e060685cd581fa");
            when 22844540 => data <= (x"a771bcd1845eec02", x"db35bf8bed9b496d", x"14faf78e24c6f2fa", x"b07762bc809e7aeb", x"467c63fd1dc9c30f", x"87d8766e243976dd", x"bf26373bef2e857d", x"1843ee100fd04024");
            when 16951755 => data <= (x"e2dd246537b70909", x"454de3d55fd931ec", x"59596e3b8025500e", x"04abeaf61b29fb80", x"78b471c6b7a34c2e", x"77e90c8658747de7", x"60d4181137c80528", x"2047c77d14fbe3ac");
            when 32227858 => data <= (x"85dffcfbde7a0331", x"e00475adcb5c5f19", x"1b9291676b5db46e", x"fb45cc34de6671a7", x"c3a2b0813576e43d", x"2863ee661fbdaa4d", x"bb3ab5ee57973467", x"02f262cbeb76e7d3");
            when 28679767 => data <= (x"873179cd8abdbb40", x"8970c33750918456", x"a73d3ffffe960b7a", x"6a560a051870315b", x"bbe834674f4ffec2", x"1b20239bf46a7295", x"70efe3f8ffe05cd1", x"62046d82dd8e205a");
            when 10198350 => data <= (x"3908fa874add011f", x"2796505a4c4b9ffa", x"f65c5c1a4a04a402", x"da7b084b2acd29b6", x"b6741b298333c0dc", x"75bebe9e220558ee", x"662467468d500132", x"74a5200be02870f9");
            when 33857880 => data <= (x"3eed4fab004fe32f", x"2ba257f2f1dcb21e", x"ac22700d263941b0", x"2acd465fc9b0e207", x"a7b163a1ea14100c", x"dc1bda46edc1de2c", x"105f0c775d39aa84", x"706f30cba0f1bdfc");
            when 29209635 => data <= (x"74de26ece210a144", x"c2b67c2c1bfbeeaa", x"e0e6b1309947fd9e", x"653bb030a35b3d2c", x"48cd9abc52377a7a", x"a52e2a1110452705", x"2d3fb0cccfdbdbdf", x"9adaafb446e6c2f2");
            when 16299456 => data <= (x"33a425215f6593ed", x"274ba09e7bc9f2b0", x"f35098feec52798d", x"f98176dc68c2af11", x"6a97554b19e1b594", x"071b4c6c5b79ab77", x"142a248228c5c582", x"4c024c7b8466cedc");
            when 33249363 => data <= (x"fde648f45f531a60", x"edd6871848883486", x"540ba7e6ab392c11", x"e630e3c7589977b0", x"ad4fcb7bc695fb44", x"7051a8de5a6d6935", x"3e4699f2a6fa8afd", x"4685bcbd1a3da199");
            when 3986038 => data <= (x"d85a8215b19d3071", x"e90ae8c10c707052", x"99f75b59746d47b7", x"47179831a86d8b55", x"c59d92c7e508c1fe", x"3a7c65f1bf45d448", x"b4272483a207d7c0", x"1af7e933f597db7f");
            when 21447367 => data <= (x"f01426f95731f3e3", x"0df61d8045e0aa67", x"2e6b5fe54f63c6b1", x"06550556d98dfb5d", x"a0a7e22a6034d58b", x"561897c1b833f7d1", x"a536accd6f136fe6", x"f328b53860b8f639");
            when 9242239 => data <= (x"9c560f49fb91857e", x"79bbed3b998e2634", x"1d75742188ca0253", x"26532868305dd965", x"bbf01dbff7f5ef83", x"5d9dc40317782633", x"5276d5eedd1b3349", x"0e16e9f0e2f0516c");
            when 21122335 => data <= (x"7c980d2d901ea5f1", x"30206e3cfd7c280c", x"af509d454336f5d9", x"236abf0db64963cc", x"42c70f46494b9242", x"d0ed9a0185b930e8", x"0f77be00966dff88", x"7be09df3d02325d5");
            when 2519493 => data <= (x"1e9e7ff8276fad50", x"f681a5243a2d03ee", x"d766dc6a41fa98f4", x"4c71ec9a61765c75", x"09009b60509ac6df", x"1d91972217298e41", x"4666bf8d4bb8ee0c", x"fc554c061c8e3bdc");
            when 2588990 => data <= (x"6a5754029ced7a89", x"80c88f55b14f59b6", x"cca4c5a1f17a2584", x"a32ca1955b755898", x"6ee3d69e1872e9c0", x"0583c2cdd9c21bae", x"00a57e64951cbd7f", x"ddaca4f6fd365230");
            when 23776575 => data <= (x"b0aa3c1b223f7d70", x"ad6c9160df3fb25d", x"97888e6fbf4df538", x"90a92e48a4a2c971", x"1318f4bfaa3d4692", x"ec9f367a814f1d15", x"e98bd5b0ad4683bb", x"d2814f393c51abd2");
            when 5435792 => data <= (x"0b067ff66c3af912", x"254a5effaeb51eae", x"13e2bebfa5064daa", x"c2e34bffe8bdd6b0", x"81bf0d7c440e9fe4", x"bb8cc550fdcdaff0", x"71ec040a17983469", x"bb1d321b2c791059");
            when 31338448 => data <= (x"454276fa72a28971", x"e9fdd6b0a0406457", x"82494a4920775ce7", x"b4dfa621388e2eee", x"72a82caae80356d9", x"1a709d712867274e", x"f00220c7a88a3d0a", x"3865c74431878d7e");
            when 21691724 => data <= (x"570bbabfe9236157", x"9153a35dfa15880e", x"a47dc7c2f9c562ce", x"2e03f27671920a04", x"6b54d2b00fd47e83", x"c54403b37abb11a3", x"c6e62d39b0be7ed4", x"a2ce498205c1d055");
            when 1501828 => data <= (x"23b1ce5f75b5df84", x"04d73e2e5984cb26", x"f6317d11c9b2b4f3", x"7215261f56add596", x"edfd76aa494ac0cb", x"12ff1e943f9561bd", x"2ff7434e6720dd53", x"ab1b003ca64b320b");
            when 2419607 => data <= (x"2f268c5dfa6c1a3c", x"6da2af796b5c1b8a", x"a26026369463bee4", x"e69e98f7321b5f29", x"dc85fe069f95bb94", x"89a87bf276c377f6", x"427d97553bfaf706", x"7300abb277e5ff09");
            when 23869114 => data <= (x"d5b99d58399c5791", x"22c0cb39e718deea", x"07f6c27c86b939cc", x"c7557a5b8568a5dc", x"4d7ff623d6c3982b", x"508850c0e32e6341", x"822abb8d74bbc9e2", x"9d19488852f442a2");
            when 33063530 => data <= (x"1811bd13f27f82ca", x"8c6d921b7a9487c7", x"069b5bf59abc8f4c", x"6a5b3e586b710c85", x"53f01398507f3a9b", x"f041104c9f43ab54", x"bed2b1601c879659", x"3a688f58c924acfb");
            when 18342050 => data <= (x"a24058172d09d8cd", x"ead62968a7872ca1", x"5d6cbd2f014d1620", x"e7b88c253fb40c7d", x"10e7002fc08f07e2", x"d2e1968e227e48f7", x"560072e60a5f1d72", x"f19a8ad502ed56db");
            when 25678146 => data <= (x"4eb5ae19bc4567c7", x"1171587845c5f0a9", x"ffe3284cd63b89ff", x"88f814587812d753", x"29eda7b5b9ab8ce1", x"0e99bdf2bdd47ec4", x"466a7fd93db9ad38", x"a17729cfb185b913");
            when 30085926 => data <= (x"7d112b1709997736", x"ac6cd41b03ed3d65", x"f5d3675bb711fd22", x"0cea9ef9a1889d1a", x"901559dd8b74705a", x"a765861f910c5a53", x"0ad698714fd91ed6", x"5ac092da24cf2674");
            when 756396 => data <= (x"18c67fec0dd3a86b", x"e5aed65a97d7930d", x"9d6f61d89b076f58", x"474b431ab4fe434e", x"792bf3318f7853be", x"cf7305fdbd7f758e", x"ba18b8a39a61101c", x"d1800d7b8d75a7e6");
            when 2482448 => data <= (x"27f27c600eb5f01e", x"131768ba2acbbaba", x"e64d86506ed51436", x"7c8257b559a38dde", x"eb7ead15549311c0", x"e9c2638b24d02b69", x"feaa95d0de818182", x"5c1772e33de297b6");
            when 12138458 => data <= (x"6fc3f675051d9873", x"ba330fa24fa1086c", x"f4e90d9313619940", x"5ae3dfb22fc2cc05", x"36eb322c8cdcc98b", x"34d34940bf9035e8", x"94f36b2eb90712ce", x"6dff89efaba24454");
            when 15252237 => data <= (x"7ac398108d3b7f46", x"75054463272820b7", x"d6a82e7e75adc123", x"fbc0fc3ce09299c4", x"c85c494c26522394", x"7c58ac2a465bffe9", x"f6ba0b1ea43212bf", x"ff67fe48833bec98");
            when 27443570 => data <= (x"a27b00ce9b7c8608", x"c51e9fa136caab40", x"f2a5d186d42eea4a", x"6e71b28b5d8778c4", x"0ea1fcc5c7d875aa", x"62c3c69846bb3752", x"59c5f066fb0cbc0d", x"da1fb35ec6d1d3c0");
            when 17372618 => data <= (x"df072fae8aed5101", x"a1a3c71dfd4bd930", x"495b4b6dcab6311c", x"10a2ba71d0110914", x"ba1bd690131f9cb1", x"5bd22727b3ead31f", x"9f39da27842ee258", x"5f5be6059f50bd2d");
            when 2045795 => data <= (x"af735eb1303cb97a", x"c35a5d68a1c9ceef", x"0ff7b214f957e8c8", x"7615f9bd5379b5b4", x"5d85913ec74899a7", x"b3342ce99d0983cf", x"fcc4bdc7a374af40", x"009b1c4d0abcd43a");
            when 1028418 => data <= (x"4f5ef2dfd5f520ab", x"d1bd4896666ca338", x"9b45d7a7e87e5c06", x"86a27f5b40686d9a", x"51fc14349901b614", x"2766f0bb7941fe84", x"1873445e61122d07", x"29c31e72ff1811f8");
            when 18586652 => data <= (x"288e3733c9dabe68", x"38b2ff8829acb4cf", x"cba1b7b70ebad992", x"6b58d1852206c40c", x"690cd5c87d7ff0c9", x"938626e631f529ad", x"ec0c7bcb8322298d", x"b565f267f6950079");
            when 30313542 => data <= (x"301e2a2c54425c22", x"3e8ac03b27654d31", x"49405e20e7fef084", x"c25513ab4dbaf22e", x"8ae6557be4c5bbce", x"762657298b7af879", x"2e5050665be02dc9", x"2a43ac2c5ab4261e");
            when 24156477 => data <= (x"cca9a4b7aefb98bf", x"76da54426713da18", x"a98ab40101cd50ea", x"a781d4b38c9c7d87", x"4f2ac6a675716e4a", x"d78e15e2ea951de6", x"c17ec840dcfbe710", x"53c760b7a5736080");
            when 19399229 => data <= (x"9a9158647801d5b2", x"5437b88075c8d8bd", x"32c3e92993730523", x"2c150f56ee6c3392", x"3fa596a2f90d5ed7", x"c30b12411c4c8e5b", x"c3bb0965a6b3cfb8", x"7348f27eff9c5f02");
            when 17693278 => data <= (x"acbe44b14212a52c", x"89696fcd9512ea37", x"ea9fb2f91eac66e8", x"92e428f0f7e3bc66", x"ec91aa1a261858a4", x"5a34e144bf9bd898", x"eaeb2f9e9a6acc85", x"2c1afc71959b42af");
            when 33718626 => data <= (x"47fb79b43ce7b9e7", x"b73be44305260548", x"2a303c2821eba1c7", x"f8d943c22b8a56b4", x"019a155dd3f864d6", x"5394b6ee46bbf3a5", x"852087d99d710982", x"f02a2fd28d0d6980");
            when 19104029 => data <= (x"b6743a5ce3fd9d5b", x"b3576fb37f22468e", x"a4f89de9057171cb", x"2a1e02d1bc9e3384", x"6e8a3e083c7ee16c", x"361146cb4c8aa156", x"6002ed8f6de46faa", x"46fbbf696a8420a1");
            when 27483748 => data <= (x"6c1dc3be454d837b", x"131a00c67e67a88a", x"6a09ebd582adcc92", x"f3faff836f75a422", x"27bd534c4eee18b8", x"5bb7ccba03944cce", x"5447cd4302f5451f", x"2dd70de54bcd5b83");
            when 16035868 => data <= (x"51e6296838d95aae", x"68568b92f2ea9ffd", x"ee45800b0e99bf86", x"729679fedc07d0fa", x"69a6f09dc08df4b3", x"dd8679878eb634cc", x"ac732a59333783e4", x"5851ac7ec3d5a51b");
            when 29078933 => data <= (x"ae1e00fb07f6b21d", x"315fb466331ec251", x"38e11884cf1f5401", x"9555a9415375774a", x"683873517827c966", x"99d46fb91486ff83", x"f759bf5d77a04033", x"e46f4d95f4375bb4");
            when 2779368 => data <= (x"49115eca3e9bcc23", x"e947e2e5de261d07", x"a3286ac9af6dc70e", x"b5d2315ebf6f2af6", x"2ed713f4f7886553", x"a73a720337eb1258", x"c70a10049e9f0779", x"942d7d0762d4d233");
            when 30074634 => data <= (x"3ecc90dc50bd8fd1", x"be400b70801ff913", x"c39dfd2e04bfedf7", x"4e4af8f2cd4ecd36", x"4e2f6fd75fe15239", x"a5ea2bb78d292323", x"d392edf84cae4b2c", x"8dc83cfc58b0055a");
            when 15369846 => data <= (x"44d4e3034a378c58", x"acc6ce5945469f5d", x"ac66f870d8552310", x"e4b8c92662e24784", x"9a84ce755b0e5870", x"01be4fc54aadb144", x"c1ba4e396bc6df3b", x"78b99377f5f16a1d");
            when 23111353 => data <= (x"56031cca83e28f1e", x"0b69206044304aea", x"2a89bd618d965eb0", x"040a0f36af965c12", x"a6e249a70cb25224", x"ef1be5476af2b8f1", x"e83e34953988c1b0", x"9108f42a5df59e11");
            when 22333773 => data <= (x"f86cbc1ad891c9ea", x"710fe3a68d8f0b0c", x"7e05b3fa211fcf15", x"83e3246e63449e05", x"c21489de7c54a74c", x"cfc01ad27be7f246", x"40a4d7a59b5382ae", x"868882aca322486c");
            when 33756140 => data <= (x"fa7d2a92b17be805", x"1e62adf4815980f0", x"65d83a36c5cd673e", x"4772b7ae12fdfce8", x"f85580f36c892292", x"0abc470998b9fee4", x"173244fd00587b35", x"feabf59e9151fa88");
            when 19820724 => data <= (x"8c0ed5ca65009978", x"d73ae05608755b74", x"b75fb62aa53ee29b", x"e51f3d1f0c35be4e", x"005689d170b9d515", x"1a07690290464fc8", x"6d1c0416035776ea", x"690f8605cfe1c83c");
            when 16611399 => data <= (x"97dd95d1cb2882b4", x"9dba62c3bc2b99a6", x"6306b1f9720bf747", x"f924147dcb3bb706", x"7a05e756bbe4d806", x"34e9a83ee84e051a", x"a6059e4747c8f52a", x"ab4ed79dd9267342");
            when 29592460 => data <= (x"8effe60849a8bce0", x"b69bc6823169f233", x"f37819081bbc8e56", x"b342f4947dd40919", x"bcf4a4678fb194f9", x"229a3f973ebb2e58", x"8b1638f45f4f7724", x"ea3f8e3f0b309b69");
            when 19289025 => data <= (x"68f6cda47e2a24f9", x"09ce8f1a2fdecc03", x"6bce9a3e57594518", x"2c56808d5d105806", x"b3be9ee08a5f3f26", x"092d9c81552f46e5", x"46b77fabb1fe245a", x"1b3ffb59b6175400");
            when 19449788 => data <= (x"bccbf202d65e5168", x"43c34e0890c984a2", x"dfffc6829d91ae9e", x"64d19a9e17be5365", x"b024295b50d46689", x"9d8247cd2b6d5824", x"e02dc48004b899f8", x"0ed3db06c6607071");
            when 1327412 => data <= (x"27e4934f4bc0b67c", x"c7887d767dcaf95e", x"1bebeecc9aefee6d", x"d26d34bc86773740", x"14f09d5db68ad3b5", x"e42ef3c1c33e4f3f", x"75f46c37d593e42d", x"d08b92be5a3719d3");
            when 22270655 => data <= (x"1d143e7c57344626", x"afbc67417e8cbf59", x"9fd874cdb56f7c83", x"a6ec54b46bdedaff", x"6f7c4d7106faec22", x"265f776e0774d8d9", x"c801f0547130f843", x"9bf1e9042109c413");
            when 22676942 => data <= (x"52c2f1458823c760", x"7c9e5b558be1c4a2", x"248a90b10bdedb74", x"2019b45b3789398a", x"2926a670d6d94529", x"cfa1f7c0d6881512", x"a9d71ce9fb141546", x"6c0edc0310bfe0ea");
            when 7379426 => data <= (x"74d4ff8f191e5572", x"400570f5dd93cda2", x"f6e9415afd9b1f6a", x"4259e750e0265962", x"43eb2afe1f5ea4eb", x"75c41d1a2ac505ec", x"3ab8f1de3a19b911", x"75e4e51866bff8c8");
            when 8896531 => data <= (x"aafdca04c61f61d0", x"48841df593c5eeee", x"fe283d9c007dc5e3", x"50519d3fba2bb299", x"b5fb96ea4e90ca24", x"b11c212b724c7d3b", x"19f7cc0407dfaa73", x"3d5227d66853e041");
            when 19506665 => data <= (x"dfec44c1bdb74673", x"537a31afd52a1112", x"b5efc8cedf3ef768", x"4f303f6b3bb51720", x"b3a3db41e53f6975", x"ad7d6545abe071bb", x"c1ca9cb2d746adc9", x"263580418fd5b412");
            when 1724410 => data <= (x"8e7315cffe7c65b7", x"7d28db75dda5050e", x"76289f549817d719", x"5068f2294d769454", x"03ea1c1a3245ea01", x"d7dc5bcbb25cdef4", x"ce846338abded838", x"6608906b44d7be03");
            when 21476719 => data <= (x"6d6a5adf154b9fa4", x"f95411a370de959a", x"e587e88a70dad546", x"30b9568cfe379c0b", x"48fa4bf9fe3cc439", x"001de0462eb3bb9d", x"70f314ba00bb2780", x"30fbaaf5126d0ec5");
            when 24037576 => data <= (x"2b580a1dbbfdcff7", x"c170eebdfc98bae4", x"333c02c4d09bf7d9", x"722200c9dd35660a", x"356066e1fd9bddd6", x"f87eca1d3f27932e", x"f8f49c507a80a8f3", x"d4ef03f299562a84");
            when 26326710 => data <= (x"4b5fdf93872c8e8d", x"0186ca2451d1635e", x"42bb4a01e329603f", x"1b6f49386b2d1501", x"d41eab9b33266f01", x"85ca77bf3ede7584", x"9cb99723ac73996d", x"3ebdd28261e62b97");
            when 30920294 => data <= (x"793ed6dd49e0a4fc", x"d3f0a2a86efd037e", x"25a5bd39dca71675", x"699fc312cf459acc", x"01ce84574969cd11", x"fc34b9cb14c3bcd6", x"2ef71f723e81eb46", x"b9ea182f6d82fe4a");
            when 9632789 => data <= (x"51f054510c097487", x"d4b590ec16ff543a", x"5f453cbe8bd967a7", x"cd816c7c25b9ad0c", x"fc240589fb89d633", x"270eb43d848b2b4b", x"b420a710e46ce691", x"d8518cd27219e2da");
            when 9849210 => data <= (x"cff82ae949040aa1", x"a74a79c4e9b546bd", x"65fb748185a396a4", x"f15e0a6bc4d395b6", x"ba26f95cada256d9", x"e03010996fb0af59", x"d07cf0f6e502cf53", x"cbfef85bdde6ffa7");
            when 3010712 => data <= (x"a4c6249a79069f33", x"d1f258a026882dc9", x"8a4a06f48ce65e7b", x"4cfbfbd2e52ba37a", x"814160aca0a016a1", x"6125a49dd998a8e0", x"45839f1899a2e067", x"e92a47d143d637f4");
            when 12783206 => data <= (x"8bbbb101d023562b", x"9e8370502e144f05", x"b247996cc894e326", x"4cee824af6271fd4", x"77433a037f5e8d58", x"341ab5b4704206d6", x"e96614d58ce33c80", x"0c67d8512a341f96");
            when 28798419 => data <= (x"285c5bab696b74e1", x"552b2f57962f1c94", x"12f02d32815261f1", x"101e6cd81b4e7991", x"615d8e0054fd1c40", x"cd9f1681f9a3d0ab", x"e841f27e03d8bbc2", x"d6daeb36a68bce83");
            when 10190398 => data <= (x"1e8ec6688b9d250b", x"d169a60b91289043", x"bc470f643ea4ba4d", x"d135954a93ce01af", x"52fcead043d33934", x"1fd0a33201f2c8bf", x"8f23512276b6d4da", x"16ab7b917af96522");
            when 10504566 => data <= (x"696f4fa4b92f2f5a", x"0f6f74e37a8ae2b1", x"8d21e6c773d754e6", x"f1a9b831b7eb3390", x"bc4c1527476bfd62", x"fd29804505d50e57", x"617f1969501afdba", x"494492b57cca91f0");
            when 23406342 => data <= (x"8b7df8bd5d3c3c5c", x"bcb14ce3e498abfe", x"bd429cfb0ba481dc", x"291e4e24b937e4e2", x"2c2188e502b0190e", x"c0c1c09ed84d6b1d", x"c2af00dc0cdab623", x"e2f0f30181cc3e16");
            when 7866336 => data <= (x"8b5bd46e0c9350bc", x"50d89586323e3234", x"55ed1cde0bef065a", x"4bfa87f1a226d1de", x"a1c9cdca5ead924a", x"ce40d47f1e61717c", x"d4a87ba6f92d1f08", x"969082aa5c8a91c8");
            when 8802037 => data <= (x"26d9ac16b4b4206d", x"538a10d235dfdc15", x"45bc2ea386ceb247", x"6cef6777d38aa714", x"7b0d8d8abd9c9357", x"2332a9174463e04c", x"19c349217f2834c2", x"ba179af646188f6b");
            when 22105590 => data <= (x"288c0889bb49f347", x"eddc9c07b73112ac", x"c91a1cdb096a27e8", x"e6ec467bee67be2d", x"0032128dc81f2ba5", x"aba5e54208782c4b", x"b5397fb95b57f20e", x"3da905c644a2b0ca");
            when 15710427 => data <= (x"6860471c3fedb8e6", x"79595d50b5176650", x"da192df30541fd24", x"918054113459c573", x"7ccaf5ac018fc145", x"3e93f0a54d8fe533", x"86d902eb6968dd86", x"cffbda2d794b2421");
            when 25157454 => data <= (x"24ea70e8d14700a5", x"7ba7afdcc8eefbe7", x"6f38cf9df3f210a2", x"9be4725293c48e37", x"6a8eecde48b902b6", x"5a9563ff1f35eefb", x"31dea171bc0277de", x"8825f22c8012bac7");
            when 8943052 => data <= (x"f8d7379f2cc3b903", x"4bf7d09c8e062525", x"4530a53296deb31d", x"c5c47276447d54c0", x"27bbbf0ce36481e8", x"207f3979ebedb218", x"7d70e704c9f35d0d", x"568a0de0708602d1");
            when 13864968 => data <= (x"95739ac61b576c32", x"ac80f76ff122ff9e", x"e466f423033df9d6", x"457a4730fcd61faa", x"8d7bfd9be56fb3b2", x"450cee5e6d029bc6", x"aa9cdeac9c877a59", x"4e790a12d29b4d8a");
            when 27624331 => data <= (x"0139d912d09eafa3", x"c17d494fdef7e194", x"3564c3b82fc4e5c3", x"cf4f7bc5d5cf683a", x"c9e1aa55298579b0", x"c40e82275e68a81d", x"4c7619414559c589", x"9e368c60b7d1af18");
            when 2265626 => data <= (x"80246159f65792c8", x"f95277a0d2054f78", x"3eac26d6fee1718b", x"3ef5772579472813", x"05a0c9af6eff3790", x"038d3769c9084c1a", x"3b8ec04872420b6f", x"01c1017e824b7407");
            when 4640064 => data <= (x"6260cc07fe8eb29e", x"1662d8435b91bfc7", x"2977a6b119e25787", x"7445f5fc71aacc99", x"a552ebed10d7d074", x"753876b00869619b", x"997bcb2aa6a8e012", x"408c5ba75fa5c592");
            when 3081277 => data <= (x"6f66a2452aa02ac5", x"c11c21402ef877ac", x"2c0dcdfcdaba85ef", x"90a5aaac3c7c3230", x"e90be77f01ab6caa", x"c7f34c68fcca4a1a", x"7453868f0194e26e", x"5dcea10b75ebeac7");
            when 28677499 => data <= (x"e3d28c0ef81e91e7", x"95df99a1c7093fee", x"9fa190b395de845e", x"59e851cdc75f8a90", x"b2f5990c63c69012", x"dabb5f077bf03ad4", x"c7e9400e4bd9f64e", x"1bc2eebb239ce2bc");
            when 22413967 => data <= (x"bd201cc932999a6f", x"077f4f1ed9c1d0c0", x"a360f923fbe3a51d", x"89f2c85e13fa81c5", x"bab547a8bfe56a53", x"a1b44a46487de599", x"19133e85e1b03cfe", x"81cef336a1db0ac7");
            when 28482146 => data <= (x"35d27e2c57ca59ca", x"72015864ba564ff1", x"25adf6f27f090e55", x"e695905eb8c455d8", x"4a93482b2f3be45d", x"0eff607dee5d79ec", x"02377ef453e8dc96", x"0ac307ac955e2d2a");
            when 20594275 => data <= (x"663697934bfee4dc", x"266c43de1b0a7746", x"da2127db972bb324", x"f45f85ce0790311c", x"d15a6138eb084ed5", x"559bdcf269651c89", x"1244c824bd627a8d", x"d1280354eafdfd6e");
            when 7403334 => data <= (x"f0174d966e272f10", x"3d68a475959212e2", x"eaaf6fcffbdf2fbe", x"4a6335debe69b63d", x"590221bf8859b43c", x"4217803e1c9be6ed", x"fef6251ae3524449", x"2b35a4939b5182d6");
            when 18875185 => data <= (x"91a4d0a77132bc8f", x"0c6127c76fe930b2", x"ac83963aadb3e5b1", x"4d34219341c9764d", x"0f730146ceb360de", x"806b740a2fa38a4b", x"91380942ea75499f", x"eb0b5c423ca3dda9");
            when 7034362 => data <= (x"c705f8a8dd876c0e", x"703ce0f5bf1c5029", x"c4b72708be532056", x"4645f53c632b660a", x"2ddaf6d9c0acf463", x"55a86cdd2836b45c", x"b14c687e6de5f1f8", x"cedb170868b5d1b7");
            when 12075929 => data <= (x"dcf3f569cc198d46", x"757207463bffb50a", x"ad1ea2aefb8e854f", x"38ae6ba8ef66d295", x"3dc90ba6012954be", x"fd1dbe5d0193cf58", x"69f58df81b66cd69", x"ce8135148f0c71f9");
            when 13846384 => data <= (x"ee43644d92837d9f", x"115f3fe2a989407a", x"1e65f2fcedb1852e", x"4133ffe5a3b07691", x"071c33345d1cdf71", x"d8ec1b5c7d4c5181", x"c94b792e1c6594ce", x"b9aa1221a886b4b0");
            when 27263552 => data <= (x"21ef3d2237926142", x"b0dd608ff8a5d1d8", x"8ef844d900c4fed0", x"ddebd3cda589d5dd", x"5b2d26325a39bc0f", x"17ee41c0b3677d10", x"eb63314fa69ad12f", x"724b66614fb3cbcd");
            when 3264913 => data <= (x"4765d04521c8433a", x"8e7da4c75c5fe14b", x"3b786707700ae4f6", x"da060f92ae537bc4", x"697fdb5ad78bb384", x"5e604d605f74211a", x"03fa017828d940fc", x"4b56ca474d9cf047");
            when 28736957 => data <= (x"6f52bd53207ba8f0", x"3ff153696834a277", x"7de3c856dba68362", x"3595894ba9d1b839", x"b2bcce4ce3faf927", x"0f8c928840279d71", x"1239040f759396db", x"bdb772b0f574925a");
            when 25641095 => data <= (x"12253c41e765093f", x"70d07e0f2293eb92", x"db414eec49720ccf", x"e41a0b409a37db04", x"cece0f521b0f89d7", x"5cd2c4367d296753", x"a54afca633a14e41", x"6d3309b2946f3f90");
            when 31948086 => data <= (x"2b84caa08ac9b8a6", x"886f3e05a3667514", x"eb060203be6b4b12", x"1216ed0af3d914a1", x"9285649e0f480195", x"e5451b03e042b2ed", x"d3beb5bb313d4336", x"fc049ea2669b1c27");
            when 23660452 => data <= (x"001516ab78dd58ca", x"8e7756a4d41da29d", x"4ae6edcb2e6bada9", x"c50738ceb2836dff", x"56f0f0882cdb42ce", x"c46319c17e18a16a", x"ef49da0684aa0586", x"64f6447325be1300");
            when 30053141 => data <= (x"1e05360d54576be4", x"ae6c69b48092d461", x"00233a5f860caa8b", x"017bdba321501d34", x"a06f857dbcdc9c49", x"bcd6d9217f0a8012", x"eb3e67086fd808b7", x"d294567321a0cca5");
            when 834522 => data <= (x"6d85a6ef745ff79c", x"20d0b03b7e35e6f7", x"c1fa66811f8104a3", x"454daae4fcd2f53e", x"5d0b00941400879e", x"3a6096534ce02215", x"326f6373d7e3a2c6", x"e5742f765d5afd7f");
            when 15528419 => data <= (x"d88620c1b70ddafa", x"2c6a368903f70d47", x"1da79a4b1319788f", x"119c2e25ee036196", x"947f77bba839ffde", x"a28341d012028b25", x"fccd49deea0d34c6", x"7562237cc202d77f");
            when 6642959 => data <= (x"6b00b765ccb7cde1", x"a6a98e9e464c8844", x"ceaffd9e694733f6", x"f43dd555a0f0ed02", x"1450e8e9a35fd0b1", x"0b290968665063e0", x"7b5a5412b607c950", x"6702c8f1bb09938b");
            when 16148409 => data <= (x"47e67ab41d36801c", x"09a8245a34075cbe", x"27d10c991323cee7", x"70bae42a51490bf7", x"2fe12352d920ec77", x"e7ad481a2ee6e8a5", x"501e1941ffc57a79", x"b6d264269f96f4bd");
            when 29212590 => data <= (x"8573ed0cf26c6dab", x"74b5e2f5757f22e3", x"8c8aadd76ce623c7", x"6462cb6c7a9cbacc", x"1138be8678dc8250", x"f21bf10afdd84c94", x"e29241931d6a9681", x"e39c132d3d04ea77");
            when 19926435 => data <= (x"2cb6cda0d79b1364", x"bad8994719284631", x"92390288bafa652d", x"f4b29671250237da", x"d5ffa6357c0ef8ef", x"71a630988f38045b", x"53d0a560229ffbdc", x"6fff3b7acf2f6151");
            when 23284438 => data <= (x"5b10da2e40d5dfbb", x"b58f303a84ff281e", x"efa922f1022eb2d2", x"e2c42566a51a3adf", x"88fcd5486615995a", x"6a2dd0a40ac5801b", x"abd6d4fd67e3ba4f", x"5de3a8dc3b870eee");
            when 7684940 => data <= (x"a40dc59950fb3ad8", x"29fed813a38ddefe", x"0074c0b34e91254c", x"c0832ea6444728cf", x"89c47130f9fafda6", x"8228f8462d979b44", x"90a8da2094ed3080", x"51aaa4a35184c8ba");
            when 12476254 => data <= (x"b2a9c4ed3f4dce92", x"c5bcff6e39af842f", x"14b63c0e67ebab75", x"0a80d303b91dc328", x"d3b0372290592e4d", x"5204cc964e6d93d2", x"74e46545f6866a9c", x"3386c884d3bbd665");
            when 29649278 => data <= (x"d5e91a0e461ae683", x"8b83f9bf38f55408", x"3cf2ae016031f6d0", x"c6a5a6b0109174f8", x"8bce4bb457772a0d", x"6bd33948f23b7613", x"d0a792caa65b55a0", x"4d303a1e4d0bfb37");
            when 573220 => data <= (x"5c51b7dc302c2fdc", x"425a3f3061bdac45", x"0e1b5e902254a8b6", x"6bac03925eb54296", x"05ddd7f17c4c6354", x"641e0139d22c8d40", x"f37e6fe49797775e", x"711cec0602a0c29d");
            when 9672283 => data <= (x"7440ba0b184f2caf", x"1dff9e506a7870ca", x"737d2426f5e23dc4", x"60d4f2f3f9a7c69b", x"e756d532089ef3e3", x"97ecb7687438d664", x"24809a43e393afba", x"38fd0fb0c5f3dfca");
            when 26696017 => data <= (x"e7bcfa9161e4c629", x"717b5af51ffa03dd", x"64797f1d98c808a6", x"1229d7fafcfbbc98", x"35af23d09822461f", x"fbb53c9b01aa6559", x"79a8d69ef12c8dbd", x"5dced78c01a827a7");
            when 9018155 => data <= (x"48d4a8a9a3a425d1", x"bace8d566e572495", x"605dddcb80e352db", x"dc62f5f0c935d50e", x"458f12385c57dd7c", x"31d6feab303848c2", x"484b752d0d75ef96", x"fb423e2347e16303");
            when 7885487 => data <= (x"129aa1dea1e8d03e", x"9dde3a865e54eff0", x"855bc41c17380b9f", x"e11dbdfe6075d497", x"8e03ac455e780991", x"85b00f60fc8835cd", x"6a5be97c18554fb8", x"21509049f6719058");
            when 25858789 => data <= (x"6e9aa480f664fe7e", x"647fcb10e94edfcd", x"7c7f3bb4238279f4", x"5d1fbb8408ed5077", x"097270dd5df10c64", x"47d94a80d92a4aa1", x"5ae78946357bf199", x"57ced976bb7ef231");
            when 2376221 => data <= (x"aa24d18c0cdfbcab", x"0b0c356c13eeb0e6", x"06c2bcf3923a6eb6", x"2b1d4a659ba408d9", x"9e58de4bc0e61a42", x"1eb050ab15396cb3", x"182758c89ec7d057", x"b0a1fcec733245a2");
            when 11470061 => data <= (x"7ad3791da518cbbd", x"8ffe4984b2e0efc1", x"8fa21ed7c1e92803", x"86e69a330c272b65", x"d4562603935e646c", x"f1964db8e80ffc06", x"548393a88b811f7f", x"bd52a89cedcaec19");
            when 27287006 => data <= (x"b2057986d503f785", x"12485ad91c43d802", x"fe338c84f402b919", x"8e73027f526262ca", x"b8905e27e10a7df6", x"60cdd1806117c56c", x"5c97317b260141ae", x"44a1538db2fcb6ff");
            when 28817789 => data <= (x"59509a2cc421f6d7", x"bdc18f1e703673b6", x"cc81f0a381e6646c", x"30642deffd5ed6f1", x"1a450c8a584373d5", x"aec20c2f8a512a7f", x"b0003544a414abd9", x"034253bd312cd8b1");
            when 15852851 => data <= (x"39ad887f55308ce2", x"b9f743ed68611e4c", x"676d521fdba6a1a0", x"4a72f7a6c018929a", x"d1eb8c88a4fa8fc4", x"767f15d00a8fccc5", x"5d51c2cdc5cb07f0", x"1ea62eedc985c3d9");
            when 29804938 => data <= (x"bebbdb23a526ea9d", x"b130fa9cd24ceb73", x"f034dd63b82fdb80", x"b246cee6ecc4d06b", x"13b55c8e64a828ba", x"cbdd92939357a329", x"543f092b88da396f", x"8a531045f5fd3d4d");
            when 8380654 => data <= (x"74130552402f9a71", x"dd759eadaaf3bbf7", x"6a5891802bd3748c", x"f3552cdd4596526e", x"ae198588ad4001c7", x"e26959ee1f3289d9", x"1408393285ea5987", x"49ce390fdc92130e");
            when 31586274 => data <= (x"e4379250452b769c", x"d9dc2e81515ad997", x"71e543ca810bbe6f", x"bff0103bab3862ea", x"75bb5baa5160aefe", x"f11bc441b154fcfe", x"7478b8922fef0084", x"25b1cfeae37f62d5");
            when 22715249 => data <= (x"69cef0c454bae40c", x"1e00049422023cea", x"e6b9388482a86b2d", x"0afd1b2cd3831ddb", x"33d390712305ecda", x"7de22d9041f35b82", x"7b471638e7682c26", x"89c47a3a05725233");
            when 19503120 => data <= (x"17ea7806a199fae0", x"7a07bda9ce7b3fa8", x"ebbe314527b59d85", x"4bdde03c7a6f9016", x"d24de2bca80d2a66", x"04b1a824af01c987", x"54e0b5d368f185db", x"3c3958d35b0ef917");
            when 15693489 => data <= (x"fac2a88095a04ac5", x"504ab3091e0867a9", x"8b695498f2783c00", x"b173d33a9f577560", x"fc608a30bb77df06", x"fbd31643fb2630b4", x"dd7642815f7d0dd0", x"8785587e89cf2202");
            when 23533680 => data <= (x"7d659feb048cd16a", x"4449246fbe2e722d", x"8ebced987bf048b1", x"13774a2f4569f1b8", x"214bd7414a7cb436", x"7455f84e29d7c381", x"0f172d3b06af55ad", x"9ae98a5150648f63");
            when 21652210 => data <= (x"8ed731917197d032", x"7d24446609a03db8", x"ab589588db7f6e7a", x"fc387b93f928ac2d", x"1457f0044b162503", x"096c64133b433a3d", x"6abc58ffc6cd1746", x"47af981c9a917f10");
            when 33877335 => data <= (x"0f29baebdc930c61", x"0bb109ebfbd4f8b6", x"6f8f5a969dd777cb", x"1a181455a9ae61d4", x"7ff9c0bbae6ef48c", x"e94c8c44df4fa04f", x"58d23d170c028523", x"6d5b2e295e024ca5");
            when 2462096 => data <= (x"262d10bcf30738da", x"fb532276e0bc801a", x"56e252300d857142", x"51b96606ad944124", x"9a38ad4cef21503a", x"75d0cd90824e830e", x"288c2db2103836ac", x"f4cfe396d63de6e5");
            when 543925 => data <= (x"fa40e915331babd1", x"6845662a41170ea9", x"66f3d50c4c86a47e", x"a65eac41a67677ba", x"17f3639bba9ef5e7", x"9f8bcfe2f4644468", x"4145cea94cc91012", x"0038529612dd3001");
            when 14769308 => data <= (x"061f0c665830886e", x"bc3d0b073ee18a33", x"47ce365d405dcd2b", x"fd1823b11bef9f3f", x"906010663dfc8328", x"d840f9d79ff385fd", x"d5f261cee48c5f7c", x"3b2c570f13d3412c");
            when 2492450 => data <= (x"62805fd98c1ceb2c", x"2c0eaca660b9fe77", x"af6b122fe231e07a", x"b0d23c60e1f2cd50", x"9337a5c42ca4e05f", x"967594ec19cbf380", x"e803d2ce590606f2", x"f8456ef8f6c80f0a");
            when 4508936 => data <= (x"d01c92cacae12c31", x"8bacbf710260b2a1", x"faac36d839c8abc2", x"eff683756a742f76", x"c98672ec9ff6c31a", x"1220ea2df76e27f0", x"c59c0916782e45ea", x"e4792eae2b67fd62");
            when 10215154 => data <= (x"9d01879efc64be4b", x"c2c6fc36b8f3366e", x"bb5f14fb690bb4d5", x"fce2aabc04c6119c", x"0c3b865f50db8849", x"f04c521c7090b4ee", x"28eb654d9ab53fd4", x"106a3f4329c40aac");
            when 1551943 => data <= (x"5e3520d13f90e035", x"0952f0f2deaa3f37", x"5fafb2ae30074765", x"4d3c384f17cc00db", x"a107d54d817d22c1", x"960e534d09cfe583", x"ade2bbf654c952db", x"adce6a3f03b49233");
            when 30440060 => data <= (x"91d3e768cbea81ba", x"1eb3f7b7b92d0f4d", x"61d108737914d2ef", x"92e1b1dba191dcc5", x"08b008eca7306c93", x"a5cc515e9a0c8a21", x"ddf32af05d8cebc5", x"f41c80d6aba834fd");
            when 7083178 => data <= (x"8f4b13e2226a15ed", x"a85d1c2bdcc5c378", x"77e9e70118236662", x"57a4c6cf7254b85a", x"a15e031366c6fb99", x"9da1433e6e9cfbc7", x"dbc40b027d7ff1d6", x"a9086c4e1cb3dc48");
            when 8103932 => data <= (x"ea84945338b21b2f", x"d45e8fd77d533602", x"cf1755586cb8da0c", x"d234d584260cb169", x"ae944f1437d0c670", x"811761cc6e5e5505", x"3e448f449723e52f", x"025c535e6a405c92");
            when 21729716 => data <= (x"857c284f7e01c48b", x"ff786feb68155bb9", x"23c145baf1bdcde4", x"2691f922a41e6e43", x"afc25a300d260988", x"5f704f6f0451d88c", x"42a4b61ae089e8ca", x"605b3240f18661f2");
            when 2644013 => data <= (x"d888847e6fc49daa", x"0d9d5fbd93930ace", x"193c6a02b1b6b72c", x"58ebee6e8d530141", x"6d57bda074d7cea5", x"63cff271dab8cdaa", x"a81dffac1ee3212b", x"ce26f40b29d254d0");
            when 9527026 => data <= (x"7219eb3e61aa80b1", x"dd5f9b5e5eaa6067", x"eae7f156d015e47d", x"d3b36a34014f6c1e", x"a2f4d4b371e992ee", x"2d052e9603ee6695", x"d47b59736d807854", x"a343e53b9cc7253f");
            when 565775 => data <= (x"60d1a222d2841a0c", x"861bdcea0ff2fb4d", x"4cf21881fb38654e", x"dcd32f101eb973c9", x"f0f0be149eb30981", x"4ae4875287f9741f", x"5f56d29aac85a0a2", x"10507dac03b58d50");
            when 20324727 => data <= (x"17d698fd0a541cb9", x"f8bc54d966939295", x"4291479735f4bfdc", x"e5a3ff37a66a7c75", x"48d63aa02974d367", x"7a98d2b1ca180143", x"05051763e18b1617", x"c5140fee026332d4");
            when 5189323 => data <= (x"a26fbe7ee8287e25", x"009e8d70409ce72f", x"59a841f695a63843", x"283ffa5a58191aee", x"83667a071aeeb1fc", x"f83e977475ca7926", x"509ec2db95155d75", x"0f869fd5dea55f96");
            when 9174358 => data <= (x"e70a5479ce803e24", x"6b63380c2fb57b97", x"f41870dc031f7888", x"0ecda357bb2a3da7", x"f3e94ee34fad564e", x"231e16ac59e68f8a", x"340c351afff358e3", x"864cbcee0d04561c");
            when 11970497 => data <= (x"4249a49618eca73d", x"2a265f0f3de81e92", x"5351620447a0dc50", x"ac7bf07ad9d395e0", x"5ba7f137d096a649", x"ec4b36e8ef151508", x"d95ebd1a629a8fa0", x"58ab42d431e1475c");
            when 29751606 => data <= (x"06139a1179b89df1", x"f6c9d254d4a3e4c3", x"4537303ac1f106ef", x"e25fed5361259055", x"c07c21d714b34e27", x"5f92a12f42de1a0a", x"2aaa62ccb8633769", x"e329b9b5c4451a24");
            when 32388723 => data <= (x"2b1da7924ac2aba9", x"dd45f2cdeb1d7bda", x"d38567424254e607", x"02486961fde4824c", x"e9dbeb4f49138399", x"e5e25da74f6bf614", x"40716a66953d2af9", x"46d0e2d014469f11");
            when 25289195 => data <= (x"eb9c85fff87a4e8f", x"0a7b2797b431e89f", x"022e0474e2b0fd43", x"ea8cdc5c157f1aa1", x"6cdb91a4f7d634c7", x"5bdaa92bcd2873b8", x"129f13d0ea1d81b7", x"2b195c9dc41ed839");
            when 11022319 => data <= (x"0a4cc2e2e68f23c2", x"5a4aeb7ef6e4ca6f", x"c176bc41c0bb10ed", x"47925c80cec05d24", x"211f987d6e08b0c3", x"f8d66cc6e6ddcad9", x"da8ecd937b1b1180", x"741a17c32ee7b43b");
            when 26702632 => data <= (x"d390163a9a9723d6", x"93243ee4029c28ab", x"4b733989184f4370", x"c358dcfde382bbdc", x"a3ece4ce264c9cf5", x"69013882e2403c99", x"9b56505b56cef684", x"f55b74f611b4999f");
            when 23285093 => data <= (x"8b9283bc857a1f19", x"ec33e07063c610df", x"1f3045d3b8d6f6ac", x"bcf23970f3aea7f5", x"58e12abcfdd85bdd", x"9ce5d71dbe67de57", x"4ea7904796cf102c", x"171fc2047ba75ea1");
            when 30718509 => data <= (x"54bfabc68e3e6396", x"7f6134b0622ce2d0", x"e5066747b07cc896", x"994aad01aeacf329", x"9191f46931cfc654", x"758982a8a33ec5b6", x"dd5828b961b73048", x"cb0f4cec233c549b");
            when 25735852 => data <= (x"c8c2ce4656544d84", x"a629888148f5eeb3", x"305c9733145099ae", x"66022c99c93e0957", x"b806b9e3514a2357", x"822d3e3c3191b21b", x"f85f960de2761363", x"86e16427725b1c30");
            when 27714576 => data <= (x"3ee4883ae3fff2f4", x"d722edbc10d19b43", x"bdff139f239c1d9f", x"79ef7a7e67fe232f", x"c2a77bfe812db376", x"2006db01e5f1f995", x"66f332b7dd5874df", x"f2dad348d4d88ab2");
            when 32817403 => data <= (x"24d4c41db98318ee", x"c5e3466399c5da9e", x"9dabaa116a70d6e1", x"30dc668b27373ce8", x"370d981e3a735c4c", x"1624e67100e60c2f", x"5711c24ea9961202", x"de3433a8c07ed92d");
            when 20008746 => data <= (x"52f5f9b3ca7da24f", x"78ce507033f81b6a", x"cf5c966d8678c902", x"ee6b86ee385154f7", x"72872bd2239fb714", x"083b6dcd380f6ce2", x"40c7b9dc27b2d9b4", x"57d8b16c847cd676");
            when 28857918 => data <= (x"88158df9d3bc9d76", x"65a9bb30413bdb12", x"f3abd28dc54816a9", x"88f0bd421ec3bcc1", x"e50c9f0bc91d0105", x"06827633dae90e03", x"b66565939178a311", x"b7c712cee34de3e8");
            when 12177590 => data <= (x"3a4cdd2f547feafd", x"90bfdb61aa446b4d", x"0aa7bd0600361f77", x"4b0c6e09707578a9", x"38a315596124201b", x"d1bfb97a536396f8", x"2625757267857c4a", x"58718ab3ee05e1bb");
            when 18480009 => data <= (x"9718d9d81cebd4cb", x"f10874c0f2d389e5", x"ed2ffb1e8cc3aa00", x"81a9277c8555c518", x"0a95fbbb0057c9bf", x"34c520981c032825", x"f5e765d19b97411d", x"2782a7adb89168fb");
            when 26568246 => data <= (x"53266b89697e098f", x"9d9debeae05194db", x"bb3c5dbce0bc4b45", x"e9251140dd9e6754", x"a5304df45cbd4016", x"4526558c65d9835f", x"c9e97f873d12accf", x"71f76e651312e671");
            when 30328079 => data <= (x"ad2674c1a470a119", x"7283981c02e54c90", x"eb648b53a618e731", x"eb6dfa80ad92db44", x"bf7d548557a0c3b1", x"46a0485e1ce41153", x"670a9f2ce967429e", x"33ba551e01d8212f");
            when 22402446 => data <= (x"164bde36827eb809", x"0a199bcab23562ad", x"6c96210c4339da82", x"6a951291196fcfe9", x"73f749d1d61e3707", x"0b29669e4653b87f", x"8d1d3ab702470249", x"818325a441c56584");
            when 6582966 => data <= (x"8f2b7af265213112", x"18d917067aea5f25", x"27dbd80069e7f080", x"af88fc0f80c63c74", x"05cc2039e713c323", x"c4e88ecbd9d8a707", x"d61d30589ede46fe", x"541effb6b6892e9d");
            when 20566003 => data <= (x"c1ad66aeae198c14", x"ccec1f53501d995d", x"c02d8799c6ce16b8", x"01727001aa4a3c0a", x"5fbaf536f3ebfffc", x"24310cb2afefc22e", x"3aa991c60bbbf577", x"5d6c2860ab5a65d7");
            when 3584364 => data <= (x"2b08cdc002ae16a5", x"c8950f4827489015", x"1d38e88d2c454968", x"20017fa5b54f05c0", x"e8a3ede406f2e5dc", x"eb718a6a97291292", x"909ccc716ac16129", x"9e2f56f306389e7f");
            when 31948859 => data <= (x"0547b320dc25c7f5", x"9106ad38b07b7361", x"e266d765b3f34f32", x"25fe133089319f66", x"2cdadbf403666463", x"a7f20c5520ae8b78", x"66a5b53aabe852bb", x"d68f2ac6911b71a8");
            when 11293022 => data <= (x"e01342a0f25d6d86", x"cb4865f88d8a6667", x"4cfa042c94c6fe8c", x"315c47118cf26a41", x"bb67a3b94cf25f04", x"24f912fb0cc6889f", x"1e06ac3fac73a97f", x"e78a03138009dfcb");
            when 14777370 => data <= (x"ebb66ff1a8399edd", x"49fd5d5042a42e8e", x"102233ce77e51184", x"898d98cc4edae589", x"6c92ea0fc7191d04", x"edd6a6cff7082422", x"0b2f887a55954263", x"7754da22135e4bd6");
            when 17230199 => data <= (x"53d3f8f0bd474f15", x"e912e507b2f86e7b", x"e7ec2c8dc1199561", x"85d90b7ccd452fbc", x"0fac6e8fd4846c8f", x"4c9e720a6e622a77", x"dc19fdb5208f86e6", x"ed94a2c95d3ca37c");
            when 15072635 => data <= (x"4205aea6e85887c1", x"2266ed33f4f079d7", x"1608383b4bac651f", x"ee6f40f2a3e8e3a5", x"68f7d24a712bfe5e", x"e02588684123240f", x"1a09298ac026188d", x"b5ad6ea6b77051b1");
            when 26900664 => data <= (x"e2c586f29784aaaa", x"e0944760a7630e35", x"1a898b66944a27f4", x"0c5dbc30e6305e1b", x"b32f080aea49bd9c", x"a13aeee39947a4ce", x"5f4277dd229c7e75", x"7b8b9c4490e4b970");
            when 4756686 => data <= (x"220de69d69058caa", x"5236f7a5fc46fca5", x"e8aa242e59ba6434", x"c1770d596b51cf0f", x"2b6e1a5dcbd55a2b", x"5584f86109197b66", x"fbec90cf5f62e31f", x"626f3c11c7382c24");
            when 9595525 => data <= (x"074d560e3f33f557", x"be52b60e819b4dc9", x"8cec226bc562f5c8", x"a9b101df683874c4", x"2f3448facac8360a", x"4a6778a37d56ab49", x"3d2345eeeb5d7db0", x"9813ad2a787893b5");
            when 3535166 => data <= (x"12a16dd85a8a9535", x"dfd11c1edba02f30", x"da1b7f25950afded", x"9837775fbdced219", x"631cba0375919e57", x"90a9a706e4e76240", x"e40c5bde44da71d8", x"afbefd9a33ef39a8");
            when 9787308 => data <= (x"412d925dab128fc1", x"b4261eb7c62b6b2f", x"b3a9c7d092123d92", x"9487bc9cd8d92440", x"b246b11e6745d7a2", x"86482e6ef4e01018", x"0b21fa5690dbca4c", x"0ee35790250255d0");
            when 23572060 => data <= (x"1a403785d2e1b1c8", x"caef2ceda960b92b", x"7073ed6f446a529f", x"a7bfdf37a311763a", x"c56b47075a1144cf", x"b961a41e25d4d5d3", x"4acc24aa2c8ce9f4", x"67a04296f253d6e5");
            when 25293837 => data <= (x"e6e2ed951f0679ff", x"79c8bf07248ba872", x"b6d473fce0d386f5", x"59c0aadcd9223ba6", x"4bd23230c02f6153", x"3fc207248c5a921b", x"ed07198ba5b47af4", x"81b9a554112f0382");
            when 12902376 => data <= (x"af5ca885da5c8a7e", x"da96728b925acd3d", x"e08cf51f335644bf", x"72a011c206975080", x"f85d35181b6e7bd6", x"483b2bf17a217b33", x"97c30f9672436e23", x"8e15c13d4b5a3e36");
            when 32983705 => data <= (x"a425828b87cf9ed3", x"b248d43cef4ea43e", x"40c6f327dc9c5f69", x"ec084474f3819762", x"50ccb9b0ec233383", x"fd2b8346d3b75ba2", x"4d2394cf3559ca53", x"b97c99b3e4432637");
            when 21810654 => data <= (x"cd4f342dc8bd7925", x"095812bfa527630a", x"6de49e0f890e335f", x"4e81d320e0259705", x"c3e37a7d9023c0c2", x"7954daca3b2f7142", x"2f04732bb24c9e43", x"573232ce19848e10");
            when 8661507 => data <= (x"437a017fa28b5789", x"ae4086a9a4be6561", x"92a5c1d3a6e32ff1", x"65dab2a52e10a401", x"76464ab7da1963fd", x"59919ef91a8e3189", x"6a5de1b32c5a5868", x"dd33c9cae61f21ec");
            when 13389377 => data <= (x"abd213eed695da8e", x"74f1b56ced8be212", x"1d134e819f358f81", x"b9811c4cdb5dbcbd", x"27b5b8e6ba71da51", x"a60ba831b6355d5c", x"f1ff6069bc954db0", x"69208613680ca490");
            when 21841342 => data <= (x"488855494222db8e", x"372ddeeb0cdfd0e5", x"e11af0a302fcc1d6", x"d919f69b0e28ee2a", x"c66f28bb5eeebbda", x"171dd14fbc0b51d5", x"99054b6531780723", x"434cf3b1362856c5");
            when 6450793 => data <= (x"971b3320a7285a85", x"aaa0176550df10f7", x"f1eef41828417dd1", x"dd98bc4ccb36e648", x"88fa27e23dc9635a", x"4e8de12a3a7772cd", x"6240d3281a49e840", x"25f410074c2cb938");
            when 7937209 => data <= (x"23e6a36004377af0", x"857d81f61bc5d6d7", x"442ede6a58f006cf", x"0df7ec077fdb4cbe", x"b4f1d7cb7c99c859", x"31cedaf4c065903f", x"1a472bf2635940e8", x"8af029a7d4bc6ebf");
            when 25646424 => data <= (x"734a9d244da3dbaa", x"60e4f892b6d26f0c", x"702e771fef1c4229", x"e318afe06cbfb37f", x"3d133037a4b9b104", x"0f295e37d7b59c3c", x"9f7fd70b20098b61", x"43a117e1d6373ec9");
            when 25275657 => data <= (x"cd61543676208223", x"66734a464d1f7c3d", x"12dd717a8c797eda", x"34c5d086992f5c50", x"4f1a3472d6bfc9dc", x"c53689314b2d05d7", x"0f073af594b0ce69", x"5aaea909ac7b381d");
            when 3614345 => data <= (x"c4fbd223c7f182c0", x"532780462cd8b708", x"ece7136e275e49a6", x"133fdb2373daf510", x"e656c4f751fb9b57", x"4e5567c8110b7c72", x"df3d8e0d91ab80d8", x"b68b2f97b883452b");
            when 25334562 => data <= (x"402fd316dfd26619", x"04f430b751fe0f17", x"baa5b45bcf124cdb", x"a4f9f2d7bbdb39e7", x"cf182111a22cf12d", x"7488a8e66e55009f", x"038fb7824a2cb14e", x"3eeff7da5030366a");
            when 7549403 => data <= (x"f0865372409f12ab", x"bc10bfbdf07d529c", x"85e7a0bd3c6531ba", x"fae613af665b7ed3", x"d6397af1d8dc5412", x"96dbac04ca55983e", x"b98f3f167c97e323", x"88bda6b29953c7b1");
            when 4459798 => data <= (x"3aaf574a3d637957", x"1d68675dde8a9df0", x"26fa51f654657610", x"17802b6dfee7f1e8", x"b5b2bee83b136990", x"fc3d0fd256bab6d9", x"61b6b6d2a49692fd", x"309edd706226c3d1");
            when 13741604 => data <= (x"1ceab2c74e8b96cf", x"8bbdba775ed72cd5", x"17ac6a6617264bd3", x"daaa82f4d78e8c56", x"2745b9fb58845f1e", x"18e1efd1d8910fd8", x"1d9131b8fae88279", x"9600a68215fba14c");
            when 24094371 => data <= (x"7868afa8227b7b38", x"8f1eeab85d93bacd", x"6758d54cbe4ca3ad", x"adaf4eae2f1d5f59", x"dd3db3907a8c937b", x"b1b369e7bcf8d446", x"e6abf3ca48e34fc5", x"dfc3df6f8f6b49d2");
            when 14014360 => data <= (x"06fb5771ecaa08f3", x"0707a269112f7b89", x"6021cda386ff713f", x"d7cc3130d53db657", x"c75e7c8806b2f51b", x"b9dc45454f42b362", x"1358a29c655fc175", x"697e4d462ed8ed4e");
            when 31857536 => data <= (x"bee7de990b6edb66", x"d9ed4b2721f015ef", x"6edfce85bc96351d", x"969b91ec69fbd4be", x"e5999f51e12ace70", x"ee2dcabbef3f37d9", x"a7d498539cc19dde", x"e9e30b3e348ce405");
            when 4780629 => data <= (x"aebaff14f607bc48", x"5fd93b7e0d8a6c5c", x"520733ac80eafe7b", x"8f196f8953bc1847", x"b53e76c94f9f29d4", x"f57c4854513df3dc", x"4cf4d52365fa5473", x"1ffea33c42f76480");
            when 30161895 => data <= (x"dab6441201dc4829", x"2ada50fa8cc21a95", x"85eeaf9e341f8701", x"f94bf618dcfa55fe", x"f9943ac62adfe3a8", x"ee0c98d18023f1d1", x"4e05448955f42b1f", x"5fe0392b49eaf091");
            when 3829498 => data <= (x"3c4fe4afbd4b51f1", x"c76dbec51dfe0698", x"f4bdd8a62c4b6f4c", x"cc645994ad6521f5", x"8bec73e6483dd99b", x"95e0c95ed82636a6", x"e9665519e234552b", x"40b6535fa2a9d5eb");
            when 2295636 => data <= (x"eafaa632a2416082", x"69995bd97d3c5888", x"940d94bccbd4b1a3", x"ccce8b8c9ddb0923", x"fa24ed99685408f5", x"6dda2e8ed4d11244", x"f94950d34406a93e", x"7639cbe95d43c1db");
            when 5258448 => data <= (x"9d5fb7eeaf42a67d", x"3534f0165048e213", x"02bf9c5ce6e2304c", x"8883e8a561155996", x"a78eb08b1eefc404", x"bbe0a1407b2403c5", x"dae9f661902840df", x"c7cab0e70d1e2351");
            when 26933705 => data <= (x"70c32098ad66e1ab", x"48d75aa53bdc0bf3", x"3b3a6598b9b869ed", x"462404733c06e6c7", x"9a10e8f46c486ffe", x"c02f8f540557c78e", x"2808a558ea018beb", x"bdba0d4edb68a402");
            when 10734475 => data <= (x"00cb197b9508be5f", x"fb7ba2aebd7f38ef", x"97cd116b09131329", x"8b759908b9bdf0cf", x"7db6d222628703d0", x"588050da32d0fb2e", x"3bc983dcdac2344a", x"da346db42cdff0db");
            when 7738227 => data <= (x"1754be3e1f539144", x"a8d0ec947af4bf51", x"fff40f39221ca412", x"f7de30e1d3c92e70", x"295a7e3b9cb21a4f", x"f711f55a9bdb441b", x"e82ad382af3e330d", x"04aa63f0966a8e6a");
            when 27644161 => data <= (x"b610d2e588edf51a", x"c0570cd02ac87a6f", x"94267d308ae3477a", x"3f3ecbda4ef10c15", x"d377acc4808cd8fb", x"d75a29c148f8ccd0", x"e6de30b10f415bca", x"b737da1733f48a0b");
            when 27566367 => data <= (x"4dce26df45011ca0", x"de75353445e90772", x"a1fbbd8567abce1f", x"f3bbdd80e2997dc4", x"25d13e97ec2918f7", x"259a15879310cabd", x"2123ae80e8554b24", x"da12ee619eb147f7");
            when 17697909 => data <= (x"3975f34524f698d9", x"c893066efedf56b6", x"600183274ca16f9a", x"715d03a0b757408b", x"b6eda3c87fda2748", x"21eb548d4a8f8ba0", x"735d41c0531521b6", x"e52e36ba04117923");
            when 15078454 => data <= (x"c9ae246325318d41", x"d374c4c168cc4885", x"9c77e49499b54813", x"92cde6560a2a1348", x"bd495ff0eb1c3170", x"c7a9b75fbee6099a", x"29b0d5015d756d33", x"cfdb98ed59ed063a");
            when 18494514 => data <= (x"9472f6b16a8d2914", x"8e41c3ac3bf6de58", x"84fdd98023606212", x"fba72aac926953f6", x"b1c2090252be9ccf", x"f7fe3d200e30b928", x"c51c0480ab37ae65", x"582efa5bd0f3e649");
            when 29768918 => data <= (x"e5478fea89da4a21", x"3569f05965b79388", x"555b37534806af97", x"206e2e0c6be1e834", x"fe78ff9023f4a689", x"2093dbbccd93cdc7", x"6d05b9428ae5997e", x"95619e748dce7323");
            when 33711137 => data <= (x"120bf05d3cc2366b", x"b2e7d3b008c508b5", x"ff8a700ef165dd76", x"ff8cc6fe425dce11", x"f6886744e9e9452b", x"c8aace1fac1c8761", x"4197a693d8caae1a", x"38ca5fa57049a331");
            when 13322072 => data <= (x"391d03b5458b38a1", x"5e9061fe399497cc", x"d52060718dbb3a85", x"4fdd713046bee259", x"e9e5e92c078c2387", x"accfe5abb98f4eca", x"50beda6fba2222ae", x"497997d254cd3ae9");
            when 18593504 => data <= (x"8d657a9d42e82827", x"833c25a4ef2a00cc", x"9a868b24a22e620b", x"9c05f5f5de3872e8", x"7f0be8ddb978ceb1", x"dbd123d28a67a0d5", x"c7c0d1e20f296dd7", x"b1fa4ba5fb17e4ec");
            when 6833327 => data <= (x"03654ef293466e1e", x"1df4e8431414c4f7", x"d1cb04a5a99023dd", x"8fa0840fc6c23c89", x"b38dbcfef8e4a519", x"bdf7d5728cd04c85", x"e9e1664d30992d1e", x"6f051cc983cfbb75");
            when 15732529 => data <= (x"26e3170faa405949", x"47ae08646bcf2613", x"1ead7e5d78185f55", x"09ce61cc35c4a9ff", x"1735c6164aa55323", x"cee85aa35445a10a", x"5f1a436d332b141c", x"4d348676bc6d0d94");
            when 2350290 => data <= (x"45fa95297c8e63ea", x"ed02a50e1ecb2408", x"d8dbaa338d37a0f2", x"aa31f35def352c62", x"8257dfffa4b12895", x"28100f987293df60", x"92e7914c5ea593bc", x"04bad7702959c31a");
            when 30947154 => data <= (x"b16d1b1b0362a5a1", x"fa1b27beb68aafa7", x"71cdf0680d75d4f0", x"1e2fe59e9a154e75", x"edd607511554f83b", x"0cfbc040b4541c79", x"1c0623eff9880347", x"73a23bb9e56a294b");
            when 19868265 => data <= (x"e798b104f2c20eb8", x"659801b0d4947fa7", x"144dbf715fb23452", x"d51d031aa6520a63", x"f5431e6af537a709", x"639787aa2bbd3895", x"7a432ebf6ce75658", x"585abc5d056793b8");
            when 10548654 => data <= (x"f09c1f6745e5392e", x"ae29d8b0bdc7ecc8", x"a565d94af0bdd4b2", x"44602925fe9b8bf6", x"55be94698149475f", x"7ed380f19b8eea70", x"e681a693427ea1ac", x"fe345d79b351b3bb");
            when 633282 => data <= (x"0552a87aa63831ef", x"b00c81c249eefc99", x"23de9b147500fe23", x"2d04c4a1c1eaac29", x"0108b3d130da230a", x"9acda7f563961cdb", x"a5b1835000febe24", x"827f3a3249e8140f");
            when 14764348 => data <= (x"6b80419070c452f4", x"aff844f7ab15e89d", x"fbcc1640c7eafc23", x"3e498c4d9e0b7cdd", x"a7cef3468834f497", x"4f4c6317805e321e", x"5083ae638fe1dac0", x"1423484e2168c751");
            when 16118515 => data <= (x"0d43e75012c8ebb2", x"5001ff2e0a7942e4", x"41a681b907affa80", x"5f49e83933b8a12f", x"6fe2f930a84eb5a0", x"42d6e90a451164e2", x"d965e7595a942dc2", x"f9b8ce11bc7c6fd6");
            when 20506190 => data <= (x"691b4abde689905e", x"5844f85eff9c59ef", x"04d841a593bb5631", x"0adbe08664e90c52", x"a4a960b9aab8e274", x"f27fb2f8e6fd614b", x"461daf31e8cd58c1", x"5785be76cb474d66");
            when 8762812 => data <= (x"6ea26fb5d98a1fe9", x"62f40c9389f61114", x"de5e72b61a6b8a18", x"0529f9043d509604", x"516c4946af450cbf", x"9161a636062ff2f6", x"f3be7abe4f4ae6e0", x"c97a530c866e9ace");
            when 11567115 => data <= (x"3a0e70ededdd24e0", x"8131c65a4aabc959", x"9601600f9c84b746", x"2aec0bf51575f8f0", x"9c1ca062ef8a7739", x"a34d732bdbbf882d", x"2a558834d9087180", x"cf34f90d80217e54");
            when 3775082 => data <= (x"04be23954487f0c8", x"079b29c68a6818fa", x"0423f58e1eee632a", x"92d2cdab5b123806", x"3ac2201e1ed24155", x"5c2d9f15755e47a8", x"596a6eb3d866ec98", x"a4827f1f4e005ea7");
            when 29348073 => data <= (x"7b8b541ab56796de", x"d4b091f356c7f770", x"538893a7e33d1346", x"0767b6afa67b318e", x"9b5f3b84718c52d1", x"10f560546c59fe6e", x"c9833511bd47b603", x"4031ccd45b4a843b");
            when 8854555 => data <= (x"0466a8a4c5885101", x"22de33c4151fce7e", x"84a36cfb1b39ed6d", x"60944e6e35f03a95", x"960b54eea881b1b6", x"3a4bbfa1433272f0", x"2684e8c877699cf0", x"5b16af93c4a11f46");
            when 11658878 => data <= (x"77993f0f5a09502a", x"ae04bba897a6ea8e", x"a0064b2bf127ed34", x"aaa63a84277046fb", x"22a651e4997a5124", x"33735191047df033", x"0a58e6245e440be1", x"7a569e5b2f4cb401");
            when 28057673 => data <= (x"cfce10a239c5cb89", x"48a46710e7445b91", x"6f9fda2c1a62481a", x"1cb1f4a927439e61", x"b600acd682ee6706", x"c0e70e1fa1805c8d", x"93d8d016591b56b0", x"3d8927e0dfb2922e");
            when 26347337 => data <= (x"cd416620bb44849f", x"b2c364a144217e78", x"1dd6ff7fe2febc2e", x"5d026c02a39f4072", x"23f8469eb170f5e7", x"016ad24c77ebe547", x"315b091b80b52aa2", x"621a72b8264e7c94");
            when 26433785 => data <= (x"a5c08841fe9bc575", x"08bb7bd6cd5cd992", x"d19214a4d37783c6", x"ac3c0c6464e4d992", x"2e59428bbf50b13d", x"1f77b0b781830c6a", x"42a9d989ad8fdd86", x"a7181f8c7a5d83a9");
            when 13078318 => data <= (x"5d619160c3e529c9", x"fb23733b7f26919f", x"699073328805f043", x"5a16a3fdf689c60d", x"3d53a885eff5b45d", x"efa8ed484d2f3429", x"b1016e5969229cf9", x"f5411c1b206660bc");
            when 22423084 => data <= (x"9125db52a229418a", x"40e5cb25d9279e7a", x"9eb4173066cfcfe5", x"8a00ea401a25272b", x"f9ad3c2f030cc02b", x"2be328085c0d8113", x"d8f4162ceda84f53", x"518f6e4624283d56");
            when 32641538 => data <= (x"48d12d9c51497a4a", x"bd3e64fc83817b20", x"6b9d0bf239f2c6b4", x"fb97f14adca81a34", x"5619819f0261736c", x"055e870300285f9c", x"37ad3aad5baf6832", x"1e0f6be3ddc39c16");
            when 10900986 => data <= (x"811a0cc02dffa842", x"a761b8ff77cdd9cc", x"7544f1911955147b", x"0a0c7ed21d5d985a", x"098f126c23426d7d", x"adabbaaf2a83f34c", x"1ce9402ae3f007ef", x"65999c261683608c");
            when 9939252 => data <= (x"e9e678446498a015", x"98c1b66ec4453476", x"85f30f5c01887b45", x"ef59cd1f1cc67d35", x"a66c509a6b1a76b1", x"bb4b8aa0f6fd1104", x"1f6418a5d0c329a1", x"cecdbf421e9b7a39");
            when 31699199 => data <= (x"05adbeceecb657d2", x"08722510be5ea24b", x"75bc036f9a1f09ca", x"47b8b493c60649c8", x"0487486972d638bd", x"0f87aff33c40ea35", x"203e5d3a60a82e8b", x"a25d3885b9e8a6a7");
            when 14905002 => data <= (x"21d4c741d1481189", x"4e37172d4723658a", x"ce8bedb691055fd4", x"ff82323d77f1c071", x"3d4b8928edaf9628", x"60aba58bd076c06d", x"54e4e9f1e4750db0", x"71c069048c4c6cb9");
            when 3888617 => data <= (x"d235db9f5635d2ea", x"4223046de77a0e8a", x"fac9a67f286d9fb3", x"a57f5b23d85a9fb4", x"476dcaaca3379974", x"2a85236639f4e370", x"3865b6d5c344ea12", x"91b0f1d25737a759");
            when 10492461 => data <= (x"1ce8e6ed9326cb03", x"8732b39bb1ac94b8", x"8cd0cfdaf410e5b3", x"3f73676a2f0a6e2b", x"139abf468af7418d", x"e367662e6bbacea6", x"7d23aa814ed4c82d", x"318177ec2f13cbb1");
            when 8796613 => data <= (x"d1cc9bb03f66ee74", x"831ae04b3b7a666c", x"98564bea5bd7c4bc", x"6ac516e7016fd83d", x"3dd5697a6df752e1", x"ef9b175f6a807074", x"aacfe825ae36b5cd", x"ae20ac22ae900d39");
            when 19707977 => data <= (x"c5e97419506f659e", x"2a0077a3faaa5b70", x"1e3dc20b7d91ec39", x"7bb2f4472caafd8c", x"32cee790eb5b7f01", x"2874c2a5a2ee728a", x"4a899512f8651439", x"a494787101b1f766");
            when 2663771 => data <= (x"86292802a88ba7e1", x"5f0091092b476aab", x"c682cde85d4e8aff", x"7d7d3cb826cc06f3", x"9c0c62593e76a16e", x"d78cdf813e24cca2", x"72110a54ac7fc280", x"111a4c4e4182b57a");
            when 7392881 => data <= (x"f07829eff133fd69", x"08db5ccdd10fe2f9", x"146b85c1a0fce8cc", x"cb1a44670ca17336", x"d87689b232ca74cc", x"b0061c759e92700e", x"8a5f25e6201e5d5c", x"8b13ff155faa45a2");
            when 13679357 => data <= (x"1feba05acaf283b1", x"565e27a0349db455", x"ec7b749a181aa2b5", x"25fe2300c3a7ab42", x"73ef121215360a59", x"1b75b3fa484b66b1", x"9148c25ef397eeb8", x"e4c8449b078f2c82");
            when 13829041 => data <= (x"26f16796db7386dd", x"4f9d6bcf922daaf3", x"db3e4ef15da63475", x"91e6f58354541e3e", x"60af3285164ff757", x"701568a084382d03", x"8a76a6fb580d388d", x"a85568df5b5c89ea");
            when 8063796 => data <= (x"40b792767a9609b3", x"ac9ede40c0d211e3", x"dd2ef26067e2154f", x"2e474dacab743e97", x"f02142b5293cac64", x"f9cec7dda7e4cc59", x"96069cb88b2de569", x"97a5011c1bd793e1");
            when 29455316 => data <= (x"cf8d35f1301276da", x"9f3521244e03301b", x"94344fb448d3d1a9", x"280f9d1e3a0c7632", x"3e440911147f7f0a", x"542cf9db43aa3de3", x"54cb3453fc93dfa7", x"2de1c27c089cbb81");
            when 12817024 => data <= (x"119237d46ff88f8d", x"93b875c8da3d1c22", x"95f12b8ec5c82fb3", x"5009b6ba2cd1639f", x"219c75fc8adb4d90", x"879577062be8016c", x"01123df3ab5ff8fc", x"c3b2dcc49ec5e4d9");
            when 8381468 => data <= (x"0c7861c882d28e1b", x"c3d962200fd31bc5", x"e28aeea5a3e3ddb6", x"3c65583a35623fed", x"06cd74283348abbb", x"f88007f0dc238f3a", x"5f15433ab11ddc63", x"761f460b9dc65f7c");
            when 8463184 => data <= (x"49bc6705fcdd3f69", x"9c167b4fced50ff7", x"5ac74247d32f263e", x"6ac672b95a6482ff", x"2288bccf47c6c396", x"0940c89acbbc8121", x"360db781987bdd09", x"37b8ed79859639fe");
            when 12032992 => data <= (x"9590c4cb6df1a781", x"f90b7511a84bea0e", x"adbeb8d9dc443117", x"93dbf98d9103caef", x"14a4660ac5b4817c", x"35ff238861200430", x"1236fd497031456b", x"4ab88a8d711f77c1");
            when 19396319 => data <= (x"6cf720b56f0721f4", x"9219afd08bac6c1b", x"31ad6aadf89e187b", x"4a7c71074651c1e0", x"6a669d7d5a49296e", x"5a9ab9ed1186a731", x"ad0ecff24df3e41b", x"b812650ae3532acc");
            when 32978289 => data <= (x"25e33bd805016ea0", x"afa76a81b93f90c1", x"ecb19b6bc59cfca7", x"3bf349732edae0ea", x"838c1fcfec3c74cd", x"640a012e6fbe65ff", x"b3de185e6a016b81", x"9346d1dba4175dc9");
            when 11469312 => data <= (x"833ff7698352bd97", x"5508936dbc0bad1b", x"a71a8ed0b7437368", x"1fff4c7350434522", x"4c5559fd07a1e9ee", x"e69bd2c7623f7620", x"b7ece5a68658aff9", x"a2a1a525fbdf7a0a");
            when 18361884 => data <= (x"76a03fcb737acf7b", x"5d6938b1e5d25ad8", x"52167561b0c5462b", x"9bc57948a8e9fbc6", x"b9eaa3b1de6e1610", x"2544ee653775af5a", x"5d7d7192977be132", x"9ff7feeab35a9f61");
            when 4365854 => data <= (x"fd4f7c424d6d397d", x"fd5fbf58551c4636", x"bd579871005a4d9b", x"0159571081873e9f", x"a0690cb2f63fa6fd", x"dc76a5c71cd07e9d", x"1aa865711376a2d0", x"06494dde0d18896a");
            when 10394846 => data <= (x"9571ea4a03a5628c", x"745a47aed4fffcdf", x"2613f5cde3a37cc3", x"e54a55e761aba477", x"5e9a802bf8dcf867", x"4cf6585d898d717c", x"f8340b176b0b1ffe", x"855ede425718d3f8");
            when 32740284 => data <= (x"a31c8b700c873b5e", x"b46512b7fb8f26b2", x"6b0de009ce9dc346", x"52e1ade8a62d39a7", x"dbc048fa5cdc1dae", x"64e25cd956c8f8bd", x"33ed359f663f3fa1", x"9a52c8a43716ee03");
            when 31700698 => data <= (x"5b8eeedcaf19f804", x"4cfc8fdc2c7a5e2b", x"ca5f21fb15313cec", x"fd8a7de5c5a4ec40", x"8106ad693039a468", x"7cef02f3c227d6fe", x"bf9c5bcedb56bf82", x"d96924949233036c");
            when 9963594 => data <= (x"b0bf68c702146a7e", x"e8aa3f2f6e032211", x"c2faba3138a64468", x"a6037eccfbbc50cf", x"1a2fd348bc719358", x"e11333aad2dea1a2", x"e81d30de68a9c810", x"4191e7e0e20aebe8");
            when 4176560 => data <= (x"460ae64b461ff85f", x"614c7a43e714a466", x"9537f4a2dd1ef158", x"4074ced4d9dc0eea", x"ce41b2e6d1dfff36", x"9ee6ae53271b4284", x"7a29add77d33d80b", x"0a1b4d5490f23a2f");
            when 22983590 => data <= (x"b61627a40f91f8db", x"b4e8e0965cdc1ec8", x"c1466d94f3337830", x"845926f9181fcfcf", x"8a1f837163add4ba", x"225f84aec4409398", x"c74e9cb1ef093ef9", x"c9a5f593f6aaeee2");
            when 12890645 => data <= (x"7e2c2c7e6a94770f", x"646e96c43ad6b6b4", x"72a0fc0d0ae3ed9a", x"5f924a83c8788e0c", x"b9e5258a33f73508", x"21423a12f5c98ffe", x"02253f9564c59444", x"346e1fcb2b71f157");
            when 24381112 => data <= (x"78b5b3bd1fb87c7b", x"24e3068b3a926969", x"2068f6a326dbbae3", x"a79d124e34438a0c", x"6c388c2632510ae2", x"c46decc7d3aaef7c", x"edf83c1d255aa7eb", x"cb5189dd9e47526a");
            when 5264707 => data <= (x"882377362d9f05f5", x"0568ebcd605d3ba9", x"08769792623e9b6c", x"68c7bc6d860a8483", x"050923f37d1b104e", x"44605851fd1b3eaf", x"cc7a72820178060a", x"271455dac154d432");
            when 4975561 => data <= (x"1448f605767637b4", x"5a7e014179bf5d80", x"52317817845f58ee", x"732dd0b1015b03c9", x"f140c5c7aa9918cd", x"f2407ef2e230cd78", x"24dd3e66480c9025", x"80c4f52fc701fc69");
            when 33181049 => data <= (x"dc9ddf677c8c32ed", x"8a09a231cd821267", x"670ee56706cc8166", x"3616896139ddb672", x"e9b0de7c38668b7d", x"d1d785f8b39335fe", x"20b60b4b5850fa07", x"544011402587e140");
            when 1819364 => data <= (x"63ddf4b6eb79633c", x"bf0b0de484a06b98", x"496566c9600b1cb9", x"7ec583ab5cd64f1a", x"e46d07b1b7814420", x"4a9f22f14b674641", x"cdea764de92ea140", x"041cd09942f5a65f");
            when 13536788 => data <= (x"3a267e89826bc6e6", x"be741b9a427838ae", x"e752976f22fb79f5", x"9c1bccb2111848e0", x"88e38cc5506c71d5", x"2b621eda1594b9c4", x"4bc890d5aef12d2f", x"3e4e13e349b0793c");
            when 24143272 => data <= (x"9d046e6a437b4b2b", x"a723f7b1242899c5", x"ccd30950eb78acb3", x"c52bab6ca9398bd8", x"03b860a5d136988a", x"02e4ea62c78cb2b7", x"b3f8cf31e6ffe354", x"ab2245809c344fd5");
            when 8673407 => data <= (x"50737930374fedce", x"d131f82d524041c7", x"24a37de957150d15", x"2047ee63f4953b2d", x"7994c5076f430713", x"a5da5e670751c42e", x"5c67b395a5e1d420", x"1802302e21e2345a");
            when 29659559 => data <= (x"d5a8b8c9671729be", x"c0dac0618bc5ef30", x"896e388060d853c9", x"0436a17f2f39ccc8", x"7daeda1b7fcb1fe7", x"256591d32e57e072", x"2d828d15959699e8", x"472ff74cf95a7a38");
            when 16809546 => data <= (x"c7d0fc06caf4bd53", x"0b0be2af138db1b1", x"2353d15cb190ea35", x"632a34148a1ca475", x"7e7b0ebd8a24d28b", x"a77fcd653d712fd4", x"270f705b137d4bd4", x"2accf19188137978");
            when 24611897 => data <= (x"1b3fa4e000bdc6ee", x"47a589c34344c94d", x"0b558dbcb49c3e9b", x"90f5df770ab8460c", x"dfc5612259fccabe", x"b58fa1c5d4ad12d1", x"914d08c4dfcbf165", x"44ffd9ee4af5b8e4");
            when 32153863 => data <= (x"4ea18d58c7011293", x"5834db3b95b682a2", x"29f2553a870475a0", x"cd59ae3dcf854d7b", x"14597a102dfa0afc", x"f3e95fdbda48e3e6", x"96580ecdfb0c5c3f", x"1897092d4b762efa");
            when 30356675 => data <= (x"a4f8ca285ffea4f8", x"9b79a318a0ef1807", x"91d637ced1cbbc7a", x"54208f15c6e07685", x"f1ecdba7309f67c5", x"09e8889b01841248", x"9d3ad424d14c58de", x"790349745a53f811");
            when 30059192 => data <= (x"46510b4af6bc7d41", x"f810a8902472e7de", x"6006022e9f014cd0", x"01fee3d8a1c212cf", x"82ef35b1ac85c39d", x"67d72ebb737637f2", x"b4289e80bf582126", x"ab3da3271748bba3");
            when 6812502 => data <= (x"a274d48e6287c521", x"d2ec58ebd74bad07", x"a7782f67a3c99700", x"acf5798cbe4f8161", x"f672ca8700066fb5", x"ec2fdfde4b87ec35", x"93f7b723cda082f6", x"602023f5280c103a");
            when 17746076 => data <= (x"9785f15b91029647", x"98421c23c51be4aa", x"a501d6d3c849e5fa", x"a4d186673384ae9b", x"5382239f0fecf519", x"1c99cf896f39fd3b", x"853216e60fb057df", x"dbc18c84e6d2ca97");
            when 17444671 => data <= (x"14cf5cbd5c8c52da", x"4cd497d18e9a80d7", x"d97d32239a73df26", x"69a7a8addfe0da4c", x"84a4b2301157c9c1", x"8667f001575fa86b", x"21adf4c36a1d3c38", x"b8e64bc38b61ca7b");
            when 6591876 => data <= (x"a297a933ac49e18a", x"83136a10195a1ef8", x"0ff466c280ecf987", x"3e224347a6c046c3", x"9b70eaab4a680605", x"bf74811e91fd7b5f", x"c513271a6be6942d", x"71ec7edf14a936fe");
            when 33946871 => data <= (x"6a75c38bdfec6eec", x"4506fa9a69d7bf4c", x"fc08964d4d9a7d35", x"12b4f439a08d9f5a", x"7c36b12211062262", x"05e74e169a974fa9", x"1394f2ff6f861cb9", x"d9bf5cf5f428cc96");
            when 13274643 => data <= (x"f4a497b2a25e3993", x"0e9a6de1e993f9c6", x"ddf7f82626dad432", x"9e73211ae1e560e1", x"473d3a10179b04ef", x"81681fbdbecc9b17", x"557c286c522d786e", x"fa338fe8cdcdea06");
            when 2691947 => data <= (x"9ae8ecd0b242e434", x"13e825b20c3a1ae0", x"a0312d29d55175be", x"a61e2bf92b8f1f1f", x"cd527a520a9625c9", x"e18a16f89609430b", x"4615c3fc926432a9", x"e3bec05e932ec97c");
            when 15433938 => data <= (x"3db04da44a519a4f", x"7c5f9a6deb004274", x"7d804b48014aac3c", x"69c606b4198be669", x"19b9029e323a6df9", x"9a0f63ecd1185cab", x"d434a910fef8f296", x"0a8f1eded478b278");
            when 16449483 => data <= (x"74849da13071921a", x"e6385c0428ced3ce", x"c5bcca6a02e5952f", x"85071c016ded7ca3", x"209ecdd85e465842", x"d3d644e10e6414b4", x"13ae6eb083115856", x"fb223bf716d091c0");
            when 3013462 => data <= (x"31ceaff74367f365", x"68ee4412c532ee77", x"656c1e05004f896a", x"50e2ecf7905de1dc", x"156268627a2e568c", x"1fabd54eb5cf18b6", x"7f146762901fd7f6", x"2c6d81b68250c952");
            when 7748195 => data <= (x"fcd903d23b47a050", x"eaa97ba29a593ada", x"20a8ec34c0281306", x"7f0bb87afbd5d724", x"21c608ccf3e0429a", x"e50f852a2f3d0aba", x"39c388461171fe19", x"41284b48d2e75cd9");
            when 3543746 => data <= (x"7bbf2d7987688d4a", x"002279be392ea4bb", x"5d63ddfc23b57a89", x"1f4172151a7905c5", x"dee09c74c2ee0d58", x"cd441b0006ff8e43", x"5175b8d661c369eb", x"add0ec449106dc42");
            when 24869961 => data <= (x"91ae770c4cbbff8a", x"c6b6460b1fbe54d7", x"0e10f9ead96af566", x"90bcb1baf8da9576", x"4d2e0e7eab0be730", x"e3b19ec416936f97", x"1e89d73f15c9b3ba", x"8ecf9049d3175d7a");
            when 11949174 => data <= (x"b7049ee9d62981ac", x"842e8c207e48207f", x"9f6682302212d41c", x"19e100bf870c69bf", x"59ebdd8808aa81b3", x"3db57a3900f378f8", x"a67b27066eea71e4", x"31f5d4e7d45c4ae3");
            when 22402870 => data <= (x"c498e12424952315", x"a829d19b8bff1d44", x"775c0b81db0d6475", x"3821246d0abfc011", x"50ddc1d8e307c78f", x"25c6b139a2dc9d08", x"afb8e50f90ffdd53", x"b88f3f5d165dfbcd");
            when 22310726 => data <= (x"e5c9a0f1624513bf", x"7a97d712f95ea296", x"b197d80e5f53c5f6", x"b2a4f35d87ff6513", x"87d862d288abbd7c", x"2a95532164beaf81", x"1bae6d8485b389fa", x"d6bb06f99e7e1716");
            when 7359456 => data <= (x"835b80ad307d68c6", x"58ba67da499e6f3b", x"d95374c018d392f8", x"adc8c233ce8fda9b", x"ba3fe1cb27cc0c76", x"e9fb52728955d909", x"42b178419d15f006", x"8be6fa0a5db35c72");
            when 28544209 => data <= (x"9a77ee9a718d914a", x"ea0a7e7106078fe6", x"de54ffbfa08c4166", x"2ef06ec5e4388b0c", x"db16e2a0ce49d849", x"be69fc30e4d2a741", x"bf004ce9b7ddd51c", x"43011c0c1455175e");
            when 27952688 => data <= (x"64f741d51251f99b", x"c0e3522dd9c5ec9b", x"6d0fba41ff9543b1", x"50db7fe6a56620c7", x"363f77a06b20dc88", x"3942714e3d02fd93", x"3b07b34b677ff672", x"fcc5993c2bca0419");
            when 29584682 => data <= (x"7694f6e6d491891a", x"5309e235b2612dd5", x"38dbdc04bc284861", x"9e6db06765308e80", x"e2be9f0babf5f60d", x"027e4ceaeac6725f", x"88541f03d316616f", x"1e8bc217c67dfa89");
            when 31771485 => data <= (x"c583757182bb2f44", x"d6e4407bd1d13be3", x"d2114fe4ba590c98", x"093edddb848f0fd5", x"fe1d2e4a10815964", x"9620c8bef3c1be2a", x"336c5db8a7dccd6c", x"cea84d6a43578639");
            when 15813605 => data <= (x"7aceeca50fdccd6d", x"6b4e0cfeee4e6af2", x"b4b9bd4cf38a362a", x"8c5e0234b05a8ddf", x"483def1f693c72d1", x"56479fb357b86746", x"1fccd5119f3e0b22", x"1f9453dec0c3d56b");
            when 2761049 => data <= (x"1c65abaf9cef13c0", x"76aaa721ec97194d", x"bd2d1535482861e1", x"4fb4fcc7dd98dc77", x"3bb648bca08d9bf7", x"0e00c227aedf3714", x"6fffd740359f22fb", x"344fddf244cff8da");
            when 26437909 => data <= (x"a27760b678e38c7e", x"44635b1d910be0b5", x"b0f74d052c2552e2", x"ec70b5b633f440ce", x"f715f10f705536dc", x"82f3b1e25a0b3f89", x"b4d2ed1e5d7d9061", x"30e60103f38f3a6d");
            when 18454912 => data <= (x"59613e14dc9a8ddc", x"fa241d9358412555", x"46c0bb430d9f2e1c", x"e14b74d5c0102221", x"253805d4efb5d787", x"b58ed77a19d6d54b", x"903183a0c23a4fad", x"755435aca742b93e");
            when 32324595 => data <= (x"c3d5eaa7e7cddc00", x"e12c29f91dfdb270", x"5e7b045751d3f975", x"f74b7971833d5d1d", x"0b11cf5c6e2d18d4", x"59133b53a325d622", x"8de6fb92ae1608d0", x"0c38fe57c7088e60");
            when 19727099 => data <= (x"ac20fb6c7b47c045", x"1329509b4330e59f", x"c3ae418261adfd91", x"4b70382c7ba984c8", x"d1492a54006685d7", x"3cde2775cf809579", x"81f59bc835a1344b", x"b6ca60f1ea2a5a6f");
            when 13075891 => data <= (x"2cd49004d8eb57c5", x"8b95bfaf90966d06", x"c54a5a9f0f26be40", x"0aaa6866e568be7c", x"c95793cdda049f63", x"722f41121613c391", x"c668196f13bf27e6", x"f8e2a238c214ca19");
            when 25698531 => data <= (x"b9d0af158de35703", x"89a39957905ffa7d", x"05b7e6d7ea4c43b8", x"b46108ddcb838a46", x"5faa6d45f9a20b2e", x"6274efb9731a5b2d", x"2ec4011740b2e7d5", x"7d139e1d81692a71");
            when 28520775 => data <= (x"9c667500ccba9518", x"5c7e2e292099203a", x"2af08ea9e6c72e69", x"ceecfcfd28484970", x"7543e88a2da4412b", x"6be8f4e283e3e15d", x"e35b2d374aec9dc7", x"aa59ea8dc1557a34");
            when 27384836 => data <= (x"7b5565b1fc082273", x"ae07ff8aa16ea7f6", x"8672f9e4a12b44d8", x"01c94ca4adf3a505", x"2dcfa32e6cc63f9e", x"a1d5d03f3f930eb4", x"5dabb8aa0f02596e", x"952b85e2f13a97b2");
            when 30928118 => data <= (x"1909ca8ad380709a", x"e548da63df303e7a", x"22b05cdaabad93e6", x"6c851550068e12aa", x"5fc01f4e1cfbdab5", x"e52cf60db480ae8e", x"18c38d248ce60a59", x"08d23f8aba314a10");
            when 22270594 => data <= (x"075cb6604db0e6a0", x"24f3e1357a7fcff7", x"e2ec29bc3b8f33a0", x"8f7435ebf1dddfde", x"1b887cbe0a2714ee", x"324fbb6899771e34", x"98c34dfaff358cd5", x"f75477f60da0aee3");
            when 26803366 => data <= (x"ceabe6fc418cf1db", x"5bfc61a4952519e3", x"1da21fc87e5e91ff", x"4d2f8a43f9761800", x"7ce58bff3a08f234", x"86150827c00edc05", x"34a66d19768f0933", x"c82beb25f6d961fc");
            when 13442988 => data <= (x"3dd84d75707c8f67", x"6e04dd6c10a95797", x"4c750bde5a461cd1", x"f5947126a882532a", x"a4498606b7cee9e9", x"2739a03845759433", x"fa850f4b65d984a5", x"de1de248e5a6f433");
            when 32702530 => data <= (x"68666a4ffcdd8049", x"1a6d4f79d46aabc1", x"16a59bc1594ad84e", x"0dbccbdfa2c82d6c", x"268cd29fb24c6fb3", x"79aa787914e46558", x"61aa5b3f4dd695df", x"f7b0e5cff1db5394");
            when 11405839 => data <= (x"cd565135be475f95", x"100b825b9fb41a77", x"667a4da1f2cbe0ab", x"31464e6e915c8731", x"82140f2f26b350b3", x"a28ca558c2c047e9", x"ac0b98179b9eeedf", x"0771d783b7c67a4a");
            when 8897460 => data <= (x"4c8ca8f491495a87", x"1c9066492fb8fba0", x"50036f3a6ad02dbb", x"eaaeaed34e4aff39", x"03046c010719a883", x"7ad5ffe5ccf71981", x"67e20ef1dff97c4e", x"f3f73515e4c1fc03");
            when 14954369 => data <= (x"50a8b4f413055fa8", x"6a395d580ba1746a", x"997072b90e8fc871", x"44c7732822007ee2", x"c187b3f2fb7a1178", x"ce8e2f0c277d4d12", x"dca96cceebeb4b6d", x"3aacf3331259bcd0");
            when 18171845 => data <= (x"0dc8fb2775c6c90e", x"4bb0603abd6acb27", x"affc013e11de09e2", x"7d0f1521782b42f2", x"34694dd508263b50", x"c503494de7c2bb4d", x"94963aaf64ce2022", x"558017b9e7a671d4");
            when 21227057 => data <= (x"8884e5423bd38f49", x"aa22c4c5a79ea418", x"7ed891596f637b2a", x"5e1c2e7d63ee1b3b", x"6daf125be57aa865", x"4d341854eb8bbb3d", x"93b4afd226ea276f", x"e80acd54e2fc52ea");
            when 14126685 => data <= (x"fcb0366c41b9927c", x"79df2ee4907bf431", x"a30893bc11edbba6", x"382825294153cbb4", x"1bb1c3826dabf944", x"c3e0a257274fd784", x"9d0ac63de6a7447d", x"1c7164839e73f09a");
            when 32531430 => data <= (x"2a82c7231cc9700a", x"b4c935c92c281db1", x"c02703fc9aa8f806", x"6d8e32576061a684", x"9ee05c2b9617da74", x"f21677ff1395ec5b", x"315c89c50d49acd3", x"0480ffdad1aa0e36");
            when 15058371 => data <= (x"3a22c6b414ab3e74", x"805b6546804012c3", x"104d805cddcafaac", x"0ef8337bfecf2515", x"9524d76fde81724f", x"5a5135b492d95f72", x"efb9198736153b51", x"675009f213b33720");
            when 16034529 => data <= (x"b1c8c21bc832cfd7", x"5ccd351a3f2e1d9c", x"5238f841828e7aac", x"8b907eb9b6faf539", x"44c29d7e7365edc9", x"eb68dbe0abd085a6", x"c6764e2583d94bc6", x"799b1a39577d7b1c");
            when 9563779 => data <= (x"2d11762ae397980c", x"78a1ed0c83f225de", x"839159155ff05fd2", x"bfdb1c6e61ed9f62", x"803e450d06e39eaa", x"7f91443591ceb720", x"cb6a7a9e967a5c9c", x"1935d573f294bada");
            when 13612057 => data <= (x"b36752a791eda2b7", x"f113944ed3a03688", x"f4ca706fc481b678", x"2ac341c6f3bc2d81", x"82ef1cb76800e089", x"ed49998656ca8660", x"023cb66b1e99b1b6", x"126a451c0357a381");
            when 10729192 => data <= (x"747584a6f90f94ef", x"833540db95c9f0b0", x"d25c16419bcedb84", x"2deaf22d9310c8a9", x"4a2fc724e51a02d4", x"779b58c8f824417c", x"575c4148ccdcdbf2", x"2749a7218806dc76");
            when 24226407 => data <= (x"e567e5c804ed6a8b", x"243391c6d4baffab", x"da9a1f49a1553b61", x"faab009aadc9cb88", x"c8f8f49d9c63681d", x"6036af28a435643a", x"e89c7d6835fba604", x"58af7cc53912bb78");
            when 30141575 => data <= (x"7bf25cfee8ea8505", x"55b973a7fe824bc9", x"20027bf9f695e382", x"3e2345b72959d42e", x"9e9dadadfaf9f0e6", x"9ce2bdbedf97eb83", x"616cdf52f98061e8", x"16e0a22a827daf33");
            when 30834999 => data <= (x"3d7e55ba3bdd2f63", x"1d6fa53f90a46f87", x"61df5b5deb6a2e67", x"0a79ba5e2b5aaf5f", x"7ba4210ad50c4af5", x"4a4e7dd6f17e9a2a", x"8813378a77da4979", x"eb28082bcb7a7abb");
            when 29716226 => data <= (x"65b440158dddb324", x"b456657c5c891fc1", x"aaac69f1ce0b29ae", x"fe95a5427f9dc917", x"3800d42a44fb94b2", x"d6b8af603cabaf95", x"be269ce14c7915ff", x"6afcb746867c3a8b");
            when 30703175 => data <= (x"a15e7c711bcf8224", x"54efd20b2644f830", x"77a74da458335f33", x"82f5666ad0245e8d", x"45b00c8c5172def9", x"2559456c75a52b37", x"b63559fa5122a7c9", x"28876f23eeddbecf");
            when 13385849 => data <= (x"974004b5637ba7b0", x"5c7e5d149aabb899", x"509d79caa8a3f5db", x"99ed8e5eb2312a14", x"fe0d1d9b8167e140", x"eb375efdf15d4be5", x"694dc488645aab9f", x"d845e21b358482b1");
            when 8231508 => data <= (x"de38b8d9a3db2d1f", x"9473d079e812c5ea", x"8de6cef550b6440d", x"0ecf3c4841270a5c", x"5a67e5dd184d19fe", x"de5a2be1bf579e14", x"891b2eb5e0f83442", x"4a8901899875b3ec");
            when 12134309 => data <= (x"ac3243974d968f54", x"a374119af242e3f8", x"a07cb90f88a29d71", x"19d3e8bd2cd862c0", x"b521edd9d5c53f98", x"431a98959720fe26", x"6c14609ce9506fe1", x"256de02dfe2eda9b");
            when 6204589 => data <= (x"e66d02f00fd23105", x"bedb214e9e42e1e9", x"6ae300f127d1ea92", x"14999ec3dbe29679", x"bfdadd967e462de9", x"31bfb098a20f4bd9", x"9aed4fc29a192c97", x"6041cff4dcf1e5e8");
            when 2153357 => data <= (x"c037460e1129092a", x"00e0435969392b40", x"77e0ff4985b57a41", x"f18efa271eed34d7", x"7224c2b69b521067", x"f06cfd1e1c5f7b3f", x"ee0077c72344c024", x"5c24945be66f3077");
            when 17169564 => data <= (x"bfeabdedc70aa420", x"2a8458bcc066e84c", x"f22234d6f94913f6", x"024a4b3e38bc6e03", x"b60c8914f9c51988", x"0de375fa6bad4cdb", x"a2dc377df302406e", x"706b5351a1657458");
            when 7151017 => data <= (x"21c537c23b21b8d7", x"4c5357d5746ab491", x"55c3fa826457646f", x"787b3cb967554c56", x"10e8230b0afdd704", x"1e1eb4f69d86441b", x"979386c34d68530f", x"e6b1630a6c0a3128");
            when 32282440 => data <= (x"acc2f320116c420f", x"4b097bbab2b5d319", x"c28d2f213a88bfab", x"c21882872bf15df2", x"e4adbd3c4c4f349c", x"d192c87143ec7429", x"e2d0d01a5a2e4f0d", x"fbcce9b6d3ef0300");
            when 11077147 => data <= (x"6960c8cc615ee773", x"61572484ac1fa610", x"9fd5ef1d3c075506", x"712eee3a660cd8da", x"3e6f5b421ba2c838", x"eee767018b12a3e3", x"9fa4a213631bdc19", x"0df45de2f56ef9a4");
            when 32887119 => data <= (x"d1942621f5e6ed0f", x"79991f38941f0ac2", x"f11e99dfb4c771a8", x"305e14339880d067", x"47c4ffd2db294496", x"ee86840418d69013", x"2ed792267a3429af", x"67737a83a89ce66c");
            when 24350028 => data <= (x"63e42209683d14c7", x"c70c9519391e4b53", x"adc06f7b38ecf690", x"d254acd8f2e1d556", x"3262340a232646e9", x"94256781e3af9314", x"1372e4436c2ff2d8", x"f6756d6657609d9b");
            when 3792492 => data <= (x"1184ecb5f6ac162c", x"4bbf7d1a5228e800", x"c574b3ab164e2e24", x"d5af2c3d8ebc207f", x"d01c93e4676f7af4", x"9ba7173ada4bc1ca", x"fa225f4a210f4375", x"8c9dc6c23a7d5d34");
            when 21531605 => data <= (x"40ce737f2e875fe4", x"adb5add998deb08a", x"0dd112990ce07e76", x"fe38ca00a0e8abe1", x"c94c33e41304ff74", x"64739ff4116b6245", x"b960a67c78bcd658", x"fd747903b89ecf68");
            when 2929738 => data <= (x"e4f219594125f300", x"121f4446575b03b9", x"afc13138180eadd4", x"13e597cdd7f7aa30", x"82444b9c9996a5c6", x"50ffa0ecc625caf5", x"e67b600641200d1d", x"22049ce2e49129d8");
            when 15848629 => data <= (x"559e9fb6bbc9cdc8", x"a6cb08401cd76fcd", x"6683b84f89d49a8f", x"b79b36f379e7baf6", x"d50b0e8767c3c862", x"6594495499d6c4cf", x"5e593bb2e9882e30", x"4a42bb95d1248922");
            when 31216622 => data <= (x"b4b5dd9cde066e28", x"81820b5947e6b973", x"8f72399a7c92c45e", x"9935431f090db048", x"370d1707fde33491", x"f24cfdf7733b2e9e", x"202f4efa2d568c9d", x"97902ed1dae6010e");
            when 32002368 => data <= (x"08fd737c34e7b120", x"cd95915735a30eb0", x"6b0da417bb2c0da0", x"afc884550ce39e3e", x"576dced7d1826e34", x"00718ae6ee4d062a", x"23d48996eee1f0ae", x"203aec237c79f19f");
            when 32390759 => data <= (x"f4fb23eb46ea63c0", x"8e94702dba8005b2", x"88b08912464f4c9c", x"77ae30bb23391b2c", x"8a8b212a1dfda1ef", x"0cb608101468a0e0", x"bb4a9859f97a79de", x"f426332b7675e192");
            when 25545041 => data <= (x"b3ae2375728060eb", x"a4e80e8eb35cf897", x"6125de6251711e62", x"e848bee679bdc389", x"04eeb9646bbfe470", x"7a53c5ff5722fab7", x"4a366dcef876303f", x"ea46f3ed584f1d94");
            when 19626322 => data <= (x"fecd511e233ce984", x"e759f3453bccf64c", x"949287c3f29c1836", x"9377e0e1b23a5db7", x"2eff36487841769a", x"ffd9b83f72cf5301", x"8119613b7f37363b", x"08fddd1fdb08aece");
            when 13716495 => data <= (x"76b140a2e1abe4e2", x"d870f74c03dd67ba", x"10fc77071b21ec40", x"fc584f64cdb6c5c9", x"edf508357ce34fee", x"c883a7fb34070ac1", x"6b464b1d6bf57876", x"cbe06dfa71ce206e");
            when 4031490 => data <= (x"06e7347d9664c113", x"3ca01e5a0026e4a0", x"91a1988666d3e752", x"f2e0794f0a725e1c", x"cb9a7b47e49f6331", x"ed82e4cb44970ac7", x"447d3a08787766d8", x"3ddf1c41831fbe67");
            when 33476011 => data <= (x"1d4b3dbb8e551ae2", x"e297789d905cf6a8", x"2a6d409ffbf018a0", x"90f470d534de64a0", x"ba05ea44bf332ba5", x"0bc3dc2546b5497f", x"e31eb4cea6344725", x"741cf1416ff72c9f");
            when 2070194 => data <= (x"a1aa9d4bf4a2bc6c", x"786210732d7967c6", x"20947c585b7df297", x"2dd4b7f91aebd694", x"f5ec0d38a7232a44", x"6e03b46758b2a8e1", x"3d4fecbfbb1a3edc", x"539600bbada02bb2");
            when 2455139 => data <= (x"d27da77f8bf98e0a", x"d78849c2ae1d5434", x"cafc071fa65f275f", x"26eec32d7ff7a1ce", x"2c849bdca8556d02", x"e5c2fe71700f5a8b", x"bdb8bee80d5ffc0a", x"069e0a7c65decbbe");
            when 21788585 => data <= (x"3db5b43f6bb4bbef", x"4ae718441a1c22aa", x"a0d4ec27b6995570", x"1f2009aec9a14c55", x"d934557b77070d4e", x"2e8c0b53eb3d5cc0", x"1e647a9ec01fd7ba", x"51bc1a8dca666669");
            when 27827940 => data <= (x"f6038f9464b0927c", x"b74d14318583bb32", x"49b795533c1e2a68", x"230cf088c716a03c", x"a1ac7b4e205e8b52", x"4929df15bfeecbe3", x"18f8ee3c96167813", x"a168741984161186");
            when 23252346 => data <= (x"4d2a4a993a5a6455", x"b9911ba6c1fd9e76", x"77417ddfb11541e6", x"cfcf706a409677eb", x"a972c6128c7398cf", x"5445f1b371b75fd7", x"f9b3147c3dc2fe91", x"e9943c949ecb6e63");
            when 15622419 => data <= (x"def6f4c17bd495ed", x"975678178d5cc3e2", x"0842e0b1f92f4043", x"0307481e6d041f12", x"fdab821c3c780cbd", x"d6c229ba290a6638", x"7aa40b326edea465", x"faef8799eca137b5");
            when 8084579 => data <= (x"98686ab3451b72bb", x"d8f6f732d88585db", x"b30a83635a015a21", x"c4f575b02e65d05d", x"b4e97ab105a5ef77", x"bf9f290b09eb7bdc", x"61821f3acd213af9", x"b03754db3531806e");
            when 29265519 => data <= (x"12b40e9c617e6713", x"432ca9f9c78dc18b", x"29c12841b8bc0bbf", x"61be6be76391e8aa", x"c1a4bfc499226e58", x"107a61c06809cffa", x"605c9b18a3ec5849", x"a8183160437193f6");
            when 6505535 => data <= (x"2e99d78deb847101", x"6b72cba684a48f80", x"d1bab7c2c36b7ad9", x"691f171475e99f32", x"bd15c20ebe52dbce", x"f3ec8206e816806e", x"ee3d6c770ccb6359", x"f6238730172e78fb");
            when 16409297 => data <= (x"83a752ddc00b6dfd", x"853988b06ea9f7b7", x"4ac15b9bceb57b14", x"99cae36a72e5e3cc", x"a43f834dd902eb95", x"fe53591b6bc3c666", x"a270bd4de1368ee0", x"e2ab6c171238702c");
            when 16391198 => data <= (x"7d42f7ad06836e80", x"ea52d430da68692c", x"fff3aa4950eacc6e", x"2c447e4beee7491f", x"ae23b5def29517bf", x"39924605f0bff116", x"f54fdf0278650987", x"b23c7b6061af8c24");
            when 28608006 => data <= (x"a018b404766a2dca", x"1b7bac759a86392c", x"0512d10133c93ecc", x"3d5e94cacca1ccd6", x"49a4e1b28949f658", x"822413c14312757f", x"d8748b5876766cef", x"46a858a0b3589b4e");
            when 9789595 => data <= (x"0103906231c9b84b", x"62f801d870753e49", x"9b8f0ee13bb4b585", x"ba459682251abfe7", x"4c950d2d9cf8bc84", x"672e5a062d7a761d", x"d89be0e08ce065ba", x"bb6e6b991eb3f567");
            when 6219818 => data <= (x"cafc495f6fb94a73", x"43bd879c7e74da2f", x"de15ba141e4cb1a3", x"c54bc45473235ef7", x"ed05c42648e9f135", x"84a6ddd91cb99708", x"faf21b350d5f3e9c", x"d84210426f620b29");
            when 10855679 => data <= (x"6898ee35875911c5", x"2a74d7502985d2c3", x"de4bf45d04f80ad9", x"de555cdea84b6068", x"39ee9b9bc06452bb", x"070aeaa41437b16c", x"c51f9e15a421ff06", x"6af18131d9bf97c0");
            when 7710679 => data <= (x"cac78163a8335a10", x"dd421b92afbfc90d", x"85b82052d3c4d36d", x"13082adf9b8c7ef6", x"26a2f15f640a4eb8", x"3248796158b53ec6", x"764479b23520819c", x"9097d00dd8bd1d4f");
            when 31240179 => data <= (x"f7675271730a9fac", x"8b57126a1754bf40", x"a8e3bfdb72c1ef74", x"b15a16fe1d875268", x"16ae0ffab64b68c4", x"0d09eac84dd658d1", x"c06dc2c1c4750243", x"180e0fdb7d245cb9");
            when 22725864 => data <= (x"b218bc8dd4941d5f", x"878859694e4cc589", x"5adf01ca78fb49cb", x"8d6c0b2c6d4c49f1", x"3252e443bfa39f18", x"378ad77569fb8dc0", x"0f2cc7a080e2a86c", x"a7369e5d185feea1");
            when 18847950 => data <= (x"f3595caf6f952e11", x"1d68eee9d232cee9", x"1b5545a4850534f3", x"f17596f8653db047", x"71f2f5c69b2784dd", x"faaf87e85374f45f", x"5acb1105c8e27d17", x"775ba5080dfa052b");
            when 975607 => data <= (x"e4f69021e4248276", x"df2b57a24385072e", x"5813b18081fa8d69", x"b9aeb46e04117364", x"e6935e9059c3449a", x"a0a2e0c44eae72f4", x"f1db9eeffa36d796", x"0f11ed8b9a6f9e54");
            when 24177843 => data <= (x"442f3b48d3c62a89", x"cd316e43965d74e2", x"6f41e660d5e0f696", x"0e2f638756539e1c", x"aca6a6031bc296ba", x"2f560be786f8f025", x"de845d104158f1fd", x"7884deaeca09a4c3");
            when 21468857 => data <= (x"16e4db6cca39bc14", x"3c4c2ef08b9f1eac", x"8077d210bee979d2", x"2ecd1552d7a4e3bf", x"611783fa8aea9b56", x"325aa1927f6f8c58", x"0f95a07b9573e80b", x"7ce53366a0e641dd");
            when 22394575 => data <= (x"7dad35ea8c3dbd87", x"21d0c6f3b87f2928", x"58d8ca1dbb07c176", x"1ad8681bce401c0b", x"f9c8f4f9b39f52af", x"113297490e2f2004", x"17d10c38ded4b305", x"f13d8c2c88f42d00");
            when 25929866 => data <= (x"23d7722c94894252", x"6460e35b1cc3b027", x"e1502df8f49d90df", x"b3768aa582bc48e8", x"097622a900e88059", x"537f83be7cb0f826", x"5a81dc23033823a7", x"5e0f890087adc8c5");
            when 1263020 => data <= (x"94d9e82814d4264a", x"497faf5779c3c730", x"60ec83ec18f3f197", x"a2af66dd52c568fc", x"e1148c744e0cf8a7", x"f6b830a873d024d7", x"1f92b5a84427655f", x"13a3e32360cd9749");
            when 5474477 => data <= (x"824a4b5babe98f79", x"f202285e12e027a4", x"00b6feba0d616b54", x"8e02a24ce64dae3a", x"b6ab8dd6c7de3410", x"12428c3af4c7e794", x"ae73d5a1f47e3007", x"d81cea956d54fa91");
            when 22641259 => data <= (x"723aa789ae552c19", x"b3e8b360ac542403", x"641c020ee29b96c2", x"68bb147bcfe443b9", x"9da4d557a67b445b", x"620de3a4d3ccb227", x"60b33657f6d2dbe3", x"6c8e5883e77840a5");
            when 15785273 => data <= (x"055a4e9e00174cb8", x"ddedc69862bc011e", x"97a284110dd2eaaa", x"90f4b620ae0b01f1", x"6ccd77ac25a401b1", x"f0decce80ce275e8", x"1992b4dedf438e5f", x"cf88a5f157ba040a");
            when 1537917 => data <= (x"ba7d4a4b3136f6a7", x"6ce4d278397ec6f3", x"effdf10d16796493", x"4642dac7f6582f9a", x"c6a86c5aea290fc2", x"f9e9bf41f00efbe4", x"928ce7d22181b1d2", x"bfc71893ced0ff6e");
            when 22280134 => data <= (x"81874a4a905b6525", x"6b59cc82e228808d", x"27b49e945fb0c086", x"872de8660d270a3e", x"40bcd8aea9d46d91", x"364f9c1076462dea", x"f44ed467ae0b55b0", x"2da7112126c7b14a");
            when 1763526 => data <= (x"ff456d13e67e9b82", x"3bcaed275bdbeb7f", x"d6962652b28c5b63", x"bbd0f66a744909b3", x"d02754bf2e3d3feb", x"079d3b6707f5ac77", x"bc74e0fbfde66fd7", x"8b410325725e49ca");
            when 5523220 => data <= (x"43698afd07b37386", x"e504c3e22bdcf9a9", x"3b4ab3f775c92b6f", x"02277665eb8efde0", x"777b2dd031d8294d", x"66bf775a2d10c3fa", x"0fd40a60cd63cccb", x"30de562b6f1d24e5");
            when 20219393 => data <= (x"0638beec17b65ea5", x"d4baa7c707abcb3e", x"81a2ec505f07c7f0", x"b326cf6d9fc4f079", x"90588e2adde1f49a", x"61e5436c96f68121", x"d69c8a8b6d664458", x"2e36aad86bf72aee");
            when 14201284 => data <= (x"e6d190dbb1dbc36a", x"c43a82d69f75802c", x"325e119b795803ef", x"4b2ba45ce352a153", x"d45777a9a9312396", x"4a4d8d74efadb923", x"eda1fce49e74a234", x"13eead6f549ebdcd");
            when 19926861 => data <= (x"06b14fa277e5db88", x"86b5281c4bf4ed00", x"3f208d9fb1933b41", x"8c6ef5c9b89d5f0c", x"5907fb3c0f1c7dc4", x"d67b9f01b6d63353", x"dfeb5ab0b832c156", x"f4b4047a4b530d3e");
            when 11812767 => data <= (x"e69d649bcc1d4ccc", x"6a3c2daa212ecddc", x"ecd19318fedcf7e8", x"d2b60008f6f57b69", x"63cc1cac16178d4b", x"50bcb345fa2736d9", x"a10aec6dfc6dae33", x"092f4869686940e7");
            when 5609281 => data <= (x"4105d90f5cdb4c9f", x"64d833d1a7c62e34", x"cff4c54da9624c65", x"dc6058c00ba94ce3", x"adabdce8f2e599ab", x"eeb208c146a5f443", x"a41b058b3f566564", x"451d2a9967ad84b9");
            when 5350176 => data <= (x"888ddbc90f59244f", x"23863d8a0a053f98", x"6320c7f8e297f7fc", x"f857e978f99d19a3", x"cdc195ec4e9e055c", x"9b73a6a3a6277e40", x"651e16665bec18fd", x"b94fcbd0637af979");
            when 19312141 => data <= (x"c0983b76226e4869", x"a900a3b36da37787", x"a5ec2535362bb19f", x"57078a63efd54f2e", x"0dcd826f58ba4d23", x"3041224960a27379", x"74026c841fc6c993", x"f82a715c6a9541ec");
            when 1498397 => data <= (x"8c783c61a954e874", x"1a9b1e6b25e8e7b8", x"13b9204e89759d7d", x"543dface12f06767", x"3f600fb895b9d751", x"d9e7f62bc3b3ab2a", x"4e91ab1592a312d5", x"cfbd772f047f9491");
            when 22247746 => data <= (x"82263dde4d172709", x"ac815f158856b32d", x"2d9b75ada619c775", x"e97b5a4601dc3d25", x"814047684469b193", x"b34a9007321946b4", x"8fe1f41ffe8eb221", x"36515e4f0b8c7baf");
            when 3811010 => data <= (x"4dc36f8158e90c6d", x"9f4970538a2773a9", x"da0a6dbdf52df87d", x"345060c2272256cf", x"777aa9d6c75182db", x"79e18eed1c472cc5", x"d3f15e782ec3f147", x"d4381296a2c4c1fa");
            when 19174519 => data <= (x"e90169bd0d68aab0", x"26d04b85be70eb4b", x"35f6cb8fe7ad9b3d", x"139cbecfbea7b7d7", x"0097a9373aa54e66", x"e808391699f2d8c5", x"658885b2fa3e4f00", x"53de431049b8a3d2");
            when 801155 => data <= (x"a5a3155dacd66a20", x"a928c87f4c9e2d72", x"3cdbcd2ea0447449", x"f9e886517351c1ec", x"4c4f163a01decfae", x"64c02cfa9d18290c", x"46a55a8af9af2793", x"758a61fb0ce871b3");
            when 28624415 => data <= (x"1b2abfb0871bfe3f", x"25f505d8dcae9856", x"d3c20ca5f56feabf", x"34d32806d23b9503", x"e36cd5bf999192aa", x"412fb09319c0218d", x"0d0d79b838ba3f41", x"cf79853a5ac67811");
            when 7589912 => data <= (x"b68a60327f32487c", x"c47ca1d20de6ac53", x"f049f1bb6bfbfc5c", x"5ac788049646ee93", x"bf84ac3152980e45", x"80bf30bd3e749e06", x"87f922988c54740e", x"97851bd08ce93a99");
            when 26955499 => data <= (x"244ffa31e97f1f40", x"382ba81664383edb", x"c210f4ecde2104b1", x"4d456915753ba577", x"71893faa3f0136c0", x"217d5cb669eca6d3", x"e486a20341fe5c4b", x"83bcbdfe1d9603f9");
            when 12545205 => data <= (x"a5977c55d86a2153", x"51c240475e7015f9", x"79e922f409455b50", x"e2b78c596ca3511b", x"8878becdb1aec74c", x"3d965351d6309d38", x"b6643425deffb5f6", x"f9981ada331bcb65");
            when 22363587 => data <= (x"ad59ac2cbe5d3e8e", x"d58117f0dbd5b121", x"dc8a569dafef5e48", x"9f35b85c1f380659", x"aa371f2429525da6", x"333ac5c2faad3893", x"76b654ff1eebd9fa", x"1f2f358fa2cc7864");
            when 30466977 => data <= (x"9ba88a2af605c07b", x"d4f55f692214c585", x"7a1bdc8260c1612b", x"2794fc042d3671f7", x"7d79894f87cfe4ea", x"8a67885cb156cddc", x"9b25fbf00deefdc2", x"1a00f4f8b4b93814");
            when 25306301 => data <= (x"6a4448cfe2052675", x"dff335be21a4bcc6", x"37970020146a3a21", x"fd74277a5ab2b8ec", x"eb61df184db5d5fa", x"b7df666e4d66abc7", x"5814bdc74d8d76a5", x"8cfda3228d8f6421");
            when 14428027 => data <= (x"27bbc58abff01081", x"97e15eb49ae25730", x"9ae12d986077df63", x"d2c97783079f7865", x"4a06b2d5e07a9938", x"fd35fcfdd2cf58c8", x"0d5866f898229ee4", x"aa364549182500a3");
            when 20692462 => data <= (x"3cbaa1994e9e0ee6", x"600724ad4c097e47", x"da61a1715936de91", x"24520525889d8d67", x"2a3287888b4d77f1", x"c3d0ff18f42176b0", x"94606e8aa1a975a7", x"cd41bc74f7c9aa23");
            when 23952316 => data <= (x"12d09ea589ae6913", x"f8fb4717af4be7f3", x"53a0fdd3edabe30f", x"9abec5aeaeeb6132", x"cb021c3c9ddc3926", x"94b8e8df0602f80a", x"6214eef8f7a325e8", x"fb81672591147704");
            when 6219134 => data <= (x"138b417f519bdcd0", x"2692e37c4313574d", x"fab0ba27a758e194", x"65f225c26d474ce0", x"8269f2a3a705676d", x"96c9af95729d120a", x"4a14c133e6bc1cbe", x"607a493040880300");
            when 28458680 => data <= (x"e980ed56f303a338", x"d22bac1e9d99edb4", x"f28714478c9a6c09", x"6675397045874428", x"a6f58e9f3e8a3ce7", x"e762a77ddfe426ce", x"f46c40d7c9d8d8f1", x"7fbb28e610c3aa7c");
            when 13055172 => data <= (x"9c0005302dcea3d8", x"ce13ba44215f713e", x"32b43dd39f845667", x"e8682ad70aa8821e", x"691c3e4dfc2a6e74", x"58651a79e96adc0a", x"6898daaddc3e6fc9", x"4879be6abd1eaf11");
            when 18623722 => data <= (x"67b7b1c49855f4e3", x"afae7cb2a0e6ce95", x"b69f6017667dd7a0", x"ec2a5b78352d41fd", x"0c5359106b1c7ae0", x"c9513b79f23a7a3e", x"1bf3669ccd64d9c6", x"54dcf4e8666f3e2a");
            when 27090079 => data <= (x"1726a7147311e984", x"fb57f5c0e6494c2a", x"c529c15a2d115864", x"69d1aa921072b6e9", x"d88a202f4e2d0a2b", x"69396834b0f335d1", x"4590bff9bd6a5f56", x"d20dbc3027b4cdcf");
            when 25839639 => data <= (x"6661943617a45991", x"15aebf770fb2cc26", x"9932eae5d4cd063c", x"8f345b2dc13cb56e", x"1ad0a17b2717b67a", x"c61be83802b8fe9f", x"a72ae585be76bb87", x"c12a7a8d9ad61c99");
            when 27028011 => data <= (x"af4abbda0917134f", x"14b88361e1408901", x"04807acf61f84051", x"18695f1b3b4c8974", x"7c836b07b48f17fd", x"001324a80cfb5225", x"eb128c2b8e7aa47a", x"3c9bc2aeec363d9d");
            when 12137294 => data <= (x"43af42f59e37db18", x"e6507b827661abad", x"3af2e03fcf3aa4b5", x"8ebb7dd746c51a78", x"d079b356f3e0e687", x"a27b13ffb5e1d244", x"3afd2dc3c98f3eef", x"ad98a9747fd4f80e");
            when 15760682 => data <= (x"42845c0b8e814a4d", x"cc94fcf72bc4915d", x"7f7d25b4bd8d3b85", x"fb8d95508b8d0960", x"6745032d1762ae3c", x"846e03e45aaf8364", x"143a1c1cb8a3d483", x"f786bb4584868f12");
            when 8740015 => data <= (x"e72f7b1f7070a936", x"4c496168834f8cff", x"ef8d419ddfc5ce8c", x"1fec8fe4d6860a37", x"74d3dc9bf662b3ff", x"34be717f6c255045", x"04d1ee0dc4a43124", x"408d22fff18a2017");
            when 21352920 => data <= (x"6a9fbeb9190c5c8b", x"505acdf16fca1a26", x"5e870a896f3e5630", x"582d2e596119b78d", x"fc643334203cbb4c", x"b0107fcfdd8cda42", x"5a6ee797a968e530", x"21825b5e1cfc7006");
            when 6382933 => data <= (x"6f05dfe5ef65671d", x"47d22d0a434b6188", x"57eb3b77915fd293", x"b4c663a0abf1da66", x"d609b6d70e60b92c", x"e37f319250cb34f0", x"19dc637091d14e34", x"57446c116382d205");
            when 7606114 => data <= (x"2740e5b0bd7e4d78", x"34a5360959f47d19", x"a1fc6ee61ff8d9cc", x"a924af16b4817bc8", x"4525db45c3bed088", x"8f72c4102db6df4b", x"2a18fbaee44d2a88", x"9ecb97de719cbda0");
            when 13643785 => data <= (x"3cbb9744c2fc5ead", x"8a867be77de3ccba", x"22f327156c1d02d8", x"f71ff3718733d277", x"08ce6e1484a560fc", x"bb899fa6125ff608", x"2a69bea1a3e1b610", x"6b1202adeef2164c");
            when 9148433 => data <= (x"99dff9946ea5be2c", x"e0878149d6d175a6", x"8fa97066b344fc99", x"1343b7b2b93b5d7c", x"73f9fc4fcc0a2909", x"be890c3bffda248d", x"40d6a06fa1cce4c8", x"0dcde67275ffd39c");
            when 22741802 => data <= (x"91b9444091447d13", x"311005eb3d71fe84", x"84b5d480d300693b", x"d51dd381f85dae3f", x"12d1f5686a10987b", x"0de147f69dda0249", x"2735e9ba70e8a7f2", x"ccdaa89a233dedfb");
            when 13637730 => data <= (x"0b05d1e534eba79b", x"33873cf390f8f25f", x"42a5c93b70b78807", x"f2dd616a036a31db", x"6935b9de9c90c150", x"fd5e0b6cdb2be0da", x"ca8aa37031ff2cd1", x"095c7c41d3648e35");
            when 19104142 => data <= (x"d2d7aed907efc467", x"4cdc3d849e8b1b0a", x"1ce3b1017c25e041", x"970dd26b854e2d60", x"8f992f31cc5603b1", x"1cb24571f928b194", x"369f29c21dd3469a", x"5dea5d4623b2b31f");
            when 12097816 => data <= (x"eb929ff32db762ad", x"e80f2fa3a53c2520", x"9f7d5b0c8580d705", x"98f878dbf655f147", x"8878693e09462baf", x"e0fad9ea677f1ae4", x"b59656db4830b5a2", x"afe2562f665d8441");
            when 30064743 => data <= (x"c772b490403eb1d4", x"81b0c3fd4df54509", x"69c79d72fadef6d6", x"06c2f5a76bc55198", x"1e1f0357ee6c969d", x"7ef7e4fa6661e9d5", x"eeafc44cc1cbdb3c", x"5d6c3b99992ee2a7");
            when 12023959 => data <= (x"eaa629e4e6093762", x"a1cefad676942d3a", x"4394b3e9bfc3ef89", x"a19a2d9c0e1d77a8", x"ce9dd8af8b9dd73b", x"5c4e9c35e1cd4033", x"2c39a7b395816328", x"c0b8e8be98975a07");
            when 11723245 => data <= (x"e1acefb56ad210fd", x"da90848ae889abda", x"ccbae771e81a6fe5", x"420725b9e77eb7ae", x"bcb1cb03a4946705", x"373479b6e863f982", x"15fe82c740b8c2ec", x"6d45d0d98c9c098e");
            when 757030 => data <= (x"4b4bd8bbada18859", x"e9f8ac93b33dab58", x"6cff42b9472b846c", x"d08b77accfa13314", x"6fe0e50a3b15639d", x"1d93cbf2680ff6c5", x"59417dce542c27c8", x"6add2ee51b3c5bbf");
            when 4358003 => data <= (x"8adadddd60de4efc", x"6ebc02f33ad2df7a", x"b6218d8931d67e70", x"8fd82c133652c3fb", x"76109bc80fd15a1c", x"980b1283d5822d3c", x"feff90bd2bdaa81a", x"5e96816ece0c6285");
            when 30729445 => data <= (x"1c4fba9dd0989bde", x"aa2ce262af52589f", x"8eec3f2a7e338889", x"cc083a0d29ef0ff1", x"65daa308774f7d63", x"fa38484a96dd4f40", x"f62c498195dac324", x"9a46a1ba68273c1c");
            when 21695268 => data <= (x"2e7b7fb1bd98bc00", x"d9021f1f1e0f1d77", x"7f99fd5c559245f9", x"956e88712a271383", x"77a65fddeba620aa", x"aff1460aeaf1dc05", x"25db5ccf479ebf3e", x"cdae48ffe7c6dc26");
            when 32354647 => data <= (x"b5bbb364e83a99cc", x"aa3f5393dac0f523", x"170d08ae8de4f670", x"ea15078c2824e9a9", x"4b1879d0160f9c88", x"700bc5d334506fed", x"cd7d3084ed5b3199", x"4d93f4046139d818");
            when 19806010 => data <= (x"0f1cb90ad42eb66f", x"bd51d81a0a09c2f2", x"a9b71673a5efc44d", x"76fa7884451500e8", x"b47443a6927f7b8a", x"b8122430f68ba653", x"061de7cf88d6fde5", x"ab563b411ad39d1b");
            when 31029134 => data <= (x"f68c361b397f4f24", x"f821902521fe06e5", x"3eaa3f241d549ba7", x"02eb4a1d18787fcd", x"07c6109159ec3938", x"761d1644deafb58c", x"6454d835c6990ba1", x"c3eabe569921114b");
            when 9541541 => data <= (x"9eb9c3a02b74a087", x"d83263e8af05bbe6", x"b4b96edf0e121c38", x"d22ef7286f84964a", x"99658ac73d096f0d", x"01c816fe3d42ecd9", x"37a984b9252b27ec", x"1a122a3d324cfe81");
            when 18474841 => data <= (x"dc192e0e85f84963", x"85d96edd3a062406", x"8128234c7aa106a8", x"294ad33216e400d5", x"fd2b603a240748e1", x"89fe1ada7337404f", x"1b828ce74a0d3947", x"011a45e6dae43189");
            when 6273655 => data <= (x"15044a35ec343fd8", x"be19ae0f707e484c", x"8ec054c1840c42b1", x"04f9220df88805fe", x"ff3c9306e771a63c", x"37576f42ceff7fc2", x"976c96dbd25f1c12", x"bb257866a75fbfa4");
            when 11336272 => data <= (x"52b0c4f1048696ff", x"351712d562c8b722", x"c011957a9d3aa62b", x"48aef7c66a9cfdc9", x"62cba4686a8d2535", x"18a5eeb791badd5c", x"3b6d8424600b7ad0", x"2be142f36edf41aa");
            when 5398303 => data <= (x"bf5c55f8602750d4", x"96e3b168594367f9", x"0b4f5f8a4f5a4aba", x"90981e322cfa7a33", x"a51887faf771c582", x"d6c07fc2c2a56728", x"ba969bc64d2efd42", x"b9e2b082e51f1793");
            when 7956419 => data <= (x"d37ed6d9cf1f2516", x"50a8500bcfb133d5", x"524b90437e5c2020", x"b218c31e0923207b", x"ab99a20a867b3b50", x"59732bf5e73cd48b", x"b4dea6836ec9a447", x"fbfcf31f0f202f43");
            when 8124586 => data <= (x"3abbd38d906ddc1c", x"88fa832b5b5c1c68", x"1d0a43f4bc22d483", x"1a315e0eae91306d", x"a53f07e4ddb2e13d", x"4c1442abd403ac88", x"f17209f6b58f85c1", x"ee311e5f9b11b029");
            when 9079151 => data <= (x"42f2f44d93d858fd", x"23a7157fae4a61f6", x"712e6b917e472ead", x"b7061c1ddef53f79", x"1eb66e54bd43e46c", x"8cc27c09b8fe7b58", x"aa3fc4c2a3cbbf13", x"4f7273cbb15fd253");
            when 26942889 => data <= (x"30b3ff1b483b47e4", x"84d52946fe1e88cb", x"13405627add5c185", x"e8cf2a84ebe8decc", x"234f78007291745d", x"174e9700616aa10d", x"06f3df77e50a8592", x"8bddca99c4513aae");
            when 12431955 => data <= (x"2e545faaf2d1c5e7", x"abffb0a888e6e5c8", x"3c571caccb976661", x"67fc1f3a6b6d69df", x"aeaf76e6e7a708ff", x"21b83b30d532d6e0", x"4fbb0bfb8c2ef156", x"be0572adef3dcc89");
            when 19750468 => data <= (x"62b73ba9c1dba386", x"77d4a185e943b903", x"1a7e83c0ad9e6b74", x"dbf2e9415453fb72", x"2020a213bc65f50a", x"cc16edefac934838", x"c75d4281d931cc58", x"984048e1ed5c2b80");
            when 33373648 => data <= (x"cda67b2660bce82e", x"5c2513235ae4319f", x"44929d98a7dbe8a9", x"a89b6f1ede332caf", x"c0fabc1129d28ed9", x"e63f696f01ba43f2", x"0313f37691644d41", x"3afee0b64024abba");
            when 30354562 => data <= (x"fd9b8966a1fb9c66", x"99b70c773df338a5", x"764ba2cb763a5297", x"d7c179d9b08f79ed", x"52668c0967d7447e", x"0bc9821a1249412f", x"5748c2ab224e4b72", x"0f0a5e382b62aa2e");
            when 32436967 => data <= (x"adf869033b1ba43e", x"1704fa1803a1fee4", x"27cbf70e29551b07", x"f0c5e12bf4151c07", x"6c6153de846ac5c5", x"adf5050ae2fd5a6c", x"5ebebb3e5b82d0d2", x"f23726e9f5420817");
            when 10950583 => data <= (x"29bf102537f385ba", x"ba81824ee410225e", x"5ea41d97c11c96cf", x"07c2326ef15b4ef0", x"7bd6195d8884a245", x"b7f91289888bad11", x"7f915a09c96d7a44", x"232eeadf598bb7ef");
            when 9608232 => data <= (x"19e11843668c02e4", x"998d88812d1e5a83", x"a8c635f2abf4f533", x"00bad428821db8d0", x"7bf6ba15e1678d2e", x"40d1b56a9f11d712", x"6088cdc2098328b0", x"c372b5800072ee0c");
            when 19101995 => data <= (x"a5e77b647cce92bb", x"472dff5b39bd212e", x"738a0d0d6b744257", x"89a20e4ee18f9d55", x"412922d7252011ab", x"aec87f2204dccff4", x"ef28715a7052c1e0", x"2293b1a8d58463b2");
            when 31506361 => data <= (x"baf002fd0ba4cb99", x"e5e2b6257ee3a40e", x"60c7c2d5f9e65bc7", x"ae445618c4f8a2c9", x"80d5083572913118", x"60dca803f0bb12e1", x"3a31b8d732f442b9", x"416659d22b9354c7");
            when 25438156 => data <= (x"ec8a8524e2984530", x"811a35d97a34ad85", x"afcedde24cbfa98d", x"cea67c38ce20c168", x"965f4c36894abab3", x"f73f1c52f3dd663a", x"975d01fe143ec12c", x"132aabc9f9bad3ba");
            when 1292126 => data <= (x"fa79e1b8db115c45", x"cf025b4ebd80a159", x"360e0f9f80d4af3f", x"37a6165a9613f9b6", x"1a7e5fd6e74dd59f", x"7ba9011772aa1456", x"897103e52faf94f1", x"943fc15a2bc3a321");
            when 7013455 => data <= (x"0eee76813c939f10", x"7a35a9d60006b824", x"cfdf3477658a3897", x"7090bfae876202cc", x"2e96c39d4c88640b", x"c8e4e422fd6e7db7", x"6ba43a14eadf51bf", x"22ef6bf53163d250");
            when 32311323 => data <= (x"e0eec4c29a36873c", x"13b44777535fc72d", x"87c6e77ee7442959", x"564edcd8fd9ac749", x"9f1aaa0ad62fcc22", x"c462f62dce06c3f7", x"b7182445c686c259", x"7f46da407a126f01");
            when 23075123 => data <= (x"e18fa75d86e40974", x"07879015962cdb6c", x"e631cd20e06c3ba0", x"4f9e2727efd9445f", x"8472a40854b6f104", x"4497a54f2506a425", x"3e2211ee3fb4ea36", x"674a101bc067ef53");
            when 8101619 => data <= (x"d9e55ff15d944c35", x"281d7dccd0d79133", x"9eabb7a5db0e3026", x"772c0c6c56f335f9", x"fa8f018120d48470", x"ab5b389f939d7c6e", x"9ed4a4ecb06bdf1e", x"6efceaa02513d272");
            when 14452027 => data <= (x"8489e4de060b314c", x"8ce9f92b2f5f364c", x"ae557714e74a9ed3", x"827b82a8cda9e164", x"36817bdbf027b14e", x"0331545c75ca8cf5", x"2ff47ee611c03351", x"9a45f3c57d847052");
            when 11140838 => data <= (x"e93f3c5ca27c78e4", x"4cdec7d69cc04886", x"e201037b137c839b", x"4e7a2f6e30b27634", x"0e91d05301520f6d", x"51b990555232b1ca", x"eee55d9963f874c2", x"c3ba4a6429c4b754");
            when 13954467 => data <= (x"e22af27ae7890f4c", x"b635b3132b456b75", x"dc12a6c448a974c9", x"198b17b0dfc3998b", x"0b2e6daa195497df", x"38bbb2d0b3985528", x"f9fcc58828694946", x"bbf00b95e2d3a6e9");
            when 33006219 => data <= (x"e6ff635f33c9d5f4", x"7cdd05b8793e9273", x"207f93efa01c492f", x"6a2b4e36e75915dc", x"27f39437efe4c301", x"efea1908e27f7976", x"7f2d9b410663bef0", x"7f51d5c6d1a9b03a");
            when 29048682 => data <= (x"b8dabc23d0caf03c", x"c0f6f883ac13cf6a", x"2c042e6b754794eb", x"a36f1cadaf44c83a", x"16452bbc330e29f3", x"98846efd0185b7b3", x"c84b02dc7363c3d7", x"2e727e07091143c0");
            when 3785012 => data <= (x"53200799941836a9", x"8da42c1f679f06df", x"b02595ca6a07f701", x"c8128ba7b749efbf", x"b165cfc6aa25d37d", x"2d579c87234688ed", x"7435b06f058b8057", x"656ab34bd1144f46");
            when 1570966 => data <= (x"325222637970b454", x"2304f5260d59c61b", x"b533c55d3e22e6a4", x"a2c9289c789bfd90", x"cff9699a9f7e66a2", x"11434dfd0bcffb60", x"6504c401f75e5fa2", x"2b88f78588c6ee51");
            when 30598297 => data <= (x"33af5a6a4961a8cf", x"546c179fb3f135ba", x"9894ff2d0fe58162", x"953ab43e35f044cb", x"abf75c94652d9077", x"a8ea115868c3e74a", x"431de10e09975e70", x"3930444a50cb4ce3");
            when 31805946 => data <= (x"52aef646cc846c6f", x"ee1af00a59bdf8e4", x"c21728e3842f6066", x"fe8a5af62c2222f6", x"535762e8a6242f6e", x"9cff6785e2f2d03f", x"1d36ca6143113879", x"8200447519b99dfc");
            when 29436461 => data <= (x"39406970d94682d0", x"d81acfd94894a167", x"9770e25797b5ee5e", x"59fe5f9ad1f08e08", x"5d2a27f2579e3997", x"6c4daf77994428d6", x"0f110cd9eaaec593", x"132b0e0125f8e710");
            when 25799696 => data <= (x"4fb675d1b91bd6a5", x"1cefa0bcac64f9ce", x"5e2cea717d46cece", x"eb22106dd1689367", x"0e4a0acef695a901", x"0f8e7d272b827484", x"a8af10ebb6d38c51", x"8010f7e4faa52ee8");
            when 32938622 => data <= (x"dba364c66024aef3", x"58ec89ec2f3678de", x"baaf6f83eab93608", x"478fc4208b95955d", x"ebca75ce97ff83ae", x"4e8228e97f53b2e2", x"40a1ef3e8a359b2e", x"9bf3830e92207a0c");
            when 16025607 => data <= (x"082296452f78b6e9", x"0c62f2c9acbf33ad", x"b161587662f168cb", x"be06f750b8b3ad4e", x"918b15fadc9991ee", x"640235d2df93c44d", x"f8dddbba77d0046c", x"60c625fbc000251e");
            when 7965882 => data <= (x"3d71541ab73081df", x"8be40d805414e9c9", x"3885f15f4a7dbd6c", x"45332af07039580b", x"1e3f83d239a1a112", x"3b499ab52d5de001", x"341ed2a3d1f08558", x"3813fbd4e5935bea");
            when 33835189 => data <= (x"bc4e6a3d221138f9", x"61558f68931b88d4", x"cda8595628b392fe", x"162d86341b5ff1c2", x"1c5b597330867743", x"9294e2eb29755048", x"9ec01042a8b9ac04", x"5b33a6dc3f946f35");
            when 16529728 => data <= (x"0a9143638d1e3521", x"69b2ab8cf20bfbae", x"ffe652e265719684", x"cd8e019b945bd96b", x"586b182f832dc2d7", x"9cee0066d0829c45", x"e535cfc92ed9f25b", x"15ed6fe8eb0fe1ab");
            when 5088218 => data <= (x"53a7621afdc6ed1c", x"496ecd53578c0455", x"966b342d5d77ada1", x"9733635613b00b87", x"41e98b2863e833b7", x"2ceaf7e644279e1b", x"b6126f676a9dcd8c", x"2ecb6f0229a33d31");
            when 11457091 => data <= (x"a75011996a1389ab", x"31bff1d4f84d373e", x"56e996b843ff2b23", x"c212cba4d689ba06", x"011d5de85eb7172f", x"2fed777e4bdf952d", x"7406ca5ee261d957", x"aa29db1dd341bf1a");
            when 10121983 => data <= (x"e3a959341f3ff1b1", x"3e226cf827dd0ba9", x"7252248812b537ab", x"04e4e29e4c0fb0f6", x"173a205226678cb9", x"0fe3aee3c955e780", x"43d35fe7dd2e773f", x"3e978e92ad21dadd");
            when 10457141 => data <= (x"26e8c11612c7a7db", x"9236ffebea55f330", x"fb5670fef7bded9c", x"9c6a539ba6c597fa", x"1dddd1a7048bb0c8", x"b1d0193316d1a2ed", x"3d53cc45b2db3d0c", x"25e7368310f709f8");
            when 30429652 => data <= (x"5709add61d8a0f6c", x"be0b73020b215b8c", x"5d810abe5ed73cb4", x"0e8e85e0db9ccf14", x"dc1c9fce7904d7aa", x"f61a07b778e9c357", x"138790e56470dd41", x"d4f6b2bca5160cfd");
            when 9172504 => data <= (x"fb554c3a07064be0", x"835485f4b54a8b8f", x"e2596b3dfcdb6ab6", x"dbbe2b87e3e62861", x"4614486e02aae172", x"c868c52e719f0e9e", x"628e09fc3b704f85", x"c09ee86a6246b05e");
            when 19889288 => data <= (x"0cd7f0866fb7ad62", x"49ef46ab095069ad", x"418afea6a6d6ce15", x"899447f2d0c785f5", x"810328db2fc819fe", x"39b1271472d3d4e3", x"e30f81d56f2cb52a", x"bdd25f71ea3c4d70");
            when 32192015 => data <= (x"817f5b6b13e2e2d5", x"1cc7e791271bd55d", x"c708690f7497f02d", x"4d2710dfbd645df2", x"8ae2ed9390bd5877", x"7e5cbeddace44fb3", x"7d2b7a7d05e8badb", x"7af0a563f73a5699");
            when 29071043 => data <= (x"329973d42f43c57b", x"f318605a05be93ff", x"b6cbd5a97acc6234", x"7c07fc2e6dd455ee", x"6f34db055bb5ad6c", x"9b18207051bdd0a0", x"a463c91edfb340cb", x"d9c5847d034857cb");
            when 24426907 => data <= (x"b442049cb43df7f7", x"78bc048d58713350", x"3ae58e8de7540276", x"577d2383313c93e4", x"b93746ac1412a558", x"9ba48412dcace6db", x"dd2bfbb811584318", x"69b853ff3514380c");
            when 22426414 => data <= (x"d05b6aeb777d0025", x"6f27d86ef5802fd3", x"3921c4beef79ca33", x"6b0cccb3fc0705a3", x"c5ab76ee4693c4b4", x"33b8b890c0a97d05", x"7009321f67e6e8b6", x"4583f57a6b9693b6");
            when 26048051 => data <= (x"caeeddf8033491ec", x"59b3cd08f93387c0", x"4ce7be6814b7e1b5", x"3ed95fb4b0bd07a8", x"29452d949150ca5d", x"c707c2afb26cb2d4", x"8409e11f3134cd2f", x"34efc75dd74d8d3d");
            when 7923986 => data <= (x"9991cd903701e23b", x"46a106ce26ddd5e0", x"f5159f06c33d883a", x"8c72046b817c3570", x"dd1efe5ad7c4b721", x"032684b2f90f6855", x"23b42cd903bc476d", x"77983a8b844fe778");
            when 6272037 => data <= (x"8c60167a686d9cdc", x"738524f32e3c16c4", x"353c00049fc1ecce", x"52e2da4eb4c5828c", x"55b9f94f06887e1a", x"f047fbf33d6bbdad", x"9304b21f1f89658a", x"807c790c479009bf");
            when 12455351 => data <= (x"84c770ade448ad39", x"1190e06f7f610ca3", x"f512d66bc0437b90", x"7a84f0fca77070c9", x"7d3e14cf1a539639", x"39bcfab90455668a", x"b720647c4825a310", x"ccc24b449b1c9876");
            when 16418262 => data <= (x"1ec02f2720158611", x"5bc6e6791f314e23", x"82ef8b14b0a75cdb", x"b8bd87ce7fd6340a", x"ada963bfe66f88f8", x"77e37f4ca8317907", x"bd8a3d150ed2f29f", x"070fb0849c971b9f");
            when 26531851 => data <= (x"597897a1c3101cc8", x"73e59d300356226a", x"584a4c0bb4d20f2f", x"6842d4fa1daccc2e", x"bdcd1b0e7796f133", x"9dbe0647a46482ae", x"269599b4acbad555", x"756339b85268ca77");
            when 873612 => data <= (x"6968d5777bc4b045", x"c766f4052aeda62b", x"999c5684826aef09", x"fc401c221fe021f5", x"13cbb8c120268cce", x"09845c3f3da9867a", x"d6720065549363c4", x"30864355ed5d6043");
            when 19003517 => data <= (x"91f08c1957fc1227", x"37697a8bfef11078", x"3bb9d045d9da2267", x"c755273349e7d722", x"0033692b4672046e", x"044cc4b5dc18c439", x"43fb625b1cb17d4e", x"75a3536daac82b7a");
            when 9491307 => data <= (x"465d1aafa8211162", x"0d8b7bf6cc6fec23", x"6c5234b3463332c9", x"9e498f9157825ad8", x"0a74b9700c80b3ef", x"8a243ac91d95a592", x"e2bff7684dc3719b", x"2ccf4af6c1c0dd5f");
            when 14709581 => data <= (x"0b4734b61952c56a", x"03d097774271f162", x"c4427457bc591b41", x"15fbeefc0f983a37", x"8631e2ea831088fe", x"917440fb55803ca2", x"660fa64a5ad373fb", x"99190a2d54c72e13");
            when 16243810 => data <= (x"63cf3fd522285b45", x"c0a54b34f3eb24f6", x"a26a47475e4560e8", x"d6635146e100c664", x"5d26e79ad52e9123", x"e4db9c20f6f62bf3", x"c8d1eae8d2ca7f9a", x"48fe02888012e3b8");
            when 17925208 => data <= (x"53a05fe9fc18e429", x"856a8471dee56309", x"3277e55ec2143a73", x"46fd5e940d2f2c64", x"47daf463e61f3ffd", x"06f52007f6ff4ba8", x"f96e8856870cd268", x"c952ec9cf6df9ec1");
            when 5894065 => data <= (x"6728c03efe146106", x"b0e862b854a89ee6", x"3fe54d469aabab55", x"90cbc9b436398ee8", x"57cbb8f2df7c81f9", x"d69ce5401302cd8d", x"129f61fe90f62885", x"3354ead4af37b824");
            when 8319614 => data <= (x"ea1ae6f92f74428e", x"b0939fb982bcf988", x"40c826d9a08728a8", x"3ec5d09de566b5a0", x"45aecc51361a4392", x"709e3b6b9a5540de", x"5be5e8c9b61a8e53", x"836a0f7140e1ce64");
            when 33441258 => data <= (x"5315262c293c3eb2", x"fb2ac6d1d4dffb80", x"21a693773ca37131", x"d7b37b54f8978deb", x"de771236f2ff9e64", x"17818741d3766656", x"e98c45e8c6ee408b", x"946aee8bf039ccb3");
            when 26453283 => data <= (x"8850a24a84bfcb6e", x"28f321329b4aaf69", x"0f801d9adba8f646", x"fdbdbb72f2a81768", x"cacbd4773f67a2b0", x"bb16bbb98e378d4c", x"03ebb7b8a3fce2a9", x"a0c0d3d9a1536942");
            when 33750487 => data <= (x"8716002e5acfd2f3", x"712fabee9cc3f4e3", x"84c70eca7cd32209", x"4663637f9bc8d156", x"76a3156d56cf9719", x"e7ecd4a668b47e68", x"930ba9bf6a3ec4f8", x"8462b94e194c085c");
            when 14757088 => data <= (x"1cf086ac4a6813f6", x"3bd3eebe2b4c76e7", x"0858e7f7870bba4c", x"03ff4b64950edacc", x"57f50ba9d880234f", x"0ba686770265dbc8", x"bab1eb281aabf4b1", x"11da0c454ba9e2e3");
            when 28398968 => data <= (x"4456e8c6904d4e03", x"e53da3c2fc95edf4", x"890fbb6530fc852f", x"9865adab8d5eab7a", x"c45634ce81bfeb12", x"1ec3c2cb7442c268", x"5953673e9eed9649", x"7b8ae93c855979f4");
            when 5855505 => data <= (x"4c79f09d48d020fb", x"f34c7bc8a08be254", x"38c90887d03ab978", x"5654290dfe4302c3", x"786a158a21f4e358", x"0b40e5eb2fa1959a", x"08498782b9bd4b11", x"1a68008d94b3da0b");
            when 1431505 => data <= (x"bda0c8b000cbb845", x"7ad91f9c7cd334ea", x"f1fdd45ace1641da", x"56c7230ffe13e035", x"824d6bd17597e190", x"4f8b6425002c0487", x"1d00fe40eb732a0b", x"0e6762e10bc1cb85");
            when 22888620 => data <= (x"8d8a60ba7df21021", x"7e684fb90e3a44de", x"7c7813adaf107bd2", x"0f6a31255fd6487b", x"9fb638b55acd0b0a", x"2b668355a059d5fa", x"545d5bb4383f051e", x"5b106ca0bb4d32c4");
            when 4765221 => data <= (x"006c05b4e7f8f3a6", x"9f9bfc8eb54e4bbc", x"51bb57ba16b52681", x"6ab34a1ea1467c5e", x"fa307ca6d83f6382", x"981b6afb511a9034", x"80d524aabf9166fa", x"05753659a763c4e6");
            when 23721753 => data <= (x"f1a85b299ef86341", x"7af261c400fe7f4a", x"8f3555a6b895aa82", x"75c651d10bc433d6", x"aefeeaf39891ac35", x"c8515b2f7a351508", x"94e3450644c61a06", x"ff224ac25bf972dc");
            when 5628109 => data <= (x"5684ecc58433f283", x"751f6e01a1c18612", x"85844579773b2167", x"5250d8510f14d32c", x"189b43f9aeb4c7b3", x"b7f9f3653b692a8c", x"f3630ee220aa97a1", x"6f553a2d42468825");
            when 18456307 => data <= (x"5dc7409585188f66", x"f8d1d51537bd2302", x"fe901f18b8a4fda3", x"516d5aab4a22d9c0", x"cd6924cc0d933fe2", x"608a63fd51fd6731", x"83ae3198ab2d41bc", x"54563b77cb7119a4");
            when 8723930 => data <= (x"96816d4d8c070ebe", x"95a5ae077fa39f7b", x"c4c4313cb978ed9c", x"e30f5515c67c4829", x"b8ec2f7343ddfded", x"16f69d1b36d1a7cf", x"a6767fb39144a7f3", x"f360a6a99051dbd1");
            when 12486258 => data <= (x"c8acf199f3945203", x"a1c777c6c654c0a0", x"f26ad66d09e02c8a", x"c862f029c86768df", x"8d208fb97b45ce3a", x"a9d6a5a7128d4694", x"0b4ba9610c66453f", x"48f45ed0ee4a18c8");
            when 8145355 => data <= (x"feac4a597350b7c1", x"ef048bdce910c7fb", x"d7b7c5a3fa68dbe5", x"422c51415a4a8081", x"ad86ca4fc8f78af2", x"d011df71f047ef17", x"c9b5f72cb6575224", x"09f005e0b57757b6");
            when 20145347 => data <= (x"b6503a8d99813208", x"8b0776ad72669860", x"733a0a741d062ef3", x"d80b8db98699031b", x"dd81b5a4eba30e9b", x"6a982d8618ae2ba4", x"4b0b08cc3b0ea3fc", x"8d4ea5a4483cd27c");
            when 21545647 => data <= (x"82712cda70334f78", x"cc05000b469ec1e5", x"5e0f3e0b36b35f2b", x"2aa10d81a946502e", x"1e142382628a7318", x"4479d8c041a453c6", x"5ad45ce8c75e1874", x"3187314027244beb");
            when 8313179 => data <= (x"3a177766dce741e1", x"09ce841b81fb8a18", x"b3bb8e1fc1fc81c1", x"481fe8ead0219cfb", x"2ecdcd12050716b8", x"93e5aee40941faf7", x"838dcdfab502b256", x"9730abb6ce775785");
            when 23055007 => data <= (x"dc971966d494dab6", x"bde6426b4d889ee3", x"b3a15411a694ca79", x"9693a4908faf6c39", x"08f87ee8b9d38c6f", x"693952aa066fc600", x"f10c6caa9e883885", x"570dbb6906a5122d");
            when 24367472 => data <= (x"043908d41f549499", x"b8be234ad73dcea4", x"bc269eecaf044e8e", x"d1038df15f73def7", x"0abf6fb62f3f9bfc", x"875157f21b03672c", x"eea7c0af9c4203d8", x"206502896878a356");
            when 14114269 => data <= (x"bae4b1f6b256e248", x"a9872918a07622cf", x"f1c61a2baf8e1f10", x"e30ec7eb1443d690", x"94d087da314cff55", x"ad3f2226204b69b5", x"44a863aec695be80", x"27602b0b1c7c1949");
            when 15745252 => data <= (x"fcc3a16cc6f5bbce", x"a6818e86ad6498de", x"38a4203d5e3788e4", x"eeac1bbe87d09ce0", x"4ac873a7c2f0bb1c", x"ac6e7192373df758", x"8934b00bc0bcc203", x"0b1c232d35bb8e5d");
            when 13099921 => data <= (x"834a02c1694e850c", x"27f4e9b0bf170a46", x"3c2213a36014b79a", x"57ee7fbb4ea94270", x"56c1e29cf6a57df2", x"e258d92976ae8ec2", x"effac49f4cd64431", x"90a2abd7a691fb1a");
            when 3244615 => data <= (x"2c2a2df19af5795c", x"30413984f610050b", x"1b0cbf59f62b1fa7", x"b11601a7c33ac6a4", x"9ec8d4a8a3b8807d", x"836ae6bf876544b6", x"0ac45d737eca0ff6", x"260d5a497b25f7c2");
            when 24063722 => data <= (x"04561f878463c7fc", x"6ee6e828706545d2", x"0504d2c0fb81dcea", x"2a4f1a48a3d83d26", x"a50d2a5e63290ec1", x"b8524d52b2663b1a", x"3061f9c44c656832", x"eff81cdfbb7eb688");
            when 28534061 => data <= (x"b766b68d6b6c92d7", x"996ac140614cbd0d", x"957e095bb1c483ca", x"0be66493884d8724", x"7619a10ae6bc49fc", x"b63ea9a0678058ea", x"ff3563003e575241", x"a673927f5a82ecc6");
            when 31094640 => data <= (x"944f451dc52069f2", x"1ebd8f6d16eb461f", x"a5e20935ab967223", x"d05d0a28072c876c", x"2a0fc5ef56cec86c", x"75933cb9ffabdc93", x"db08ae24989429ba", x"ce2489325d41190b");
            when 26264932 => data <= (x"08c88ba5406886b2", x"4c3bec90d7337b06", x"8588f46029bd9539", x"2325f8815644b6b8", x"e25153f44f18be73", x"9111dd819ebfe65f", x"9c5362dc42168123", x"4e62273c8e43230a");
            when 25864277 => data <= (x"72193784f02ff055", x"01b1e93e3bf5e847", x"87bea1a5b764b0f8", x"d257e3177fd7d214", x"67c616085b7ac1e8", x"6dab9389332c0cd0", x"70d1e5bf7ab2431c", x"be4aae40a0dfcde6");
            when 22762355 => data <= (x"bc834c0c0ac405f6", x"c467c39d9e30402f", x"868e3453e551932d", x"1581f352225bd6f8", x"03962580e3de1345", x"39f7af06cb46e07b", x"21850d122f42675c", x"7bc165dd08ecc99b");
            when 20721732 => data <= (x"b5243cb60e1ed1c3", x"5b01c6de6ad50f3e", x"156233f718b2e678", x"96f51e3ac7e41d52", x"0f7db8a98c62d1cf", x"b3d3315650ee92fe", x"785baafce647f528", x"0632248991d0a406");
            when 27756503 => data <= (x"de003a477e4190b4", x"de08afaf579e7c81", x"1f333844bf5d660d", x"72853aa7e9211f5e", x"22b6b213c408224f", x"8d893597f987e065", x"14746c8c49f44a9b", x"3b6b1a646affdb66");
            when 1240034 => data <= (x"321e28690cf15a2a", x"c6176377ad303def", x"223b30d13c4c6942", x"60481deccdcc5d66", x"a0b5334222009bcd", x"0fba50556f777196", x"cf2b46bbec0a2d7b", x"2cdd210eb1b4744b");
            when 5617573 => data <= (x"741ff8b7defe0dc4", x"5c98c8dab1ead6e5", x"a4e7a0191d61e5e2", x"60aaf4221815f73c", x"8c1448f421960126", x"94f4781dfde2c0b8", x"fad88312c347662b", x"7758fcc32b0b61c9");
            when 20547535 => data <= (x"6088991e97088455", x"35b09d79e5d3bffd", x"8aae0ad62b1ad772", x"ebcdb63558d4dc00", x"7bdb5104df32a299", x"4a6876b8c0aecdb8", x"fbd2b3856560fc26", x"136c34b19f48c96e");
            when 16984351 => data <= (x"a45f4e5d02490050", x"8d29fd5071969152", x"244e788b37990607", x"da9c125208473171", x"24c5e830402f9921", x"e27bcb58c7f994cf", x"3341b238ff736592", x"7283256f8cb55017");
            when 6832168 => data <= (x"11856c119121b442", x"ff2b373c02f9926a", x"3d4faca7642c5c79", x"d61dd6dfdda44b3b", x"da01f2a879a63fff", x"8d9fee540895e1da", x"a83ebc79b3355341", x"362098fa5adcc36b");
            when 3695231 => data <= (x"cc20a2f44628007b", x"d612aa234b2b0444", x"ce071433d302217f", x"b4fee435eaacc2ed", x"2c05acbcb23bb29e", x"a80b6264e920cdf8", x"f0b57ee472c56b14", x"d3629ad27e32da65");
            when 809007 => data <= (x"0a7299eaf13050e2", x"b7ddcc47a254149d", x"66faa94e8250620f", x"3b999534cb4afccf", x"a4eaad847f7bd60d", x"b4c3b780425ddb1f", x"42ccd573322ea2af", x"302c752222f3ce5b");
            when 26210815 => data <= (x"06ff15e9275bf704", x"8c61de769537f1f1", x"4f3e8e0f7385ab18", x"58e8901cca7aa0d9", x"993c90320a1ba6d1", x"665a3f457caf2cb4", x"0feed2021d313189", x"a6388b1a44bbd7f3");
            when 13531547 => data <= (x"d05bdc2ada6f35ff", x"d1f3a09f770afa79", x"75f06280c1a52e36", x"a6d3fe1360944a97", x"65dfeb3648559bab", x"2cedf3704dfc8921", x"ecc393616f53e56f", x"e617d8780ffdf5dd");
            when 11468782 => data <= (x"9f6445f37f81d4d7", x"8041413af7e56024", x"e6e670618df37fae", x"cb6f440cfc081b66", x"0289fe4990987b61", x"94fd1375046e7014", x"592d748af104f054", x"ab152ec98215c202");
            when 1938809 => data <= (x"1fefb76c6f76187e", x"c70827c4c905ea39", x"d9c88110cded3c5a", x"fee475f8f6ef75e0", x"55161bc87f691b0d", x"c1c4494cf9afee76", x"bfa26d024f721192", x"159358628ab18f67");
            when 24558000 => data <= (x"f9295b3acb9c0601", x"34babed6914c5dc9", x"3d6cff91282f52f6", x"9bc66f03995c6373", x"9df527cbe11bf321", x"2a65200ab0add710", x"8f92b907d9186e7b", x"2d5f4773cce94819");
            when 4618370 => data <= (x"c2f238db2dd9cf44", x"b0499d5cb5d6c6ec", x"66496f3e4fef5303", x"7fa80527f2d24e10", x"013acc1613436892", x"980a8fb0a78e89fe", x"0b49492b6a302571", x"b48426234b6c9197");
            when 30548003 => data <= (x"97db2d423f7d00c5", x"77e662383b771f43", x"c76ede30e4c09c91", x"88fae792dd49aad6", x"6e08649d162b1939", x"148a0c9d9475ecac", x"6a4273d518ef3964", x"2dd4a769380ce9b2");
            when 8393844 => data <= (x"eb6219732907b540", x"906122d76dcf7a9e", x"8e82086c30285ef0", x"1a3525728ff316d3", x"ec6874479d0488fb", x"af78f44bc6e29bec", x"1b09949a241261e2", x"0995a74f6a3e497b");
            when 6019395 => data <= (x"3eb6c219a400e030", x"f952d785326f0046", x"d2ed288208fd064e", x"403d72e713c932c1", x"df26536519846f2f", x"5f76840e8c7735e5", x"a745e937ff9029d9", x"dc19a5b5d1042479");
            when 30760203 => data <= (x"7ceb93a6c519e061", x"0310d889de1dee57", x"642df5e64d1001c5", x"b271ab5acbcee9a9", x"4989d1b6da746f7d", x"6af040f06575a046", x"602d2ce5d6ed55e4", x"7f7459ea2a2b2208");
            when 19097587 => data <= (x"b57b7f8d08130fd5", x"dab7b25eebd248ea", x"11b33d387dec9ee3", x"4407db2b2f03db9c", x"e59fc3ea8e203bc8", x"7451d98a0bf83334", x"4d526dd99be52201", x"2514f24bc9c0f67d");
            when 1587209 => data <= (x"96bc3bf412e38cfd", x"2f30d84f63f938d3", x"c91791b4c3d83758", x"78130728fc01faf8", x"de0f69af18b36b12", x"6bbbbabf5899e53c", x"ec454229e05170eb", x"1aca9451155d1263");
            when 31453405 => data <= (x"3f388f49f7974289", x"08d755dad27162c9", x"55d69237b5d8ca7a", x"b16ea16d76d0f3a4", x"8addfb4abf71bd94", x"4feb3fe071e7bb91", x"476c5ac40272d4bc", x"2d504e999871b58a");
            when 12428912 => data <= (x"eda71ddfb3478316", x"e2d4c19d1b3805f0", x"a20a461405e8312b", x"9cf5b9a6da6ee4a8", x"f864bdc456f8e771", x"eb9c39e455923041", x"6267496d73eaaf10", x"617c0ee1213e8523");
            when 8127857 => data <= (x"76166fa7d1067de6", x"8cfaedb6e07d251b", x"e156cdc29f0333ec", x"0d9f31b3593e31f8", x"d1571496e7f3fbc6", x"8c760a29ced9308e", x"70a926636baf5485", x"cf3923d4bdc6ade9");
            when 33159840 => data <= (x"0e80b00fe5946d3f", x"efa5a5738bc111bf", x"8a8fb78589a83065", x"3cb64a12c25f487c", x"45dbacac44c2f51b", x"be6b307802920e31", x"1c0b21be34aec7db", x"83981cec3f0aeb68");
            when 6689035 => data <= (x"8ab94c18cbc237bd", x"919c4aa21eeb66f1", x"010e2b76f08d83b7", x"49a29b4ae7b73547", x"c1526d4a97079220", x"5090f4627b621866", x"b658b3de3f56124c", x"1e84a815916a0a04");
            when 31574557 => data <= (x"b6fb0bbf3945f527", x"50f17a7dbfd66b9f", x"3467cb805f4e9eba", x"68e0ee6b4137c518", x"b218bef4f0987176", x"72a53e9c8695168e", x"2cd0fdd0bbdba68a", x"5dc054312be13e51");
            when 18360505 => data <= (x"62f978f802dd4aa6", x"66dd01a6fe191b7d", x"bfdc1a54880d4cba", x"6d4fdeb4cf1ba46d", x"08bd2ece45203539", x"bb2e8463b5f1c170", x"ef1db7e50a41cb5b", x"01bb0b951b11fbcb");
            when 15169588 => data <= (x"ed98a4777637ef37", x"8a59432a4283834a", x"85faa3b13602b6bc", x"ed3869095676806a", x"90b52668381cbeed", x"508a9ba02b054b51", x"c6375417a3fa1d9c", x"947a0bb4da67a74e");
            when 22753987 => data <= (x"746daec8feb7d18b", x"943104b760b138cc", x"e10cbc3cf46aa29f", x"4b1f7a0c7510a638", x"8e6d0a826cade573", x"c2a545fe88559d99", x"acbb8e0ea175b3b5", x"54e6d79e057c954a");
            when 12664712 => data <= (x"ac07cfe3c8c54525", x"2f1aba7eecbef1cf", x"3b611617bf5c11fa", x"0b09413450f96e98", x"a8685f110cc698dc", x"70d0270f2cf22c22", x"aed145a43ed40691", x"3b223c3d2c23068b");
            when 26831916 => data <= (x"df7552538e97f46c", x"71aac8e404e51e4d", x"86649ce21edf4c07", x"e6b1855ff167b05c", x"9debffd1bddaed45", x"a7f9ac8823dd1432", x"c6f5bcf1dedcdedb", x"b02d824403dbf24a");
            when 14716410 => data <= (x"cacecb5a375e2e57", x"49cc865025975b63", x"dc0aa8f50c7b073a", x"edcf9adf46b188f6", x"f223c9e22be665c9", x"53b4d689f4ff8526", x"662df2f757ca7c62", x"cebe2795d7a532cb");
            when 24217294 => data <= (x"1eee378916ea7b99", x"f692a2e6bb8a6e53", x"4ebbe257ca44a860", x"a5af228f8083cc65", x"44ec645d42602e6f", x"842d2823f5f32e4d", x"7d6ef4dd394b871e", x"cf9a4371b090b30f");
            when 1812069 => data <= (x"96776a8adb10e214", x"b1bf0cd2a0cad945", x"a38b74deece5bbf6", x"1471d86e417692c9", x"0724e92e82d0fcf8", x"21cf01f57b6f427b", x"278f7bfb3881003c", x"a889d407ef1cb4d1");
            when 22085898 => data <= (x"7b88ac21e120a0eb", x"76d7304b42b01fcd", x"85e23a88efe2f47f", x"3ee9326c3969d453", x"fdddb2a69cac4477", x"398d515a6ae955a6", x"ba6005918fb1b1eb", x"bd013ee5a680570a");
            when 23082425 => data <= (x"111c7bfbc4b2874b", x"ea55fc44b9f73c8e", x"250bb01eef8f3b9c", x"e4dc1f0fad8fed80", x"5daca586281c29d2", x"5a94016630761e5c", x"d1427e096ae85fbf", x"0cb5628cb7d76336");
            when 23394650 => data <= (x"31d2e519fc284cb5", x"8eb153e909e32576", x"2bb184ee83b733c3", x"beed24c1246b5648", x"bcfeb0aeae0d6f20", x"7a4a39874e651b77", x"ff2ed5d8b3ed83d0", x"d4924e8d421aef3a");
            when 20833444 => data <= (x"4bdc24a9aa24ed19", x"e2cd35a0c2e50387", x"1e04568e6e9ab58d", x"78e240aabeb14751", x"5a1977f457f52e3c", x"3faa4efa8e3a31ac", x"0b9fe221ec84685a", x"f5b88d849d510fc1");
            when 25047600 => data <= (x"461268567baffef5", x"adf21972fad4eda8", x"444264f80d56b8f3", x"6e3ed69bb79432f6", x"04e5a8ec19b56a07", x"f13e8796368d581c", x"97b4b840fed62012", x"a04f723c31aa160f");
            when 26301367 => data <= (x"f4add5a22b9b29f7", x"3120b49dbc0b4cf2", x"b16e3d982824fb7a", x"0df55bea0b6c1856", x"e993f5eec423fe95", x"3f66b41337b9e924", x"055956213234300c", x"daf64c8b44e18a0a");
            when 7313806 => data <= (x"c1327f520f32d6d8", x"3eb3178c9928b0f1", x"b09fbf0df60b8c10", x"6c705795474c6b18", x"398bca6c0b38d230", x"f74b6c670d0583f7", x"b9032baadff17828", x"daabd886ef2d0acc");
            when 29960066 => data <= (x"1ba290a179f81e11", x"2a5391ec805e72e5", x"c2d9ba12792c22e3", x"c1943b27d3a1091f", x"ff5535a884402f07", x"22de3b579f1ba59e", x"90d9cd0bc1bbf3b0", x"51f2a63a3ca2a6b3");
            when 30659014 => data <= (x"2870a65d9a75fe01", x"2d4e5948be5354ea", x"ff4b09dc040f5bd2", x"0b2f934c25fbf771", x"2c77fd9e71cb0287", x"33f04079d5659c9e", x"faeb3b8d4540c010", x"eb9fae270551accc");
            when 13609936 => data <= (x"d522546935c840cd", x"8019570913616f58", x"1e2a3f9e007cbb7c", x"337397dab07a83bb", x"8a807945a87e950b", x"1a013a1197f0a642", x"e4c20d5e32a12370", x"69864e817d1b9f00");
            when 22858884 => data <= (x"2abba678b0a93630", x"535a073356a430a1", x"db70b825d10fb4ff", x"b05152cbd4f341c4", x"38596c9ca2c508c2", x"ffb1dd516117632a", x"9d4301eb7a86e6b7", x"1249970673e221a9");
            when 29593784 => data <= (x"849d33160642749f", x"9a3fd6e579454e64", x"f857c52a2e97d3e5", x"006fbe6fa7001817", x"026c14454a4d8633", x"376796ff4b1be446", x"e11a5528d3243cb6", x"d2c2f43f586a73cb");
            when 29419351 => data <= (x"89c4194b53ab0b65", x"3eacee2203b09a9d", x"ebc4775acb347a68", x"32db0ea2ebcee3d2", x"a23136ff7ddd7ed4", x"0ab18d79f000156d", x"944d407dd020d464", x"d79354265821955a");
            when 32635757 => data <= (x"cc70f8a51b25547e", x"523aad5667f8b33c", x"78357a392f1553c1", x"857d4f1b40902f87", x"916501a1e62c8c28", x"676c1d5d0860d4ff", x"7b70f65ea775a39e", x"77f40203fc73d80a");
            when 2433182 => data <= (x"f7d14690361a761d", x"cd5b84bdd202f47b", x"9ac1a32558b95c12", x"8b99717edb290d06", x"0494ec8a9fe5b990", x"71447cc22fd8eb70", x"a8cf027d14bbfd0b", x"a0af4f661a4408c1");
            when 6946425 => data <= (x"ca0508930694bd22", x"0d60c15789eae900", x"45d500d127bea26f", x"4198506cb8d92829", x"b85ae3f90ff5782f", x"daf1512eb99419c1", x"86a70b10160f3508", x"9ee75336f9b1f45c");
            when 615636 => data <= (x"7e94ca4e8709ca39", x"31f11aa82fcff863", x"40520ab7a0dea2f6", x"70f1580b440fda0b", x"8e63f468d6fcb738", x"59aeba81befb8790", x"df91b7eba3fdef48", x"d8432b9243a35560");
            when 2672725 => data <= (x"1a1a29237aebfc94", x"05a84f4d2f12a3cc", x"78ead2fca5828d5a", x"4680f551e3312ac7", x"a518cbb948ca1e6b", x"7dbc5d170980f8fe", x"ab27c1a817c7d5b7", x"d3a8402a3ce408ae");
            when 8920001 => data <= (x"74572962599248e9", x"0e4c9b8d45489d75", x"29a64744ecc0d2fa", x"7171a35cb1b277e9", x"86389e226abb01eb", x"e4560d72518f259f", x"5e04cd24a92b4614", x"95d56e5ab02ae3b1");
            when 13045657 => data <= (x"4617892593708065", x"8802ab574574bf7e", x"4d75ce2dc153df7a", x"e18dad50f59c9247", x"2c3e3385a24ec0dc", x"56046d31f16eb4f4", x"4c9081122dfa065b", x"21c1fa6ed48b77d1");
            when 20059933 => data <= (x"4e5314630e9a4d07", x"98fd5cbd8ebf6474", x"cc5cb7c9797540b3", x"41a594fd02942a04", x"0bc8e7faf2b8be7f", x"3f0a87d763c27307", x"6e052202b2e20e23", x"332f6ec359e38dc3");
            when 20260020 => data <= (x"e1b635d3b7d1f565", x"33f4d2bf17e03595", x"869cca2fd1c6e768", x"2fb2bb3ba01c7d1a", x"5c67ce5b95ffba32", x"8b93e373dedec683", x"035a21439808b1ce", x"36af7b59343140bb");
            when 20274798 => data <= (x"8bceedd1ac556d33", x"0b32c4b62ce96fbf", x"72c983de633c7325", x"c6d121f44ee61e14", x"076a697b77a19b63", x"7c9180cf9238a81b", x"2b6856954bf9aa17", x"22da5478f4a7ca20");
            when 30685312 => data <= (x"ebabaa53f7c4223d", x"55a10c835e908f24", x"0d391e3d2858fe63", x"cc203784d3d8ffe9", x"51266a22f135f82e", x"054cf24403bac9e0", x"9d37bd2d95dadc77", x"9af5334bd955f6a9");
            when 25561505 => data <= (x"6cb14f7e5dfada76", x"f43ca7f65c82acaf", x"7cc6e606308da8a8", x"880a1c043bd48b35", x"c3fca3125e2d49ce", x"5481ab6f9deae6c4", x"cb36638644c554c7", x"fbd9cdbbb0d4f9f5");
            when 31935992 => data <= (x"3a9f1c116f2030fa", x"b58d1c932b001363", x"eddc6b454b0e85c7", x"679aca6b9b193c66", x"7afb4290ce826770", x"c2f44156745cba82", x"a95d9d7f755179be", x"f3709e005741da78");
            when 24137668 => data <= (x"dfb8b9cb0dece1e3", x"23ebac285bd750ea", x"b9e6f29c670dfb5e", x"124d6093263f1957", x"3fb8eb01418480e4", x"17e082144b01dae1", x"52e731993db9c8fb", x"022b13d54e2cbdeb");
            when 17095619 => data <= (x"fe99bdd43f8bdfdf", x"bd68514c74f13c33", x"62d448df82012c7b", x"f5ad6fa90c86debf", x"f4315eebe2c88bc0", x"407c11f38b00a712", x"2f57281e6f4b3fc8", x"f12a3d9ec37546b1");
            when 32472626 => data <= (x"e66de86bc96daf28", x"c63b4b968fceb668", x"3f3ef0753595d436", x"3099720b25fcb091", x"82edbd6b664593b7", x"caa98ce88609a482", x"4a99f9175c22e6c9", x"108a6420f9a2eb66");
            when 11059473 => data <= (x"76ef27701a3436c0", x"0ea22fcf186ff6ea", x"eec467ba30b1def0", x"f7c37fe7d61dde9d", x"0b92dd8bbfc93cb4", x"42c255c546809733", x"ac76a3eea8dd6477", x"09862c85ee3f2fd4");
            when 23239005 => data <= (x"1cfbe429ce794b6e", x"5cb9c2ddfeed594b", x"742a3626d87e240d", x"391e764cd2b640fd", x"ba2ec1dd409fff0c", x"761beff9e7d01aad", x"fa7fb9e9b6d88a81", x"bc564ef7bc5581be");
            when 2348350 => data <= (x"df2e9865b266c70c", x"7e0189d2df77ee1e", x"b629034fc2d7a907", x"cd5ee8aca32103cc", x"28edc8ae69eeb8e0", x"dc88697f1587dbfc", x"5b9d5642748120e8", x"37ff98440d8dc45c");
            when 19709126 => data <= (x"f5d2726d4d3ff886", x"c130b11aaac401d2", x"c6e85158a916dad7", x"2de4ebd0cf8b4456", x"7ab776ad7a3f3a3f", x"3b28ddb91fb7bab8", x"41502e7faab0e61f", x"5ff2ec807cfdf120");
            when 5572961 => data <= (x"7a08cf386ed4a1cb", x"7e209f212f8b97e6", x"537c3473f3bb46df", x"42df8d698d46e21b", x"4c6ec8ca21330a51", x"1f1f7dac7c3b13e0", x"5e6dea01240a5423", x"f91212e1aa5789bd");
            when 8435150 => data <= (x"5ee33038b4c4678f", x"c5c1d40b86fff348", x"d1534c699255a154", x"492e395bb64f3a13", x"ef281bae443dae6f", x"1d425d34f25e8b5a", x"53b40e01714a9ddd", x"000a3d6c4363555c");
            when 33578494 => data <= (x"cbe2408d614460d3", x"43ff990ca202ccef", x"beea84c3afa0305e", x"b403297e684b088d", x"aef0834c13daeaad", x"9218df23588d0764", x"9b81774f3b11d2cc", x"08e47831f0a342af");
            when 13338091 => data <= (x"ed2145074c253a75", x"f0c248b14183acba", x"4a9686f542c99b0a", x"60bc0280f6a71df2", x"18fbbb793e4417f6", x"54f5319267edbe1f", x"af42a410bf3a163b", x"3679a7f7e0b08cc6");
            when 24987203 => data <= (x"329517b0a693c9cf", x"42701f52346cd6a3", x"e32b294bd5d5eede", x"a01da8c957f55e2c", x"1b8737a6a91e779f", x"daeed650373503df", x"537c1831b462738c", x"1ff9d923fcca9f31");
            when 15356843 => data <= (x"780a3007d007c61e", x"fa592e52cfb2c9bb", x"25e3148c360a37e9", x"423ecdc31d8ad560", x"103b3ddf3c980e21", x"87f77fefa45856a6", x"09daf6a5e5d1c363", x"4b9039d0af0bed11");
            when 2488801 => data <= (x"109a60f0d70eb308", x"373a0c66a460f8ba", x"c552006136f8b09f", x"aeaa529b62ee59b2", x"703ab993d2e2fca7", x"635dc289a7cfb6d9", x"fee3e44308cc9a6e", x"3801bcc2ef0cd318");
            when 33885987 => data <= (x"0d90ea7978da70f4", x"aa5680ef4e7ecf93", x"0965ff928400aa3d", x"a835f3fd3d5af5ed", x"3bfe514072ff1fbe", x"4ce5ac78b52acd99", x"8ca9d397c0820763", x"5fd3831ea4a8f22d");
            when 18090189 => data <= (x"c6285aec34cf0f34", x"825c136df6ce9d2e", x"be3cd024f2da9655", x"2ce0e2a8b02d06cc", x"f8cd507817597227", x"70c7d4162b86d53a", x"00a14547ef6d98a1", x"80e4aef139339605");
            when 26931223 => data <= (x"3eb234956c6f74c8", x"043f78fdfd02858d", x"e151b627dc7ef2c9", x"88e7e27398ce4048", x"83e3a52388e94ccc", x"721009155f4a0f4f", x"4beb72791696fc5e", x"d3badcc94fbfbc96");
            when 26936026 => data <= (x"62345c05fdc3ec3c", x"cc5491135af0225b", x"4c85c9858990d1eb", x"cf8dd13655fae4da", x"fdb1469383630dcf", x"380b5d9d9db20b05", x"91e517a3db14baed", x"b18f3e933deec735");
            when 3584604 => data <= (x"e65e4c0705b2707c", x"b9a16081f091e861", x"e8e63c1cf3a8ca04", x"4de8fc68b4067217", x"b4cb6cc36e90fa3d", x"cfd2e51027d9aadc", x"e521461dc67539cf", x"8a6763e84660f949");
            when 6542521 => data <= (x"54f6cf22f7751eab", x"c088858a7e974f15", x"3645241afcabcaac", x"1cdab4af2187444a", x"b5340cf8380cdb5d", x"2fc8cf6532d4b604", x"4e81e1206f771fbf", x"2c42072fac4b61df");
            when 23617487 => data <= (x"1444130b5a1d42e8", x"efd06afb18f327ec", x"4195e70a63d10228", x"7d872a681f347e4a", x"dbe4ac083aba8f15", x"69543b66f54f0f82", x"440f1b95ab397a15", x"daa1ae62d593c4f2");
            when 33656330 => data <= (x"630b767ef58bed59", x"8652d2aeea0f2c92", x"14d9cf2084d52428", x"4959389868a53f38", x"52a35f46683f7891", x"8828653b0c4821dc", x"c2eba04e78c894e8", x"bd3036b7f18b729b");
            when 9188952 => data <= (x"8d103e0cdef7b776", x"ac85b7680f864aae", x"d29531b19e608f10", x"78212b23dc86b651", x"d57cc4662a439cb0", x"08e588d2d2179f6f", x"1f22b5b7db784ada", x"42610b56f3afbf55");
            when 18472206 => data <= (x"47c8200374c31e11", x"5a5885b0d186c9b7", x"54e5fd8aae6c9c35", x"b9624c4b20f65a7d", x"81eefc4b3388de00", x"c1fec8e9b362d651", x"086a233dbf80460f", x"de8355f637d3d499");
            when 29220323 => data <= (x"1605d27737863bc3", x"5b1401f17327fa69", x"3f845ffc087de554", x"511e526aba43e376", x"23777b7e34390a52", x"f972f9a261d256b1", x"44f228ab57c97f99", x"3ec9ce64eb1d00e7");
            when 19771647 => data <= (x"5bb4ca5d4263f3a8", x"78b5e4346492fc82", x"e07a1d3b2e5ff652", x"5f04a2285f97c898", x"57a11c67cb03c897", x"785514df3e30e200", x"069cc9c9be99b806", x"99517495d8709326");
            when 16053262 => data <= (x"73dca20dd391069b", x"fe75a8ea75087001", x"eceb184f99b0332a", x"a18eb59b1204a7a0", x"61262486deb71540", x"e5f5808a8d26ede7", x"5ae98552d509c794", x"6abaaa24885b2d88");
            when 26657012 => data <= (x"f6b3770b252be294", x"6c1955a287ed9597", x"881d21a9049892f8", x"44c39857bb0e4fb3", x"ae0f10a5946f431c", x"5a5f1b9cf64cf7a5", x"2577f81a06795ae7", x"c5ce51e8e24b1b89");
            when 11136200 => data <= (x"51711af9ee1d9894", x"27721072dc7be58f", x"3da0e0ac03776761", x"1790f83cff293aa7", x"4fb702071ec0a79e", x"c90d7ae1d04ce082", x"7b8e054c9f58657e", x"df950ae7ef7b0c1b");
            when 14559024 => data <= (x"1f7719237f746576", x"203d8f37eab49b3a", x"b89b6ee2a7eb0cce", x"fca41089cef7fb4b", x"c3a858e46f7bb58b", x"e7450b03be377048", x"c75e64785bb1b342", x"d83f0b6bc4dad62e");
            when 8287684 => data <= (x"8031746aca3927cd", x"0fda694c80156ac7", x"7b629578abbe36e5", x"a5bf599e5c350815", x"56c09b6e1d557188", x"9df251a7c4398361", x"22cb37df25a11072", x"a47dda3dfa4a58e3");
            when 31876876 => data <= (x"d11b01a5e8534979", x"a2d0e10f376b6095", x"3b157f740edfc81c", x"73eacf6facda31af", x"c0f903667ddc7c9e", x"38e30c1ac1759a45", x"996571bb6f16f57c", x"b6d80d81f490ec9e");
            when 15540854 => data <= (x"f47f97a75a4ededb", x"cd1c0ad561c7e17b", x"539056bb8c13d660", x"076a47b5a4c9b6ab", x"143755472ab3ffcf", x"a63cf9ebc248fb63", x"d06757428f84e255", x"0e44d5371de63e1a");
            when 19444407 => data <= (x"5353f07a77c6fd96", x"df03ad2360a76d7b", x"a2ef3e0bba6671a2", x"14aca97fa64de885", x"68522e54ef13af15", x"4d3bf4b626fedd4a", x"fcea2f1db6fea1d3", x"1c52b3a0969856fb");
            when 12791921 => data <= (x"bd9ab1108e6b4dce", x"6fa319ea952764e8", x"29cf1e6cb1041d58", x"1bbaa8e815813f98", x"0bf332cb57042194", x"5a75af56ea4ba8dd", x"ab192a9e15d50400", x"a1b204612c61b896");
            when 1801800 => data <= (x"abb4d1c384fd083f", x"7adfcfbc0eaff1d2", x"6325821263758c60", x"c1d637057f249461", x"2fa83f3b8d863a87", x"7de8d4581f7f65e3", x"19ea92bab72b2c77", x"81bb2c48a885aee0");
            when 3786402 => data <= (x"f976aaa9d394e114", x"a07138f759566ce2", x"4e77c5267b419033", x"1347eb52bfc1d878", x"c2ebc56ebb4942d7", x"7ae3358f6964da88", x"00d123ed781ab89b", x"7d0c3d287411ccdd");
            when 31478344 => data <= (x"675d0483c611f587", x"f5ce1832a75ed089", x"6c4d622c650131a4", x"2fe50ff993b27740", x"bb0c82d11245b753", x"f1836998ad5f54f8", x"8f5455fd9cd3f7b3", x"3119f95472bb7902");
            when 9222810 => data <= (x"40330806fefc65e2", x"8c1a1ee6d409edfb", x"56155f960ae0896f", x"a3a5f88c55c75d89", x"b21599f57de4f7de", x"97f85c7e3a507e36", x"354661ed06421e77", x"c4b83162e84f3b97");
            when 28069990 => data <= (x"15e817725e09305e", x"abd89c867a1112fc", x"df00490a44a40f96", x"9a9c15bbd06d4625", x"967afbd756273905", x"1f1ee8990ad2bf91", x"d7b0874ce6a12125", x"2b0616f74eeca2a4");
            when 7073541 => data <= (x"1d105e63ebf67e96", x"740be7a13710ad65", x"2b9282e374242539", x"22944d275a614750", x"c735bccc7dd794b7", x"dd135c0c74df58db", x"435f62b97b20b15b", x"e25f28e4cfc36ac8");
            when 12835436 => data <= (x"06699a5cd439de48", x"6e1064b252d5a3d0", x"323edd392fd786fb", x"ec4425dbe6ad3031", x"e53ac2ddbfeaba2e", x"83656f956dd87010", x"89206ac2190ac27c", x"0838f24d809919b7");
            when 2628665 => data <= (x"2e6b97d1fdd7f9f7", x"7de4e76994263b14", x"f45730ebe39bb075", x"8d3403a285c2993f", x"4188b4add77e87ce", x"fa978dbedb70c900", x"8dece317df4171e2", x"dadd25a0ebe4f87e");
            when 33298800 => data <= (x"0dab124ff7768c6c", x"518f0643c380ad50", x"b98b46106070a07f", x"e747c3d90b61b646", x"91d29e5ae04ae9a9", x"6f0a90785baa3b80", x"09682ee4bcb31fbd", x"1cd0a6b813322fd5");
            when 22539818 => data <= (x"b41cdc0d4477480f", x"809f0ac93d2838b2", x"961c9a2291c07777", x"7217c7826fc240a0", x"ae53b43e87294137", x"167ab64c28cf4726", x"5ceb578b5ca7d4e9", x"81816a2e5098e583");
            when 26274050 => data <= (x"daadf2d656bd72b5", x"ae8e0fbf3c9d70e4", x"ad4b2ba6f607bcf5", x"ee8d0096f0dfdd7f", x"655b9e6926bff8f3", x"94e304fa40597c2f", x"ed6b62812899d7a7", x"206ceb16c9faf96b");
            when 18838099 => data <= (x"a09462455cd55567", x"6ca66c7ba7b39b98", x"775560113a2a3b63", x"3fb23faa1f14cbee", x"16a54c3582ea9e6c", x"cfafed66f83245d0", x"1357c026bb2d61a0", x"8a0ff957bda9a929");
            when 3009290 => data <= (x"c48ce3d7ad40e97f", x"4da4799c3b04cac8", x"c742e93cd55a54a4", x"9d537d21fac8d826", x"861e1f5aa960c845", x"e643e342a236ec5b", x"62bf83df2e83617f", x"33b9d95a9381f623");
            when 26500428 => data <= (x"ce598c5dabc0fdb9", x"c8ba50c2262a0eb1", x"b802419943081373", x"e576c03b4864b8f9", x"863d4d5da0801c24", x"622bba19c8d51b00", x"8e5dc5525b705e3d", x"af4f7af1e485f008");
            when 15968113 => data <= (x"a8727db84f6c60a1", x"00f4afd5be354d2e", x"a7a297d758224695", x"b2000a0ed3611c02", x"ee4aaf5d2833aaec", x"7b52d3ecd042d0b0", x"5f4f1c3987160808", x"c38e3fd5f4605764");
            when 2027691 => data <= (x"bff5314bdf92ea77", x"a2d38e17631a0b9b", x"49f87950f60e151a", x"33fce19001d7795e", x"33f4bd2af2e9b7f6", x"f067d4aa39c489c3", x"73ddbc366fa5b5cb", x"8bfba3fe967d6a35");
            when 32804652 => data <= (x"ba1fd524c5b80c6d", x"6d5e544155c586fc", x"0d8a9f14610d14ee", x"1d171d1304ac7d16", x"5aaa350e5b85c299", x"8c6bfdd1ea5575df", x"6711c9d58db2ecb8", x"d45634b20358ce07");
            when 21112909 => data <= (x"77da92d654ab652c", x"9ff744869beab297", x"24847e8c1a13c90d", x"25bd52cba83929b7", x"3dd34bfbc0b8218d", x"a5f7d5a27ce3aabc", x"b9702325b47ba55b", x"548126d554377263");
            when 5559660 => data <= (x"957c6b96f2066b71", x"a3b97afa2499355e", x"1f0faf6f3930f1a6", x"2c931bc579865e2e", x"c2fb77b5d3f70a2a", x"57bc7b29960824a5", x"b85455f19ae990bd", x"79c8eee44656e668");
            when 23243987 => data <= (x"e2013d4ff4ed2c09", x"daaef5a2ff8dfef8", x"0995452f476fe7a1", x"6366b08d9158ca10", x"92e2879bb85bb559", x"ac7ab852fbe352ff", x"0cc68944ff4aa4af", x"542728c89062f189");
            when 18782196 => data <= (x"425de994b90159e0", x"2c7908ae9fb26700", x"6ce3a4bf473033ae", x"946ab0ac7e0b6454", x"78b2d5cd6822bcbc", x"8c57536ef89b74cd", x"d5d92956f6742b25", x"46d206cd47ec4a05");
            when 12783783 => data <= (x"e657932a8427d155", x"36aacfa94ea7a8e0", x"7289a5c0fd41aae8", x"c52c88b1c71e4425", x"c4ca8a49a1086f13", x"c5c098b9ec4e7797", x"7546d22f22071817", x"cb18d1c39690b393");
            when 16236979 => data <= (x"4e918756dd2e0c3c", x"a0f259648afc3d76", x"5a297819a0753b9c", x"b20b420beea70cca", x"4bda5fa45ace9ba5", x"93f33e8b6684baa0", x"a751f043f48daefc", x"7ae444636030ddd0");
            when 4645460 => data <= (x"4534b8783a72a117", x"c72bfbd6c86986a6", x"b764e59d9594b01a", x"9dc0513b12d89896", x"1687366b465f1e7e", x"0b7d63797642eba1", x"f6d3778de45385f6", x"3694ceb6a3ae5c3c");
            when 22277839 => data <= (x"138a568412b3fc61", x"c64032c04fc6eac9", x"13a01f65b453326e", x"1c01c20af7209866", x"5b5538e3717f5b80", x"5d1b6ea417e1e0fc", x"672d9854d150852a", x"2d946d874e3a77be");
            when 15240007 => data <= (x"e23c860929ae3fe2", x"5e2f8a75b9db48af", x"064240fb4ac420eb", x"185873162ad106b5", x"f79f6b1e832147f5", x"a221b15c5b675dab", x"09fc2cf632fa06dd", x"517b58d205ab16ac");
            when 19489160 => data <= (x"2cc3a33d14d79a11", x"f2c40ad4e2aa4783", x"56a87a2d18e93569", x"a146614bccb2f102", x"6048995288a5ba34", x"42e213312fbdc897", x"fe2d2c342e2086d4", x"d4d3db6f9b15f590");
            when 23080250 => data <= (x"2112f0226fe9f4e4", x"dbb592a4005ec4f2", x"9f72d0b3f24abe19", x"ab8a1c0fd274a8df", x"8350d03e086977a7", x"85b72052a7995ef0", x"d73c15303e383cd5", x"c8f6fad5292795bc");
            when 16528409 => data <= (x"562efa68c560c44e", x"afdf14bcd59d7d75", x"5cb8eef0b23b6503", x"f6388808fc1b87c4", x"df8040b7a7a546d7", x"67b7c919d181ba8d", x"6fa6144b9e2cc912", x"44f1b28ed9d68efa");
            when 24631619 => data <= (x"45f76b8552a5ddae", x"cfa8e47aff94dadc", x"74c071ea4d267d5a", x"5762852b1a7a0a37", x"6ffb64ace3d8872b", x"aafbc1c815713727", x"99a5173068296766", x"ff5e2fd3ba107548");
            when 12861967 => data <= (x"512c5476d5c80569", x"a770dd05dbf4a8da", x"c1136abc490d9b1b", x"5a11ca12e57fd503", x"43223bd4dff02cab", x"fe657e3cf98cc7fa", x"59f7c97fa75407b9", x"ba0793ebfda96e49");
            when 3443646 => data <= (x"654e3190d951b471", x"893393cf71d8e7fd", x"4e7c8acb22cb6a2f", x"23d8e2cbb4fb45d8", x"531fd371e2e2596b", x"565895b81db1cc69", x"9db502c796a321c4", x"91323eea7e2f498f");
            when 3571469 => data <= (x"e82b191b587b4ae1", x"c28a588cdc423e2f", x"c691eb7ab8277917", x"b2580cf7fa316c51", x"81385ac7c56dbf69", x"40ac05f48126a710", x"8b5b848ce4532266", x"173e2c8450bbe78b");
            when 6233009 => data <= (x"52e099d43c49431a", x"7c0e89d5cbb3ee91", x"5645019d37d3d01f", x"af25880921d31a52", x"c952f2e6494e1de4", x"50746b9db2db73a0", x"5a7915d8ae51ea7a", x"e5ae40bf58901202");
            when 26329918 => data <= (x"96e5c8ae52c415e2", x"724c0a255fdb8dc1", x"9cf23bfcb7b53e42", x"59c30b0fc5c855d4", x"f72dede7cf25aac4", x"ca18d6f43216aaf6", x"2dc42f65ff2f832a", x"e82ab028ff68d1da");
            when 10740723 => data <= (x"8c7676cae8a535b3", x"c55d08f00471d0cd", x"76133c6c2e807d47", x"33f149b79e1eb58d", x"578f5b70ba09be43", x"3b6ef8cad63a640e", x"01070b44298888f9", x"64950df7d4916659");
            when 21956184 => data <= (x"dd6aee31d33ccbe3", x"a02cac259415dd63", x"338d30b583cee568", x"514a218a95943d28", x"56df6d77ed36b018", x"5b01092f177f2580", x"8f547aa09f980e8e", x"eb5483cc431792a6");
            when 30292818 => data <= (x"15be7d1cb5f719de", x"54b28143836bd888", x"743f9a3490fb01ff", x"307422d576c5ce22", x"97ac778239773f30", x"74a055269354ba1f", x"597385c2a1084a5d", x"6ffc3c6478e8090a");
            when 29947658 => data <= (x"0292879944cc64fa", x"1b01e97af5d7900c", x"26ae2117a06175d2", x"40efed5b215d19cb", x"057adf9528c0c7d1", x"08fa74b4dde4cb0d", x"730b66985d7f4c3b", x"bad05684a19b546c");
            when 8234166 => data <= (x"ad56c0213a3a6032", x"4b78cb6d9ab6e72c", x"01694f33a852c465", x"5018a5cfee2e0fdf", x"e2a96a8405814469", x"21f3ccd3d37203e1", x"ebb13127e613db9e", x"dccd239fa8d7223f");
            when 15951730 => data <= (x"d752148dfb103d95", x"472fef70862193ef", x"bd601b38c944ee19", x"2f14b00d4b3bb1ea", x"4fad60e4239339cb", x"0a1aac8d06198a11", x"bc37ff228c93c7f2", x"8373146fe84f6e0b");
            when 20335215 => data <= (x"7074d7641cf77ca9", x"b745023887eff80f", x"f32fcee64c24be29", x"d119faaf504ecd35", x"ad1471a444ca87a6", x"5d5f9e441f0f0df0", x"86f3d99d9ed3b6b4", x"0f00acfe22179616");
            when 30411626 => data <= (x"7bb46dfdae9e327e", x"7b77fdf86dfb7897", x"c92ccdde164175ae", x"0175f03b56a44edc", x"77f4cfcaff3ecf7b", x"ca12bed3bab564d0", x"bfbf7adc204ac45e", x"8381eae375c6b23c");
            when 24501997 => data <= (x"581844608fb0dc93", x"2dcac8544f92176b", x"58268748f945c24a", x"949625e2da3453a1", x"c7055a4e7424c659", x"58ae0f36ebcb7b65", x"39965f59c8df5697", x"44cd4c9fadfed47b");
            when 5799131 => data <= (x"d516d8cf4fc5bddb", x"3b903042007b48da", x"6a8795e2c6864505", x"402dcea04e6f2d28", x"3baa3828dbbf6443", x"3432d6943a41c559", x"458874fbe7d93a25", x"a54d521221d77054");
            when 24574470 => data <= (x"630b2f57bd645d55", x"4b03daeea3041223", x"c40102c9ff8dfa75", x"0f382ffd8ac4794b", x"a80c7dd32dccf8e4", x"329a70e7d3166ef9", x"5e04bfdfc41c9917", x"c31430d4dc8e9e71");
            when 33741724 => data <= (x"d5b74055ac72eef9", x"18a84f9665d06008", x"6e56af02c912fc75", x"04a360f297efe769", x"b0830f1379da9f74", x"32f32a9c31da6f15", x"fe35befd616a4d57", x"d707e183e83fa3ab");
            when 32616867 => data <= (x"4ed284f05cfc3375", x"2b91200e34c5f36a", x"37db564ebab90b48", x"ff9054d7229e354d", x"6236127e788530c2", x"b276d2db1171011e", x"b8ae71dfce9951c2", x"4621d2d96c0865c0");
            when 17147029 => data <= (x"04498ad2c2822b76", x"a81710fe2273f547", x"883319e21a48119c", x"334ff3c5c65ac635", x"fbca14907fa96458", x"706eb3c1ce99f3d0", x"b2317a2b2e9ae8e4", x"cf8d1f7b812ea712");
            when 8623489 => data <= (x"ffcf3114f290d770", x"1c739d8088b45b51", x"618033810c52287a", x"2014962520ac5f69", x"a0f907886d539f3a", x"b7f05aa67caefb08", x"a17e1b9f4c0d5352", x"d358f37a26b6b817");
            when 31508854 => data <= (x"f4b5ab8b4b172f19", x"ab25774baceeec69", x"d07fbca07924f605", x"09d680936fe36d1b", x"2bfa54e8a0720c57", x"a1fe68001fe88be8", x"739305e872715b8e", x"b483840772f98d97");
            when 23021163 => data <= (x"fa87e61712af4f31", x"df009a1003d75367", x"e75f887e804be2a9", x"531d07365d59639c", x"b3e34cbe24a57cee", x"e1559023f0aa6e2c", x"b9ecbf7e7f2d72fc", x"0c0f3186b3245deb");
            when 25847528 => data <= (x"6038796d42f30f14", x"decf72642e2dcd83", x"6616376f73347acf", x"3a71ff1a40d75e39", x"815386c014b43410", x"43222c2be7a6c316", x"15b0b1e6a414d9eb", x"218547d5d9447e79");
            when 31038163 => data <= (x"c6c7c137e14ddf66", x"e41379abd667ddf8", x"aa57cd87cc8f5f07", x"ff4f12403ed9acc3", x"dc8d56cce024f5ae", x"1302b38ab16a98e7", x"9f2e4055041924d9", x"ca6692799bdc38d2");
            when 6611793 => data <= (x"24c9e615074831b3", x"c9ce679d79cf979f", x"75489716ff481cf1", x"c03aba22d1fe94ef", x"26a7ea1689cabb06", x"771d13af9ae1a968", x"c8cf1c3e4b3445a5", x"709f0eee50f6ae38");
            when 5507217 => data <= (x"e266505bca3ef9bc", x"87f4084a2c1f0318", x"5be1e9ab169914a3", x"a9154a3e1fd1fdf8", x"94e87e4df4b3197d", x"1332548b0bd22cfe", x"cdd8d6fb6409ed2f", x"cdbd440d48cc4e03");
            when 24204345 => data <= (x"bdbdb8dc19aaabfc", x"8bd76d88cbcb10f1", x"74678023413aa4d3", x"19f4815d32e6e721", x"c951034e20a4dc63", x"3c63c428209ea5db", x"424fd7fccaf7c518", x"a1591f61807f1e7f");
            when 12460407 => data <= (x"cbf2f8db0ef97a32", x"c99ac8ad52e583e6", x"3f34b4baafbaf3f4", x"1539f08b62f4a605", x"ad38f598768fc253", x"656729f0df80e937", x"3cb6c47e30a7d37a", x"2c36755d9985602e");
            when 23376313 => data <= (x"b539e3c782ab12a5", x"1cde74f2ec18685f", x"2e390291690c7f65", x"126ff5c67840df25", x"c1f189bbe0e0236d", x"dfd35409c1ae6721", x"283c3e24176e2364", x"85788e7a6b7ada70");
            when 22247730 => data <= (x"e6161288d2c0afb9", x"80ba752f633b4e66", x"868c2a46206930b1", x"f7d4a6cfbba79560", x"adc9cd1a4b08f009", x"367a059685abd7a6", x"f2d975ed6e6b6365", x"1285a7ced5f853b0");
            when 1141597 => data <= (x"8df9c533fefdd2ed", x"0548d4be027d28fe", x"5003341cd04242fb", x"a74bc59505c1ab60", x"be6bcde11675a922", x"ae20709cd5a3a720", x"5f5b1d2d5d681a6d", x"19c2bb5375edd8c0");
            when 3453969 => data <= (x"db9ba3dfb4ab9fde", x"423bc7764bcedac5", x"75601d8c3c345cf7", x"748db5b0be15a936", x"f902c2c5882bd2e3", x"3d899c3e00f5b7b7", x"f4993d97a2c81b22", x"36b7952e89b4d88c");
            when 33233063 => data <= (x"6b73c75c47c77987", x"6ba90f8caa12a856", x"674f0e2a0d31e8c7", x"3ca2414e414fd61c", x"6daee4c6c4a17331", x"c598069a8f3e06e7", x"f4f18b080afa2baa", x"16f8a540ef6202c4");
            when 18715406 => data <= (x"28244f6f5cfb229f", x"aea192649c92476f", x"0621d56c44db47f9", x"1706fc5d4019db88", x"5465788cce30eb27", x"1e9f5295e81ab9be", x"4f9a76f737f0d5f6", x"9e54b938f42d4d5f");
            when 5502213 => data <= (x"c030ccfccd2d20fe", x"2b7acad809c6984c", x"058590837c7640e9", x"1df683260f51850a", x"f51a0b86b0ad6b91", x"eee61d641337b367", x"e52990a254027e48", x"164cc892ff69ca3c");
            when 33705162 => data <= (x"8cd5578f62ef444d", x"65e1e8016581f2cf", x"70f51152909c7767", x"8af1ff3d2dddeacb", x"0b241c2ebf695c17", x"3ef7f6dfba559b2b", x"080509cbd7cd70dd", x"f6a9b4c928ef8aa2");
            when 14918410 => data <= (x"3fccdad6fe7cf6af", x"f59264edc5ea17af", x"6724f57af3235b1e", x"22aba617c396ba19", x"654c3e0cab0cb444", x"bb02d4e5e7815c1f", x"7700ec1a42c52b8c", x"8978ea15c0f71df4");
            when 13299599 => data <= (x"3a9fd4c531f78837", x"1ad5b7d9742b0ec3", x"2fec6138edfe7fc6", x"947c8cf622a7ef95", x"6f357899b15001ad", x"47af1cd715524530", x"1037e543b3e1b618", x"e7dc11b104f5bc06");
            when 11993976 => data <= (x"7e630b323eba3f6a", x"eac97021914135f9", x"78fe1ea7890a8e14", x"9bdd48e8a63d5eda", x"cc3145e88d6f3a49", x"2319362ad2e3ecf8", x"8ae77f0c863a3ac2", x"2f326c7ab7110103");
            when 21610107 => data <= (x"e746174f2e7861de", x"294c3cc791e7f4c2", x"3c8a57e5a80283f7", x"39339e125c5de865", x"28ee43fcc87fe602", x"60d536e7935c2c02", x"d8904aaff3bf5da2", x"648ed2335610c54c");
            when 27120232 => data <= (x"14d3ab4fc8832f74", x"b8523c768e6572fb", x"5311b69b5ead6b11", x"65e3690a00a38a38", x"fbbc5511b85da74d", x"ae6fbfed962101e5", x"a67ce91aef7a7e24", x"88295e215618f1f1");
            when 16089547 => data <= (x"48e670391d8961b1", x"30d153c9ed3c5e43", x"134a96c8a89ce59d", x"3f218d61c743826c", x"e85277fe0783f5ba", x"ad8aa10a0cd647ca", x"b1db67880fd73b27", x"bb29dc2217e6a74d");
            when 907660 => data <= (x"455010bd7dfec2f4", x"5f2d8693bc8482e0", x"c72191f31051829e", x"e1cfc72b889e12a5", x"592b2bf6db420894", x"cfc41315e8349f13", x"6d40796dddd94143", x"c54873450b022f37");
            when 26856774 => data <= (x"31c4c3e5553fd17f", x"b4ed22538943d30f", x"40564e58740627fc", x"623ed3e64bedda5f", x"8b2494dc1145b228", x"1127884e0c39d8d6", x"0f83756dce8d5c07", x"16281004a7d55ec2");
            when 9415558 => data <= (x"9d532e8965e1c18b", x"8fc3d6319de1461c", x"04440e915aa96368", x"c2af2a83e3401544", x"cf8ac5bec3aaa4a8", x"8478ee88f26605ae", x"5ae84c9b754acac9", x"404315a1e4a466db");
            when 417972 => data <= (x"054be958ee1c578e", x"79369fb6df9c81bf", x"e3fb7e9196e68a01", x"12e4467bd1e15e87", x"a73b8b60ca12dfed", x"1a376919f1c6a344", x"332d5e66edd10c29", x"ef78f6e5ad9b76fb");
            when 8292197 => data <= (x"5b3ec042552b8aeb", x"53e181ed751f8dd1", x"469726831f026aa2", x"c8f3e8eeae47e4ba", x"ed60746de826956a", x"08727bf4c4efe461", x"2c56ccf9c1a54765", x"7df01e2824f3835b");
            when 4155043 => data <= (x"84cc2c1255d5dc3a", x"4e84e497546c196b", x"334a132092fbfdb8", x"fdd6c9ff87062022", x"a6cf6ed3b65c7119", x"0ab61e858bc6bea6", x"35cf397552e63dc2", x"75a34b1274926d9e");
            when 14478654 => data <= (x"962bd9d4065f1dbd", x"eae12eaedad059ca", x"9783efb9fbfddddd", x"6651e09d1280188c", x"641d70e9a6b48652", x"320f62590fc40904", x"6f54cd9846f244e9", x"c31c8f011a1f2a38");
            when 20359868 => data <= (x"60e85f8104d784f5", x"6b3bef524a199726", x"9338ba32bc00cfdf", x"867e0226d6ed0306", x"e153684785273439", x"c4c42d221b64cca9", x"e231d57805b09c71", x"7cd609a901575801");
            when 768899 => data <= (x"0549e0e308116153", x"6f9b89554c658ee0", x"e939dd7380174e26", x"eff4a6741bee1ee7", x"4b2285f180bd9296", x"17124fa863a1a831", x"011268305ec37f15", x"824db69cf071a017");
            when 693413 => data <= (x"90a720b0c690376d", x"818b28c8a733ec05", x"ab00a21f4f6974d7", x"c3626e70517702fe", x"311c27a87366078f", x"616b6937495d963a", x"d9962f814b49224e", x"dc84dbd9cc30b170");
            when 15989593 => data <= (x"d1565917308f480a", x"27737ef10cb5f179", x"5eaba8f8629f8ea6", x"ecfb0f8d7b46eadb", x"cfe26040207999d9", x"abe7433f5e737562", x"7fdcf64e0dd13ebf", x"7c58cdc06b356ebc");
            when 8928570 => data <= (x"af354cb37296a3bc", x"ed636e6556ad50c3", x"2c0bc69415d81181", x"e79af22d463f4d32", x"8407521336afd8d7", x"c279c209671c2bfa", x"dbcedbe9e7b432ed", x"51e930165d929f18");
            when 7330282 => data <= (x"8aff053db19dc2e7", x"f0a0b7edf7b2a0f3", x"85f519c71882acea", x"847b2d3b163c85a5", x"6b78ed9626039988", x"d2005c69711e4661", x"adcc1a9dbff6c634", x"67b4127b71fad777");
            when 5783598 => data <= (x"5ab46d4d73dcef99", x"fdb9d6751b6e70a0", x"a0c5e29b1e72176c", x"0ff83ca845697728", x"349c99a07073c10f", x"28eb67c6095d671d", x"357808a51911875e", x"b8c4390f5357fb8b");
            when 29282924 => data <= (x"a76d505457050743", x"b5cd5bdc764bbef0", x"53dc2dca64227093", x"083eb6e28cf71073", x"fb7edcad1a3c059b", x"8b15144db7cd782c", x"7c806ab2047bbc3c", x"1743c25e8d0c23f9");
            when 11330832 => data <= (x"50ea748f440a38af", x"9413d22bd6f45343", x"16b548a1707be5cc", x"d277d607e1be4e37", x"05f640a56dde0fa4", x"63888828c1cbe03d", x"c140454b23a47616", x"84dcea4e71114db0");
            when 3267427 => data <= (x"3ee6877d3bbc4d37", x"642c1ed8fcb508bf", x"d9fccbfed6650e20", x"b3870832045ce98a", x"8c2606f2a206ed03", x"1859cf24419b262b", x"43aa4a1029683105", x"1b9fdf64a4c04cba");
            when 30983962 => data <= (x"e91877dc6eb85a39", x"8d5d3cac43850455", x"3aac8f618a8f5fe6", x"447a5297d0a083ad", x"9a3cb8367832a396", x"56f0c0408d05b7aa", x"f542708cd0207544", x"939f2ee002346b39");
            when 1229128 => data <= (x"0375c9e321961162", x"cefe4e36b81cdd70", x"85ee5f79ad024af5", x"9889bc2a4215d139", x"dc884b4c6c2a3f05", x"7548d82121f7b5da", x"723195e43bd5585d", x"9be3ebb48c59dc36");
            when 32206455 => data <= (x"06e975aafa77f982", x"315b437023bc763e", x"f92da9c5509df4ab", x"33ec561eb66d8f78", x"dd28aa1ca507ff18", x"6475c69bd2d5ba6d", x"a0763790b4500ac1", x"e0554403644ef42f");
            when 1281039 => data <= (x"09a1425e5b16d72e", x"28067f407e0ff3ac", x"f29a28f3ff07d83e", x"d5a9950812f8de80", x"a7c086556b682321", x"8c2916681fe09b8a", x"881198c4654f58bb", x"f90320a21c4036ef");
            when 10312791 => data <= (x"5769796b14d78b88", x"42372e5f73fd0ff3", x"9a0ba9871d391b40", x"1afddff388ef91d7", x"d1caa4489258bd3d", x"d0b0a0e7d7f27a5d", x"d723cfb1b9149683", x"3fca3c032c374077");
            when 11371471 => data <= (x"9f7470470d6cfb97", x"417af7fa4b9be6a1", x"25139e720c60a501", x"2f60562a6dc868fc", x"9d1a12fc7fb6de43", x"ed694fc1d2adcb78", x"385fd586a1652ea0", x"4063ade68c6bd27c");
            when 15115967 => data <= (x"536bc48a7ab7523c", x"1e02e5ddb6da61e9", x"ff67db0033b7f105", x"4c8ec4c96272029a", x"9b966dea2c2c4c2c", x"688fbcf51001830c", x"22fc0013dc6c420f", x"99d0a143f6195837");
            when 4012369 => data <= (x"f85b6dd89e6324a3", x"f3aca8c0eab0e0ca", x"571c10b7a654e05c", x"ab23c44a6ba2d255", x"b865c670aa59b09f", x"a4f30fa93301a551", x"68e6ce1a10df41e2", x"44d3f330be105060");
            when 16793132 => data <= (x"4e8a511cebdf689c", x"1eb0602dbe20a9da", x"e5b8d998ab7d9ffe", x"8b0fec4100cbf781", x"bc129b35ea3c1487", x"1f0f7b7139e16a9f", x"82481bece3d932ea", x"4f5ad640f8602ba7");
            when 29684366 => data <= (x"866bfc1e0a68988a", x"2e1d525cc0facdba", x"8c41dc13cb200560", x"320f6262d7121722", x"d0bd3021ee363f15", x"18032aaa223f1138", x"dad736bd8cab5267", x"315ac9c4cd42a7b3");
            when 12848007 => data <= (x"7834c7882b911568", x"bd216b559cdbbda5", x"fea1bb460b580a48", x"71e02ebfd8a0e171", x"b687011e076c0680", x"3a2fd9a4c55993b6", x"d7e76d3e17b562d6", x"f649bd965ceb1ead");
            when 13180900 => data <= (x"e29d87c8c33e7492", x"227b1dfc8804cc1f", x"136e048aa9c607b8", x"777bba1f5d443ce1", x"36053eb73737770e", x"9a5679d861fd6a83", x"adaa3d0fe03965fb", x"d1b441e5d2fab191");
            when 24709303 => data <= (x"20789b39128f2f59", x"c54d11b1cf48e3c3", x"caae3ac1cbea8978", x"fb63ff860224f738", x"21047556be55c906", x"9df6539a25ea39c0", x"47df443b15196295", x"aa7e03362df24a8c");
            when 4713952 => data <= (x"c01a8b6b3d691811", x"bd7801f31a07e161", x"dd706165392e88f5", x"db0e5cd400ee66a5", x"88153f38e482bd87", x"bec4e949b297b24d", x"94d3d8b0726f6a1d", x"aaa7c2ed1185e722");
            when 19823188 => data <= (x"7072337511b1461a", x"01636d9e88c93915", x"03019464466e6f31", x"4572ac0bb36a62ad", x"c6acf8a241b8b50f", x"9d0faf3bdd5441da", x"907f000548038622", x"c1f97aea12907491");
            when 22479854 => data <= (x"fdebac6239c561bb", x"093534f1751a59a7", x"927a3e2894d143b1", x"42e3f6b5587278eb", x"d8ccf3e51167e1b5", x"177552f82f757d86", x"df1f6b68ca1f5507", x"46b61e8609a22d5c");
            when 13139658 => data <= (x"a5475e1e86bd5b2e", x"3e3fc3ee81eebcce", x"3cad4a0b0c1eb249", x"1262fea7c5761cb8", x"25facb51b3c1cc6f", x"ed6826d34165b2d2", x"01384bcac46e3673", x"efc05683ec006ef7");
            when 31860799 => data <= (x"969b9f1dfa031515", x"3f47f729262b59ab", x"062dbb423557b65d", x"e265b052e5298818", x"422cac53f6c05f68", x"44f71624a13e37c2", x"ac004e64587d5947", x"8074f7a17f6aea52");
            when 27060266 => data <= (x"becae3ee032ed165", x"864857278b748ba0", x"b93b679b9ec141ad", x"6dea12040e49638a", x"b2e28c665ec65015", x"87af4cbb29c74e51", x"67bbe175d2bdde2d", x"4f19e0cf8d187768");
            when 6450167 => data <= (x"4867280d6207556a", x"1f01e4bb7eca7caa", x"320ca56deb8cbc05", x"15dc3e774e205536", x"8ebaf69ef8268575", x"6809691898b9d2d5", x"3ac3520870d6ab9c", x"ff7db66d86e0818f");
            when 15857402 => data <= (x"cc3bdff7130f763a", x"d3dd278506c80900", x"05420eee0da52de8", x"998bd0ff1c1faa04", x"48ed7839534945b2", x"58be107d23165689", x"e162551c58b8e20a", x"97b9127062a19d63");
            when 7003186 => data <= (x"3018d8d0879b8c83", x"ab2da19d0747d25b", x"cabe759623532f45", x"ab3e9788a60cb322", x"14ce2120760754b5", x"fd542426516231d7", x"d64c828addae78e3", x"5bf91123c4775637");
            when 14594294 => data <= (x"770c34195875f35f", x"1c4cc6f87b0dadc7", x"42528ba53b5d099e", x"383c19bcb7f5d89d", x"93add8f58345f815", x"945427e53ab837a6", x"a7897009d03ff379", x"a91821a9fe00a72c");
            when 4512203 => data <= (x"6a6f92aaf887160b", x"1f461a3a382b5043", x"33a62d8e4369f5dc", x"bf038f35f6bdb587", x"9c171b399806ecf8", x"f38701dd53df3440", x"9f2042ef9f86fba7", x"0a50d610ff092b40");
            when 9319488 => data <= (x"220c67ce201a1152", x"4f6a2c6382688e0e", x"d34a87a90fce09fe", x"ca040c3db29ea386", x"e7d65057927a3954", x"13e943bc11462f45", x"45685a97189578b2", x"ae79555dd4c30601");
            when 12481030 => data <= (x"9a729f07facde7e9", x"a3586da3302dcf23", x"9fc16548d217f5e5", x"03a5ee9a63e8e496", x"6de68f0f3f488018", x"027ea7181d0480a9", x"b269fc215f3817a8", x"c04eb2d94a30df8a");
            when 24895783 => data <= (x"1df6b7e77067bcb1", x"6705b9c66f17089f", x"06eab8e8f434f12e", x"3a7a1c2bec94f0d1", x"022c11f095d654c3", x"16648f0c313d70ef", x"ed666eebe9d45300", x"6bfd513d30ee457c");
            when 9259444 => data <= (x"4f2fb6402160d0bd", x"c85d2689f98b6c35", x"0f86c0fd959446bc", x"cc3dc34766765bf1", x"43ff0a5346c3e4a3", x"9c26f8ae0b3e96b4", x"43e6c0fcf2e097ad", x"87403a132b918251");
            when 32516049 => data <= (x"b56449002846d636", x"f1f4cff3651d61b9", x"506d8907053bf46d", x"129cc46731248333", x"9ff6e174ebeae52d", x"5a515c01fd76a000", x"3f898c878f83d7dc", x"b73872abdd179662");
            when 14647060 => data <= (x"73fa9790bf447c82", x"aac21aba04308111", x"ec2737dccade7261", x"27b840274e57af85", x"55787c26061520a5", x"2cdacb1c93353ab9", x"b833b78d2afcf780", x"2be524e55c168caf");
            when 17205276 => data <= (x"483de172978a6379", x"ba09139c5e7bd2ec", x"77092b91d46ec61f", x"ba409d305da81fa1", x"06b43bf05a2ec974", x"b5912be2b7ee5891", x"108a844a30f83c44", x"a5557e964b948ee9");
            when 28136868 => data <= (x"2984c7015aa25abe", x"db351bd5abbe83ac", x"7e77e76262181199", x"07aeedd06485ca1f", x"d02b86c612f638f6", x"c0a77e489ba08783", x"f1bdeedd5556e3af", x"2e597cd309413d5c");
            when 7986122 => data <= (x"934e56cfffbfb142", x"1e3b4df4feb7c1fc", x"0af7013563192b55", x"a3622cc92b8cf7de", x"161e8708c0eec1a2", x"340d8cbb5cff16eb", x"17931c6ba50f4a77", x"68bab28f503afc95");
            when 30461225 => data <= (x"98fb68f138b9db85", x"c0664aed14ac2916", x"0c9d39c7521f7319", x"c57d8db38e5e18df", x"ca2b17dada1de8e8", x"c3f6df49f8abe027", x"27943a4655f06420", x"8ba17ed9bf31a57d");
            when 11815142 => data <= (x"86b644bbe6dc96cb", x"ab285da81effc818", x"7ce77e457d694a25", x"8b20528eb907db55", x"f0732a92d7274e88", x"607dc4a075600ea5", x"48e2366c742c8f2a", x"5f531e40205202e8");
            when 13706062 => data <= (x"fcce48fda9f3780d", x"63208430a7f520b5", x"36e666d1f9638c66", x"2649447a8db83038", x"35b33d9aa671dcd5", x"75970604a5afd700", x"8779b8a0758bacfa", x"8d705d3540722314");
            when 16315941 => data <= (x"1bab39f68306dc01", x"09aac5e0296f73f8", x"299ac5afb4d3a047", x"9820b53371325255", x"8d581e6eafc2c425", x"9197ddaf93775449", x"b6ab160cdef57710", x"cf83e5b4b344e1e7");
            when 24271062 => data <= (x"7f56f77dece4f83b", x"ac65c4ac779cb2cf", x"80f998e4a02b331b", x"04a14183c9bac831", x"203d271cf5271bb8", x"99a4553412059b9d", x"9bb1eaa282eac297", x"5501f961c0beea68");
            when 10027118 => data <= (x"ca7bd6b0bcc9e929", x"de734435221cbabb", x"622bc44a7766b9c1", x"c4eb641ccf1287cb", x"e38e0a9a0ea9e44b", x"4c823ebabc8f38f0", x"41af85866510bba3", x"d581dfdef7b54efd");
            when 26022585 => data <= (x"af785395f4be0515", x"3e67d800edbfb743", x"8a3a933484446860", x"0cc465af994788bd", x"41fef3c410299cf7", x"9c0bef6784371fa1", x"154baf5cdb2bada5", x"bea1e73f88c7d62c");
            when 25448237 => data <= (x"1301c9681613b543", x"2f4617cfd5f49c3a", x"8d64cd204c6e2da1", x"8ac406af463e54b8", x"5457989073149c4f", x"187207c5879bc303", x"4db6b55a05bf407b", x"d1b42153255fb77a");
            when 19329494 => data <= (x"d6e20b082723265c", x"619fdd8877b5d275", x"7ca2fe8ed40051a4", x"54dc3a2935b9cc14", x"870bb3acd7077bfa", x"61d982800a764a23", x"8ceef49787697af9", x"4f7f38d5b24b99b4");
            when 9307622 => data <= (x"017a971704f94faa", x"0c899572496d981d", x"db36ab7c96d84846", x"0e710cc8118a9d01", x"5642d0e08416b38e", x"c8894c5f976d336b", x"693b5dd3e2759155", x"cc0d049c38abf13b");
            when 25730423 => data <= (x"2a108bcc367ec76e", x"cfeea54fdb465fce", x"755d3aefd6fac354", x"ee609fb6f3986d33", x"1dbca38a77b0da4e", x"cfcf5b0b10836018", x"2223800f6999d619", x"8396e8fc583bca0a");
            when 3847531 => data <= (x"7730f0a47b382d0f", x"7cf6d88e59db96aa", x"232667e6a9c08131", x"c84513a5054cc50d", x"d67a0982ec2ce6dc", x"d4e30c58bf6db007", x"3276a9e40537448a", x"6f3355357c58e7c7");
            when 31164648 => data <= (x"013d5c435334295f", x"747f2d1a4a409fe1", x"db4bfa81515a5f58", x"dd98256aa5f9ae7a", x"d0ff93512393a7d2", x"8aa282ef07d1be27", x"d1a17793daaa082b", x"dc50fb17e52fa318");
            when 15422415 => data <= (x"a475dabb6648f546", x"28b90e634809453e", x"8b8405a891128efe", x"e8fd4d9ce01c7461", x"52e72eaf828fd803", x"362a4c0ba2f7ab68", x"bbc9abff6e9b554a", x"181c1cad405d41c1");
            when 5523088 => data <= (x"4a2adf4d0591c1b2", x"184eb36469baf0fd", x"40a63ef8168b4bac", x"ad2b2f39d8efba65", x"22a731f4bcf260bf", x"cee07b2e42f45971", x"9a6e3f66327646ee", x"d00000ebaa4271ef");
            when 12345949 => data <= (x"c9b012b0433addee", x"704c7701fd1e5c09", x"d34640a2b8ee32ba", x"993f560c597e8d11", x"d6a6bf3d35b543a1", x"352f8096dcf21448", x"fa03b7c85c8912d9", x"605cbdbd6b96f652");
            when 25782708 => data <= (x"188c582d7a1e9e47", x"d03a67f1875d6c4f", x"0eda0d8f5eed940d", x"a5f6107395e4ddbb", x"e52c20d89cf557c8", x"f17d2cec69f69974", x"f7c42fedf7a712a8", x"ee9030a48de7ffb0");
            when 15701820 => data <= (x"3643d1d0cf91c632", x"68c7063a3c2d9279", x"dcf226fe47bf93c4", x"2a45bfa486b1e447", x"effefdbb8dbead00", x"8a81f7b9f37836b1", x"4e836d4f4112008b", x"7cee611f92e423a2");
            when 8349780 => data <= (x"077be89b5f161bdf", x"b8f065988f2b995f", x"8085a4590c6c312c", x"5c97dceceb280ef4", x"5ce1aa955de9b6a5", x"cf6bc145246db061", x"797ba570ba0223f3", x"e7ef0b07e413c205");
            when 13060930 => data <= (x"0387667b3099deb3", x"910be8f42c6135f6", x"8f591eb2c68697f5", x"0c2505cbfe6ee9ee", x"7ee19b051d869b14", x"5ae2ae2e82438072", x"bc6d1a1bc5755e4b", x"8750ceb830b29a91");
            when 33794443 => data <= (x"e757ce7d3e102eb6", x"9ab118476b3fd503", x"6966eacbab1e8ce2", x"7b945908e7e616b9", x"4375ff045e080c9f", x"31032c7de63be36b", x"501c48ec1103c683", x"5980decd24cbd97f");
            when 12790325 => data <= (x"1e776bf1fe95e240", x"366fe672a891de6e", x"a0eea3b27933fd03", x"b6af72ae1ee8e039", x"aca5ede2884698fd", x"6b053c21f0165068", x"cc79ceab755362e2", x"5a3574f1f379ef6b");
            when 20848982 => data <= (x"a9b7fd425382616c", x"df53a0502a7f2498", x"4a161c33bc378002", x"edb777ae069c18a3", x"4947b48d952db6a0", x"1ba80ded5595f071", x"c10eb2979b82cd24", x"2892b581a7293f7d");
            when 9122367 => data <= (x"b08842c458a7e876", x"4011fd37faf30343", x"20c993bbf30cfd84", x"ad0119c97a9a0e1f", x"382a08bdbccd295a", x"f154da605a9e537b", x"fdf56c20a00165e4", x"a376f85b06c50b2c");
            when 17261279 => data <= (x"9d4afbb32791eb93", x"39d9b3efb105ff32", x"59e994aaef57da38", x"25c726d317410c4b", x"1eed0f9e233f10b4", x"0735b639c9b3376f", x"467552ebdad46a6e", x"948af0ba7a05d751");
            when 12796651 => data <= (x"c3da978a541d51bf", x"22e92734ca126768", x"e49eabf1c1cbeaa0", x"94ccb20febf78c90", x"6f4c0124d915888a", x"bb61bbf3e59e9738", x"0a2c9e3e9559afba", x"ceef2ad4232076ef");
            when 4007823 => data <= (x"8d84629c9a67babc", x"90ce7a6863783e69", x"0b35a51d2e087aac", x"c26032ca0e2c254c", x"90532f79462232b6", x"8a3ab9791b7c6082", x"ec36c94895473358", x"6a06348576092d87");
            when 20283426 => data <= (x"69bcfef97bacc4c2", x"f361629f82a2e241", x"dec7b186e723f30f", x"a0eda34536731c55", x"4f1fa537d7303385", x"9b87bf4742431050", x"02eb2a919affc6b4", x"b58f70bec5310bd8");
            when 9378138 => data <= (x"3a048c608e241ad7", x"f96ed74bd10c4399", x"0c41b8f9bd7ab7a0", x"0adf85a433a1abbe", x"e4616aa548473eb5", x"aa6c3a248a87301f", x"3e1dc5bfcc26827a", x"15eb96e786db8306");
            when 25447627 => data <= (x"36581d81f9cb4cd4", x"fdfb9bb5845e9b32", x"3ed8414ddb1e6c81", x"6aefaef19b5e2e3f", x"595cb7c02065a7d7", x"e25014b0339f1e30", x"36245a12e70d0c72", x"cd0b9b4e8b78c6c8");
            when 17871306 => data <= (x"f22152c5f380cb94", x"6aa01a5ccef4ed7e", x"b53f3569bad64b8d", x"49e36fb12ce9f89d", x"864beadadb6744c8", x"d4443c708e3a00e9", x"6b6afe9a139818c7", x"bd5b944e3f33803b");
            when 26432673 => data <= (x"19d2f5f5edde801a", x"6e90bae113c9c3cc", x"85e6998394acfa08", x"b6f71631473721a8", x"35e1e25c245ad750", x"b7cc8cf04c2db179", x"1b355d6bd5a189d3", x"b3cef0bb90e284f4");
            when 28046345 => data <= (x"a6dc527360647312", x"aa225b91d04ec674", x"d727fa3af00a5ac1", x"96853c3520ba4412", x"b35711ee987a6172", x"64a1caaf85f1b890", x"45122caeb814dfd7", x"bd2e855d20edf6bc");
            when 28898493 => data <= (x"be3cb88fc02b47d9", x"9cd6091d110552df", x"8353f712dfda55a2", x"812d6749a4a2ab6b", x"8b58021fc70b186d", x"ecec179e34555dd6", x"656af3684a1a57fe", x"b3c098bacec5f197");
            when 2134527 => data <= (x"7c21239e4a5f8019", x"fd839cbc1851fef0", x"055f831962865e2d", x"1052cd3ed686519b", x"3279bbbca0b49222", x"4298ef6a95aec047", x"6276da74f76c46b0", x"e82440a30368204b");
            when 26330156 => data <= (x"0e28c30b87c0e9c1", x"be8dfb87caec7ec8", x"626f935bb1d5a6d3", x"1e961a0148c7a7da", x"af18cf57596b765c", x"182115fe903ec900", x"c704b621efbfd7a7", x"b07c0d3922f990f3");
            when 28317899 => data <= (x"283d880546a304ac", x"ee39d658fdf1fa08", x"60d4ace847e1a22c", x"ce8abef359912fef", x"0f635b58000c3576", x"9dbf7d55bd30d2a6", x"f63b76da078929a1", x"785c131b072eb2f7");
            when 24687962 => data <= (x"8b9bac553f452e37", x"8ac2b7757ee6ae33", x"b49b3b5a4f1b60c2", x"5c44396a0b08bca9", x"f990b6039caaa608", x"d818226b58d92e9d", x"c9a133bf595b3190", x"438dc616c7a6be8b");
            when 16979957 => data <= (x"85071e0da2a038b3", x"faa542e8fbe02dbe", x"72b3a15584a3cf85", x"5f472d902e0f642e", x"6c539ced2a9b3606", x"1d4a1305afe79c4b", x"89e657305b76bdbe", x"442033cbe0507393");
            when 12534538 => data <= (x"5bd31ded50b05ddf", x"3d97e2104b05b077", x"92f54133ff27a830", x"318904fd6f321abf", x"93c4010e76bab2f4", x"e45f529e18721d20", x"e713330d20948879", x"039a740191c1dc83");
            when 27975425 => data <= (x"5d868b9a16563f3d", x"8c17102bf5e3a624", x"63201f70117bb71a", x"3a9b8155b79546c0", x"7327ae17e11d9e13", x"dc0bf148e4495636", x"1e2aaa4104e942f1", x"5e18c544b4ca1f7c");
            when 25122686 => data <= (x"b2893404518e0585", x"f9bff19e560af4a5", x"71ed462bf8c5e2ae", x"3a470f886d5aca29", x"2e9286e08c0c653d", x"810bbfd81ede88ce", x"dbbdb6fc77fc5afd", x"c13be3f291a839e0");
            when 1419130 => data <= (x"767d97386e62b7ba", x"11d5696b05ccc843", x"f7fab3d6ec984cdb", x"0f14e65911afcc16", x"a2ec03c6b937d34e", x"b7c40821af40546f", x"0ccd889f25ec5a83", x"1a68547ab5e0c817");
            when 7008321 => data <= (x"dfadc79d6875c7a3", x"3872ce4a560ae8d4", x"649e1f6536bde6aa", x"4339a43074399e54", x"e788e0d6a56e3272", x"afd9569ec37a443a", x"0b2a132c44d1b62b", x"f360347955eb3711");
            when 28629644 => data <= (x"eaffe8bf2da6cd8e", x"6f0ad2108bbee163", x"f4d2835d155395f1", x"07c3ff213aec0750", x"fdcad1b06f872b1f", x"5f7f6ebc2714480f", x"d59786219d6aece0", x"1b941500c3f8ed9a");
            when 32210807 => data <= (x"2eae0f02deca92a2", x"3b8b62f8b78c425a", x"4b91c9ba52d21573", x"900fe85d9b72ca29", x"8ea158534e0ec0f1", x"e31ac100fd0d5c8a", x"d0dac5e54793b281", x"65e16f245b3ca2df");
            when 15172569 => data <= (x"e167822b40728a37", x"b8e6bf9846f81d37", x"837638bc20cca5df", x"dd07322ee6266943", x"43c61182fb532b70", x"4b4c5cc0b72d9710", x"bb5a10931feeb37d", x"0e6ceaf2ef0020b3");
            when 19970153 => data <= (x"c64133c13eb3b1b2", x"8717dd6de2d7e85f", x"2808713793399fb8", x"9607da56fdb5db75", x"9742637618d8328e", x"1bd735c7eb8b8320", x"dd306800fc433499", x"7be7b9e2d0faf542");
            when 7819389 => data <= (x"ed63f89afd0203f3", x"72899d3b0f634727", x"06ca1d879334441c", x"ecfeb298de6126b6", x"e05b1e3e01b495ca", x"a0bf4e229540cf41", x"4b7022d9609ed271", x"d9f225e685e488eb");
            when 20783808 => data <= (x"1de9411eeb3469d7", x"ca541d3c8e0a0384", x"c50bd70cf944de19", x"8ea1b7bc62bcd93b", x"9cb7aeff5add7aaa", x"2ae5afab8fdf4c1c", x"ce622e7da4135787", x"f8bed3f93cc92610");
            when 859896 => data <= (x"e6cb7552fd008ca5", x"8926d5c121f8dacc", x"03b3f09b2c846675", x"4f8f825aeba3ab79", x"77b715ab003303d0", x"b49d6949a6aef75c", x"d89049d7bcb5901d", x"ef77ea5280d2b00f");
            when 33330927 => data <= (x"607575478f6f379a", x"9c2ed2697b6f88ca", x"ce3ec16d161fee1e", x"7442c1d8ed35cbf0", x"8611514272b5840d", x"2ae00adeee1f306c", x"5a63ada636ea7e32", x"1097cddcfe917778");
            when 11015924 => data <= (x"b6e121bdda01b6f8", x"3bfe4bca1503ae32", x"c21e2bddb45879e9", x"4e16b70eb0a746b5", x"6069e6ac4fc036ff", x"ceebd5f89cd6be97", x"b3920935439447f2", x"d94435f1e9c940cc");
            when 16594274 => data <= (x"77fc4f2d4292af62", x"38a590b28b30f773", x"9c84d1c90efbc9dc", x"85e96138f3bdc6aa", x"338b06e6d7d0a28e", x"aa02037688e560bb", x"45e223d9080fee70", x"57ec82a6e30f8ad5");
            when 33246450 => data <= (x"bfb53729f4eed0be", x"18cdfd29c0762b51", x"43770e2ae72b147f", x"338836c33c06cd3a", x"038442bd8811f5af", x"8e032d82d468036d", x"1f5b54aa1b06e83f", x"0c5ec15013195780");
            when 15663896 => data <= (x"d226c5894d3e274a", x"9c2c13e9a879e436", x"141cf30efb2a6e15", x"2e608acb24de4fa9", x"7fcc20ed442985af", x"653c83d24b76b27f", x"29ba281225a5056a", x"92f57250b2941d38");
            when 22955915 => data <= (x"ccbaacc3bcc4a507", x"2723a45d48412285", x"a15195876128bea6", x"94c015a1b3555c3b", x"205b2bcb4d74acc3", x"fe5f417e463f285e", x"85631b09cce9c976", x"0e9d085e9421e1d2");
            when 10566268 => data <= (x"e16e8cd5f2db0626", x"36b1f9ba84cb05b8", x"f36771772ae54709", x"405b2fa20f51f815", x"01ebd4108cf31671", x"2eb965029867113e", x"754241beb1bc9545", x"9d27ed5e9bbe8cc4");
            when 29301460 => data <= (x"9f884e88b59cb3ac", x"f4fdabba4b68fd9a", x"0fd59f669b8dc04c", x"139ab56f05aed677", x"63d7eca84986b2ac", x"fe22e635c3f1dfc3", x"6244dd97004778c3", x"4c2aa26d323b2dbf");
            when 11342198 => data <= (x"c1ae3fff0407ecc8", x"faf937a321f39403", x"537376ce0d673044", x"d32c6dbd7840c237", x"386e89cd6fd3e7ab", x"633f256475bc6dc8", x"f00cc0ece5e5cf2f", x"6e65b3668dbc04e9");
            when 19921914 => data <= (x"30d0c5c3d3e54658", x"265e399fe2a9c9c6", x"836106a83953415f", x"717da5449d66b519", x"e4c384a75cb64b27", x"026d6928b44b1bb5", x"c478d9352532aaf3", x"0e432cfb9220ab85");
            when 14595847 => data <= (x"4d324ee73a7ec96b", x"07b15b7b44c556fa", x"2dc2c8bd7707b320", x"25f46f37abcca063", x"2238dac13da15a0e", x"53361430d052584d", x"5065cb4b0f70b34c", x"9f8dabf6df5c4882");
            when 32036498 => data <= (x"622a6d57d3191296", x"518fc731d2b952c1", x"9128edf3a7a66689", x"c37a906e5617288b", x"376f8801fe598981", x"e2f03507460e23a4", x"ca24b3cc78cf04d7", x"a3e85d2f1d71b543");
            when 2392340 => data <= (x"5ee9d0ca04eb126f", x"5357dae076d60c11", x"e8c17cf62045630b", x"6de1348c88427e48", x"fb1192b981f287d2", x"dd33b0c719ab0a0f", x"f1f5b25c9db2b3f3", x"80703cc0376a566b");
            when 7735068 => data <= (x"f47d1681572efbce", x"6612a4d7092bb3d9", x"a841d2e1f84cd3c9", x"4364f7acf439a8df", x"4975f8664a83edff", x"39802d2d474f25cb", x"eb1c6e84cc81e1a9", x"cc7e8241e2bb54af");
            when 25280483 => data <= (x"cbfe5fcd45daa7be", x"a782489692361e21", x"48c95a4425c17f51", x"3765d2d233d96c37", x"f494b6d79f7b1e70", x"4d4d2d11b20d3ff1", x"d42378759aee987c", x"24b0a5d1cb85a708");
            when 26755808 => data <= (x"48ca07bd75d24604", x"9f1eb21393803419", x"dca0f0a0c7ef0cc5", x"8d5c7f7071b17f88", x"a409d1b333f382a3", x"3773f4ae161554de", x"0ee094d46f20f610", x"103137687265e574");
            when 17418376 => data <= (x"6b455b1e37eb24cd", x"22e1e946ae8e2739", x"37b8884c67c8a599", x"23a67d544513ec1a", x"8d17e89e25a8f4a6", x"267677237d3fe21f", x"5f1b51ae3a484d1b", x"d9a346a4d7db724a");
            when 27868803 => data <= (x"e330e462e63fc536", x"5ed664eb3def7f70", x"e915958f31eeb86b", x"7c4b89583b8a87f7", x"1b42328dd5c9ee7a", x"de3c889a6354ca03", x"a959aa1480ca0cc0", x"3dd7c93ba68a5104");
            when 18065799 => data <= (x"966f04e4dadc9233", x"1ef0205b029ff6af", x"483406a7c135a745", x"967bf299bd962fce", x"b8a59bb8a48be3c5", x"1eb9600e1b49d213", x"d4f6cf42ea478f60", x"a41cfd93ee413ec7");
            when 30096807 => data <= (x"00ff9cb684370166", x"9c596ef60522f264", x"a8a9fa73968a2864", x"17bdbe0c6ec019c1", x"51007aaa1eec194a", x"6907602140383aa4", x"17cecb2f6112710e", x"8b1058764f2bffab");
            when 16638001 => data <= (x"20bdb8838a35ec99", x"55c297dd408e0092", x"095e41f0a50ae7d5", x"37c1651103eba402", x"c46c72c9dfa30c34", x"99a6112794cfb28f", x"66329fca484cd6a1", x"ac9fc88b587426c1");
            when 26916412 => data <= (x"935a6725fb844d8d", x"fa5c654d126e9e62", x"b5de9435a0ef4096", x"7d678fe37aabe642", x"cd12fd0a5fa25407", x"4cd1d5aa53572ef9", x"0d5c30eded1fc723", x"2eb05a1911c67c29");
            when 10776930 => data <= (x"55621e8dec2394d3", x"d3ca731a2a9d05af", x"80bc6d28e7af71ba", x"73539ae8b58f5baf", x"588d148e79ff6cb7", x"b306ebf1c74f7fdd", x"cc06bdaafadd39e2", x"b88060270b2cfdca");
            when 10290559 => data <= (x"b09b03d8c4941b1a", x"022cd91b2ba0633e", x"52da7f4f03403e49", x"141c68908ea9c9d5", x"a3133d7dc0085804", x"c1ea185e23b99558", x"c2989ef2a4f6cba4", x"098d290f57b82413");
            when 31849053 => data <= (x"d39151581ae7f5e4", x"2a14b1e3ba9e78a4", x"d6c00710f957efd2", x"378f9b79c48b7b19", x"658233c7cc1984ec", x"e47f42720828a5a7", x"7b95f07df28f0480", x"adb1fd7c51989461");
            when 16264390 => data <= (x"597711049525265b", x"0944b279e6bdbafa", x"f895845e3aadc8cc", x"f7ff1b8016f6149c", x"0f22116495f2fc34", x"4170ea43c7e7119a", x"9621dd3914fd2fcb", x"c35757f2f6fd5295");
            when 22503101 => data <= (x"dd39d14c48ac50a8", x"8838a0ad98d90c27", x"f5bb57473ce2f8a6", x"676736b5b6969279", x"795bf50c165de539", x"9c0a91ce7ddecdb1", x"f79c21bafc5a2cce", x"570c8a59324a6418");
            when 32510270 => data <= (x"c8618422094e748d", x"73d71f9565469b18", x"b7c492b8a2792be7", x"fa6f3110959a1b76", x"bb6944b8aba3171b", x"24368cdab511fbed", x"770a69e38192f70c", x"546b34374143f1e2");
            when 31762662 => data <= (x"5be1bda0fd23548d", x"6973b6f394279006", x"2e62eda2120d40b0", x"9dffcc0ca6708da6", x"3994e129c90213a0", x"67afc37bd4d0cea9", x"6a2fefce42d52dc3", x"22495f243ea26af7");
            when 21909962 => data <= (x"5be1ba1b85aa3ac5", x"ba536605a2ee652c", x"8c6cc15247d053d6", x"c74f49861956ea63", x"fa8b1d2f50e2cc6d", x"c267aa7b066f760d", x"8143c5a5c0f2fd70", x"c2c8c5f302be9a23");
            when 466944 => data <= (x"8802411b898af2f0", x"7538e6a8380665ae", x"d506010d8ca66915", x"13af575262d58e35", x"cc46539d10908381", x"65056769d230b0a8", x"080d94e3cf8b9c22", x"51a815f7621a9238");
            when 9232832 => data <= (x"79070fe57a409451", x"0d46411c64f50223", x"eff24691292be2c9", x"87c5b3a4fb5b4212", x"92da65f72fccd274", x"15365006b4fbb717", x"91039872f2e83675", x"96feaa27584ef81a");
            when 753103 => data <= (x"a45c53bdd3209502", x"6735e2ac5d35e904", x"c673704fcd5a77d3", x"b338a1512add96a1", x"317cee044e3b8de5", x"f1ff25ddf34fa19a", x"9c962e64408285dc", x"b8c6f0ee09d43103");
            when 13815072 => data <= (x"3ac18fc9072c0f99", x"4b2df5e9e08f2b52", x"58162003eca75fe4", x"cfe105a8ef17436f", x"968190b15af615a1", x"42ca113581d16145", x"cab0689970bd4939", x"07ac5683a6e3fdd7");
            when 5114241 => data <= (x"545960db3ffe5640", x"f8e754799a7a4db2", x"1f5532b52741deaa", x"d06fa38a9232ae3e", x"b3739d759fce1f54", x"d6c96a24ea807707", x"6c29f8ee221324d4", x"43bbc28d2c8aa83d");
            when 25881246 => data <= (x"3f6c0e86d73d0da9", x"b0432c6e76e6ec14", x"b249e56ab1c9a9ca", x"df87c3f4f8ce470c", x"05ceb6ca5300f23f", x"b0f3bb23217dfe49", x"46a8b4153cb9f785", x"0779eea53298dd17");
            when 20917410 => data <= (x"b97f61f81850f919", x"25c90977e080e001", x"194e67397e39a510", x"9da3234cff402573", x"5aad2c6027540866", x"c5e5a3267d8a3a30", x"06422feb97e3f3d2", x"b88681904049b690");
            when 9999784 => data <= (x"174daa853871354a", x"17c01678be8665f4", x"2c8612015a50e829", x"5b3bced8502632a8", x"f1c279783b7808a0", x"ee2384c0dac5635c", x"cf3bc7154dbf0ab9", x"b271c47017c42ef9");
            when 21225630 => data <= (x"38865c9c3d953776", x"7ff16fa88f96af7f", x"ed1d0369f26fb4d0", x"562fac457252ebb1", x"11a48f587758d2db", x"cc7c2aec67f65ad8", x"c49f4fbcc68b0f0b", x"9cfa7796b615dcaa");
            when 24915522 => data <= (x"8dfb5a4b4d83872d", x"c223034025c9cf0c", x"b2e359f5bc63c45f", x"2decb947684ade9b", x"cf7f115b9a373597", x"d41d590d62a28e0a", x"2fce7983c1d3f798", x"1b385740d84beb0f");
            when 28195281 => data <= (x"c2c29445d8bfc195", x"333d1fce7fa6d887", x"4fb231870f424b9f", x"8768048227183e0a", x"bc7632908af9441c", x"13fec3dff7f73b9b", x"8730d7f0da1bbdbd", x"730651fca1abed67");
            when 4823130 => data <= (x"aa03a9cc54f2ade1", x"19f7a02b37b996db", x"479ea0c124f29859", x"99eed169c077898a", x"913b20db8da9c8dc", x"93ed5f66c9e19436", x"fe5dd2d5733e0f10", x"eb880499564201da");
            when 16057628 => data <= (x"7ef6187903a7da4f", x"7f4e1b5712519c50", x"95cde9225b1cd1b2", x"c5128e6527ec53f7", x"9b5c879c0a136cc1", x"db7c14033935a512", x"40c674f5a979d749", x"d4c6ced83d0099ea");
            when 15903631 => data <= (x"47ce6645a4656309", x"fcfd9440890f6a95", x"2725b2550ed9876f", x"d9bebc80b6be31d3", x"9aa8cf645dd83533", x"1a0d8d28561aea8a", x"57adc2035074906a", x"61fc5291c5a4e274");
            when 22734027 => data <= (x"b1bcd2b168fab215", x"5c96c541312f1d37", x"9c66b565f1d8cc8d", x"9dc6c5177caa59ce", x"c2aee2ebf53f2ade", x"716bdc9488280a7b", x"83ba8868dee05a8f", x"5900e857e5afad88");
            when 11313698 => data <= (x"c9a1956de0afa58b", x"a0b57d49e0fd2131", x"003b35c46b2c1b4b", x"8939bf5e5747aa75", x"38e0e0b2f8209942", x"3afd400e66d25b75", x"98a588fa6791fc7a", x"502cd1d77c28dd30");
            when 675456 => data <= (x"8029d7155680723d", x"a0363d4a8b363ab2", x"73df7e2a891d0c7d", x"3bbfd3148749ff2a", x"4122ebb41e26b80b", x"285c44185357afa1", x"088abb4464057282", x"8dbc637aa858213e");
            when 10987096 => data <= (x"47ee584f1e0d4a6c", x"8d382987ccc76c7b", x"f00a1db5719d55c3", x"9e1834ea8f7f574f", x"c1289707ebc45ae7", x"e9e1984fb81e13eb", x"9246213957dbac26", x"34b0001eb4a43bc8");
            when 26391626 => data <= (x"80f823965865f4de", x"35b0f1f665f6d8ae", x"76bedd1fd419a3fb", x"f6693ce5de367465", x"137da7e23aa2cebe", x"1cbc819507d7e751", x"8da713a0dfe028a2", x"296758603aad115a");
            when 5491987 => data <= (x"9c1a4dcdcc5fd98a", x"4a4c58801ae9c7d6", x"20994acf97c18050", x"c9b54be284600afe", x"bcc33c6d95a12c66", x"96192d99114c554b", x"854fbf5cf09eb958", x"5c43dc7424cfd87d");
            when 28309242 => data <= (x"c93298ba1649b01c", x"3aef826232def172", x"699b45d782e66f9a", x"a816d71eb392df3f", x"af4004691d9f00c9", x"7b48652aaceaed2a", x"017c41bea1fcf95d", x"1029d6de8dc29422");
            when 19558391 => data <= (x"32bc9437be92f841", x"4e0dfdc5c3e00a04", x"1d26cc0ee0d73c5a", x"7d02970a28e9cb9b", x"c13684481d9df07e", x"94cdb5da2cc12ad5", x"5e73fa7614dd73a7", x"b37c22413b1f3a18");
            when 18514517 => data <= (x"864d3a8082a0edbc", x"e48a2a301a4dcfea", x"07b2d60963b43c75", x"1a43580594facd0b", x"11ad8b262c01e001", x"dbb9fc8d97aff553", x"0be2396f1eff57c1", x"192c3ade387fa6af");
            when 13391120 => data <= (x"39f3ca57b81a5c14", x"552125161158d457", x"6e4a701074b8b3b9", x"aa93f8d4ad9c2ae3", x"acdf5ec1d75b38b8", x"3b486ef6da12df9d", x"9fd45906742720f7", x"516233dd76c6d57c");
            when 14073389 => data <= (x"752830d5b4a68427", x"d56f90879e1e513a", x"71e1d69db18ac567", x"6567bf2e6a830ad7", x"0216a0547e03774e", x"09ed7fd09a523393", x"5819b594750d97c7", x"bfafb9ca43b0022c");
            when 15244178 => data <= (x"9293929cacd5b184", x"69646e8263d22503", x"6b52748850d64c80", x"e47e87aec614d674", x"54c5c12caddaf91b", x"1e0bda9ce13edd19", x"a31c94e85cdfae76", x"b66c9aca6de5655c");
            when 27774891 => data <= (x"1a83d2b4992b7bc1", x"f62c3c5dac6d160d", x"91efc4255fdb0bc3", x"3d7b1047e735bfc6", x"a05a14413a037dcf", x"006fc4c3ca7b755f", x"30ef14da76091572", x"cea925e41638ffe2");
            when 29583768 => data <= (x"250784886bacc83a", x"e5a3c2e372f1ae27", x"eb9f7494b85bda19", x"404d514ecc8918a2", x"65ff14f024f15e1b", x"2b33f53796b0a0bd", x"8bd773d17670ad5e", x"e7443fb29f91bbde");
            when 8123774 => data <= (x"dca386e876a44a76", x"4575d187cfd38d4a", x"56a04d4a8c3ea718", x"1cc7ad78adeee349", x"f7ee83f0661982f7", x"d5c85b59316368da", x"7153e9855bdd0183", x"e220e03d056fc1a0");
            when 24660208 => data <= (x"e5f6a03f9f8e0bfa", x"0932bd6f23890d63", x"a18a55afaf4a54ee", x"17999e8b35b28188", x"02fc34f3b70461c3", x"06db24569b318c2d", x"7daf8d34e7d31c6e", x"d1e7a3b4e944183d");
            when 29065054 => data <= (x"1935eacbc6865b38", x"dd91c325dc2c1609", x"44747ed3c63cd5a1", x"442e19b6f3a4b419", x"75d639695c7bb420", x"c11ec1d95911eb1d", x"b5946ac1c5cbb612", x"4b29232a7f0e36c6");
            when 25371682 => data <= (x"afe9df331c598fa8", x"316cb47865ad12a9", x"40279af5ade2f902", x"42d750a34faef957", x"5232d2d5c4a68bd9", x"2f2bff11d1586ca0", x"9c59ad34ec15fd07", x"7af45691807b7196");
            when 31833349 => data <= (x"8089928a9b5b8075", x"95924ba57fa4f987", x"f99d4e2fd0c84e24", x"e338fabc052684c3", x"f01a465e5bfdd480", x"007b77a6ead0e8f3", x"1be7a08c53f19790", x"db5db71b5bd2a838");
            when 16525202 => data <= (x"1df54a0c256ef0d9", x"32fb0cfbe0ac5301", x"0b4289deb18b315b", x"fee78c4a06791970", x"e72509941b99895e", x"e2fefd7dabde83e2", x"3d804ffb7dbbfe64", x"51393568960d3a24");
            when 15640120 => data <= (x"f9fcf7392e0ebf90", x"6fcf84ef3a7202a3", x"8ed33a62083d0c53", x"e1c41bffd3fee32f", x"f3b9b316152dcf1a", x"30ca94dc281ca80c", x"2a1380008feb45de", x"d3a2aaafecedb3be");
            when 21249482 => data <= (x"d12382e6f41d03ff", x"fe0b9329073e8855", x"6f14c7633b7475da", x"c33b0facd11cf3a7", x"4755478269324f8a", x"e23b20b45261af37", x"262f65633084fb0f", x"e8c1e20dcd4eaaa5");
            when 20091013 => data <= (x"a1c19a77529b41e1", x"f48b0d5996088a2a", x"dd5aaf33507ff36f", x"b5a2eefe4d4929fb", x"4692c556b16b0a33", x"f04c641ab78b4977", x"c35b6710681f07b5", x"ea95c50965ba1362");
            when 4358633 => data <= (x"f4a9c20b7adc40d2", x"d8ddfbdbb033fe4e", x"48ce5b47bece9ad1", x"bc174f4723e4c7bc", x"396e5eba15bf0fa0", x"2272a9147e6ef620", x"d71c56207340cd26", x"831706af88a79706");
            when 31514501 => data <= (x"9ef335796cc24905", x"805b0768de38cf6e", x"f9e7c366d5c3805b", x"b1ff18258b67bb3e", x"fdeec40169cfd006", x"4632e504e7d5588e", x"b8b7fddad3e198c7", x"1ecc373d0fe30a5e");
            when 17651790 => data <= (x"9e5773034965c949", x"e8cb24e674155698", x"27ef1142282ccaa2", x"7239a70f48a40d06", x"50a07c0de097b2d9", x"64f32c3a8954dd59", x"883418ba10af2852", x"32d9e24a13407a2a");
            when 5726544 => data <= (x"d0a45a0b647d50d9", x"77526ba04edd1d89", x"162565d7ff243aa6", x"cb7241422b850616", x"38379ac9706af99f", x"9ba9d2fbae4a5b3e", x"73a34cd44ac62bd6", x"0f2392ee6ec44102");
            when 5950851 => data <= (x"b44a4ec08a091ab5", x"9b9489dc320a0934", x"88291ecf4b41d874", x"9035ee5cad6c75bd", x"faffde05232a5412", x"359836eda83e4686", x"40d51c6e56c65b6c", x"a3ade43ac49301a0");
            when 16265347 => data <= (x"6737be591fee24f9", x"e18cfce17a8ef984", x"2922f1b0d735e8f8", x"572bdee17ca7361f", x"1f138eb70229376a", x"a4681feb97db0b06", x"338192f678eac0fb", x"1bb97385936b79ac");
            when 25618007 => data <= (x"09135b0036522c5d", x"ac9ea594fdabac83", x"0424243575085001", x"28782dbd1c76370a", x"7699c9411e675040", x"feca031287601b18", x"733606a9b09c7ecf", x"a7b34985298d0fcb");
            when 849239 => data <= (x"258918318df96a6b", x"0df3efc17a33b1e7", x"043b0f17bd276513", x"7c0e9703ca0cfc46", x"3372011fe4f9b72b", x"9fc8363c0a8c7018", x"f1d2ead204632064", x"69427564b3448326");
            when 2881794 => data <= (x"0e7b19dd0df4a34e", x"956155bb304be90e", x"9e92188caa1d52f2", x"0830543b6db001be", x"9cdbfa830b43b60a", x"442673d8dbbc5422", x"fed6af2b9c016649", x"7e2d365dba1b665e");
            when 25015644 => data <= (x"c0656e093dd304df", x"d7b02a1bcd383947", x"966d1a2cab039898", x"c2e971779fb1bd4c", x"a5e304c7b284cc52", x"27e916502fa95f5f", x"34b50ffdaa610b9f", x"71c39aef316d09f7");
            when 29635562 => data <= (x"c7b397dea458c005", x"6e0a672f61022285", x"9dc9bbc11a34dcf4", x"d0a8ba21532346c0", x"d01a7e878fbb96d9", x"b7a5425a8da9fcd8", x"cbfd7016c68d15ab", x"471d3d94bd220fc6");
            when 10993841 => data <= (x"56ed55db0edaa0be", x"365c7acdfe7aae36", x"84bb8087286919ab", x"c4095388d74f943e", x"2c5a9e34249ab7cd", x"58134c0b6cae9a6e", x"fce0e81af8323b78", x"3a196254ce717a99");
            when 7637749 => data <= (x"408f4009cbb325a8", x"279bc7853537fe94", x"b9847d31aa4be474", x"e739216564751af0", x"a10b25a5f5ba7369", x"61b3db79028623ff", x"811a00e8382586d0", x"0ee3b47503b7d7ae");
            when 26817421 => data <= (x"77399c6004668e31", x"0df055cd14549f16", x"97bd67bacd7180f3", x"16035b815ebea78b", x"a61576e3270a11cd", x"5578d1a6a679175e", x"aeb1698e1a5e7e09", x"c113e5190b4601d0");
            when 1760211 => data <= (x"2b362a57fe5b2551", x"fd077f3686f193b6", x"edf20012cb62b3be", x"cfdec6c04d0eb940", x"1b99dcf0dae6e77c", x"af1150d0f62c9416", x"54ffe6be10e9554d", x"0b86950353975fc5");
            when 24325368 => data <= (x"661983994f76878f", x"ac80bd339b8714df", x"666d53a3404396a8", x"0eb3550a3234527f", x"63afa0724dc5440e", x"2e4bc78e07eb84c0", x"0546f9c87f0d453b", x"ad4535b652b7b021");
            when 23184667 => data <= (x"b44e1fd3b828720d", x"7825b180b7890497", x"f0fe955a02af4c60", x"82134d295f134b45", x"0ada3660daef2500", x"2b1e853e09770b7b", x"b28d8d8f71163c86", x"cb542cb15b9bf7ed");
            when 21884433 => data <= (x"b5f5d1487f221f0d", x"868103f9736fc31a", x"fe434043e0ef61a9", x"3132da84f55f8779", x"c56dbbd7c3d8dd58", x"7b5e5cb08b0d8e62", x"74a8d3d401d76f4e", x"e84a6c1ea3d9f4c4");
            when 11170200 => data <= (x"b8c0b69224c163b2", x"ac00851ff9db24cc", x"8cdec35559106ca6", x"64b6e66bdcdfc6a9", x"0d7bd3b60f08f7be", x"ac2da78852298fd1", x"985ef4cbc370598a", x"68b8bd0818a4e4b9");
            when 969921 => data <= (x"0c4d6a527e856a1d", x"50fbd2bb7e80713d", x"86a22ecd27d41fce", x"6cc982ce9f3dc820", x"52d2c3368d4d2449", x"baf9919f3047f0eb", x"0fd2913cd68de8f9", x"32649aca209c56df");
            when 13670832 => data <= (x"6d38960586cf8275", x"15f2a5d0d1b34a60", x"c7a7910169593ac1", x"1ee0540fe3c9fc8d", x"e5b7e747a45d35c7", x"ede963ec5dfbdc06", x"6f7533c39d2ff56e", x"7dcfb57e045b9e41");
            when 25134696 => data <= (x"2eff9e0d63b25c9a", x"1bf45d42f09aa2ce", x"b2c11ce25d032875", x"e617ab77caf7d9b7", x"3801b42e848148a5", x"12317d94df1f2340", x"299c39a3d4d64f9b", x"e55bff6731574227");
            when 1194633 => data <= (x"ff33cdeb58e205a4", x"05a3253514ac0f22", x"6ed818a6cc1df48f", x"628540e1352509a4", x"4403da182fd99146", x"3679a9d0743d8bdd", x"0974baf7c4f8b5cd", x"a13ab4b27289aeaf");
            when 23271998 => data <= (x"6432f4097e28fb54", x"d13f626569ff81e0", x"9d6d89cd7be702e0", x"9cf9159a05e7c260", x"f24a42f4141fc101", x"f07a4ca24f8cfe70", x"5f18e32135603573", x"425be90e98714137");
            when 8811083 => data <= (x"4368f207b4d09bba", x"988ec77722fdb1b6", x"06f9b88c4559756c", x"4f84f41d22125e5c", x"038da4db5c174bdf", x"274dd3f91c91b1d8", x"856df2f0b6489329", x"bd00d2444f41d095");
            when 25647818 => data <= (x"4a27eb5c3759aae2", x"37e590cd46803b01", x"b631ca5a5dff6cb5", x"7ab34eb5bfb33f4e", x"9200329eb3622660", x"2f50d29a12867df1", x"255ced3f3e17dacc", x"3720a98158ba005f");
            when 6023449 => data <= (x"1bce479b0f06e385", x"e3dbe1a05b4f0651", x"2ae433020ea05644", x"9c03ccac5af31583", x"491ef3449a569d7f", x"b14ee6cf80fd53d7", x"a59c7cb771cc8da2", x"e1bc635b9766ef71");
            when 7789863 => data <= (x"5ab075fc386eca44", x"d7675a280d5a30fc", x"b418cb0577dc82c8", x"98e050eed8dacddc", x"f235c64628729838", x"484cdb30c7ae4a59", x"9726034f2d20dacf", x"b6ea74af08319f16");
            when 18407727 => data <= (x"c6607785674cc7bf", x"461234d2c2b13dc7", x"95be8fc46507a6cb", x"886346e8b387bfc8", x"a3464e28346ac1ab", x"3c4764455459d204", x"ac2f729f9b4443e0", x"5418f1960e8473bf");
            when 33596042 => data <= (x"cd05f9c4c1974e40", x"ac5dfab0662c3c51", x"88299a6043097dd2", x"45308ab55d93de41", x"d20cc1a04e87a82e", x"171177980f803635", x"4143c3a700463f12", x"07b087be90471310");
            when 5581388 => data <= (x"004e22e687480c34", x"68606e349b1b0a84", x"0f9d701846d227db", x"ffd6917c47740260", x"fe36647721f69ca0", x"786b80a58de578c9", x"a4f57e01fcc4b0b1", x"3fbe4e728b6a1b20");
            when 9313519 => data <= (x"d51fdb5122a75881", x"330d693a29229eec", x"ae9063a1b70f677c", x"c0a4067db3d74244", x"c1544a24e921f839", x"6d39d62b99e0529e", x"366f4f5f49ac16c7", x"cadd23f875e93426");
            when 27792923 => data <= (x"d797e785132e2998", x"277bd8ad517afaa3", x"85bfc98ecb4e665b", x"9a5993a842920c20", x"dabfd192d6b7e64a", x"61a65ede9671c1d0", x"acaa71aaa8e34fe0", x"bf7d09662fe41632");
            when 27115321 => data <= (x"ad28958c7aa705a9", x"eeb96d45325bb40b", x"dcc81c8e5f59a591", x"a7a262f610258b98", x"0e0e52a2cf6654b3", x"fa322598ac73ec56", x"8d9c5735ea63c39f", x"c9675b82a172c60f");
            when 24975596 => data <= (x"b1eeeb8b94cb0bf7", x"24c42d3f6b58dadc", x"78d0708365402430", x"0b80ab498659dd72", x"513be51b9183e594", x"067e9833a739dba8", x"cd4a45bf6134e0a3", x"4cb7e2a92d583af0");
            when 923520 => data <= (x"18c8a56172ea9ea3", x"777adcff27ecc365", x"600c9eca2438b036", x"293dde99dd2026a0", x"47dcd0b532b1ebbc", x"cf47263675544920", x"24eb82645a67b22b", x"3cd59e49ec791943");
            when 16277302 => data <= (x"114eb39c0ade93e7", x"1e860f5dc99f4238", x"f615ed3275ece820", x"b90a268bc33f6b51", x"c19328eec5a18048", x"c5bce5c5b6fa2080", x"04d2f9f36facca63", x"4a318548faf8a4eb");
            when 33255108 => data <= (x"1ea92d88f6dfd34f", x"c2ecf3aa664b4241", x"42105af4e432be09", x"59809e265e192c5b", x"27a6ac9bda308bfb", x"25a6559994f77c76", x"3f01c79033b75d30", x"c8634bb5ebfac495");
            when 12002399 => data <= (x"69ddb0535b3a7401", x"e05e5c31b087e812", x"79dab73d37c63413", x"45bd0908b026215e", x"3f8c53427d45b6e3", x"da9f472e4004e045", x"62dc8335ae5601b5", x"48d7ef4fd5dcc7d9");
            when 14565621 => data <= (x"0e765c250b1546dd", x"539d5eb5dc4a20f5", x"5872d912af53b3f9", x"d4e8bf2e6424f244", x"e1d63165392be14d", x"6568936373e12ed4", x"6b610e9a2395966b", x"d8ec541e54d9d9ad");
            when 8340108 => data <= (x"4db43d850691c5ed", x"30300356258a2e36", x"82e873b59c05e349", x"e3a7e6b25ed51f2f", x"c50683120ef85971", x"79123498711c0af7", x"c967e3f7c60960c0", x"126684c8a4da6cd4");
            when 5111993 => data <= (x"bc4e7b6153f3020f", x"0a76ec0e5905a6ec", x"6603701e82064ce9", x"afae7e9f54ea1555", x"e7e8535024891936", x"4bb986c1fbeadbf7", x"39e1183db6442602", x"75181217007a91a9");
            when 11736156 => data <= (x"035ad23ead3d620e", x"0c8c762373e55e0e", x"60209a518380651b", x"089afdfd0726feb5", x"45967a7644befe4e", x"0176e337d722f3af", x"8ffffc678081ef47", x"58d43809b904d861");
            when 8289544 => data <= (x"64d36d0c1f81e8d1", x"ecc64433db4c9065", x"fe8974706a75563e", x"879498b46fa23d56", x"3fa542a35582eb44", x"6a84b1c330445f19", x"d31fd806583e081a", x"133cbd74ed0d3c77");
            when 15680993 => data <= (x"70ea6a51405478de", x"8f5d4e86e8ab26e3", x"f806dce03a177fd3", x"978d6dc9ac869d3d", x"fb0254bdf1b191a2", x"61f841307982bd10", x"82f275a634a47d24", x"5c39dadc824bd71d");
            when 845997 => data <= (x"07919f02ec088aac", x"a584f48a884748b5", x"00ffb7ae28f07ee9", x"168096cef9dac4ad", x"3bfc8c0ac0e3e32d", x"33cd5818ee0dc70d", x"31c62f543a1ec393", x"2b424fd8dc9eb297");
            when 12849110 => data <= (x"f1a0d3bdc93b2134", x"9e2e9aa2f2296e4b", x"a88d55029876e703", x"2aa718447ed68a5b", x"cd12f3e18be62171", x"d057c4c9dabeb5df", x"b227f20e15e69afb", x"7602261e6d8a0842");
            when 20915454 => data <= (x"d6964d7b08e7770e", x"babadebf7e3846a5", x"6bce2910a0695188", x"e7ce28c4ac81aaf5", x"0a62f93d58abeb22", x"65187c87370a34ff", x"3025d60dc5b14d4c", x"a2d000467a475ff9");
            when 20661737 => data <= (x"fe881a4d7b9784d8", x"f5f465fc7a4cf7fc", x"e981e768d9314a45", x"5f9fb556565d2d6d", x"a9ea42ff3702d957", x"cda24f395ede0620", x"bf2d8200c24c701d", x"8b3e0b1fac322a0c");
            when 25430930 => data <= (x"7e6dfd731b7c1dfc", x"a06553337c4829b8", x"6f7eb34e6c708dc9", x"fa29d2e5e0540302", x"19771e94a6e9bbd9", x"b36646c948948f3b", x"43a6dbdbb63307d9", x"1c51fda83949dfde");
            when 6277205 => data <= (x"b4a6dbc578f71ebb", x"be95fcc409e39e1a", x"a0766be5abfa8360", x"7de1e2060a8ecd73", x"b66456ed3f303020", x"76d81197d91caaec", x"32f3f3a821fc689d", x"ba266e6de0938025");
            when 19076044 => data <= (x"cbf9adf9241dd4d5", x"79dcdb9191a2a5d8", x"d5b200957355d97f", x"dd45558c687bc8df", x"2e128f9b98f5b4b8", x"cdf9952079c8c3a0", x"f3fe4776b7782ce2", x"e3c684cf44742803");
            when 7394187 => data <= (x"9458e44e7581dc08", x"c052291d6a555c52", x"60d68ea483ae02a2", x"58b15f06ef0798fa", x"1aeda99ecd638a88", x"ec6da6d31f58ebb4", x"19cf537535cafc9c", x"5327eb956e1ee132");
            when 10983759 => data <= (x"a950260a4b5f49b3", x"79321526677ead23", x"d2cb5f8331b4e8f4", x"8efca6bb2791f581", x"10e73c5d42be6bbe", x"c2b8645e8d858358", x"9bffe58831711d5a", x"512835d3f269ac0f");
            when 594125 => data <= (x"4c0f9a444bf39174", x"3edc5ded40d5d744", x"5e2eddc1228d9d6e", x"5667ea491428fa3c", x"6206b59158ae1acb", x"56ebaa16232e126c", x"a4c11dfcdca0e67c", x"a26a90215ddb770a");
            when 19427730 => data <= (x"fa27ba7e6319c6f2", x"20cbb864f1bd0257", x"03b8b6a8e3b393af", x"81ebb905ccfde810", x"c2944760c953b825", x"1b14b4f7f3423903", x"8c6db2300aca346c", x"7bace1d6ef4fd187");
            when 23505672 => data <= (x"8856ccb6ffd4c6d8", x"8053ff7480ec0da5", x"a061a42549d7463b", x"813ab4545213a82c", x"e1d3ff57f959ac24", x"17a53a08f548375a", x"65b249077c6f138d", x"0cc9067574718143");
            when 19232286 => data <= (x"a46079f6456498e2", x"416ef3e8e57789b2", x"afecd828b6e6e1fa", x"c28cfe6b7da3793c", x"c3141e1f0f2d8cce", x"ca99432f3d6092d2", x"c95060db67123d1f", x"c0efd28bb27d8acf");
            when 8571350 => data <= (x"b52f39648532a5a1", x"f05d41b6607760d8", x"658b6db9416fd89a", x"5917693fd42391a1", x"de04268049f47f9a", x"99ecb08ed5f270e8", x"73cc86e23745892f", x"bba2f6737949ac3a");
            when 18087073 => data <= (x"69a3ef112cb16dc2", x"96e980d10dc9b1f4", x"d323d7a3bffaaf23", x"4f3422bdd38dd4f8", x"f34f3dac6e492662", x"5f8937ccebc09713", x"5987e3df3adc8d32", x"b6182d8247ee726e");
            when 31509968 => data <= (x"c8022b92b9fadb61", x"3905d9d7bf8e39fd", x"454b82be8f8a86a5", x"e353d1fc0f9b4e87", x"a0085eca70e5f1fe", x"ba895c6046c8ace0", x"92cf753b5f08b29d", x"4958762fe3ac7dff");
            when 32612189 => data <= (x"2d65adab1bc77b6d", x"f20d1bc3c41f7826", x"9bc7fd3c417b9ebf", x"f64f6eeaaf7ce9b0", x"df45f37f4ad94e9b", x"214371bf2304f995", x"dd9ababa5aca7393", x"611833294fe6d7cc");
            when 18732795 => data <= (x"4d24d791a578b0f4", x"f15fc124d49bf4c5", x"a154817d27afd9d6", x"ff9e0ac49f1ed44a", x"98c9bfa8c7cbd46e", x"240bb34324486930", x"e6a8d5f049c1cc35", x"fd80da1cac715ec2");
            when 18134559 => data <= (x"d62c168e6118345b", x"125dc213176d380b", x"42709bde79b53ed8", x"d6077aeba40acca7", x"4d80899ca9d05c6a", x"73821efad5d9111c", x"7c226193cb904587", x"ff81eda267f5fcb9");
            when 11749237 => data <= (x"dd2a885ee8ca9e37", x"9955d8f1152e9d77", x"e7accc478b870e39", x"1a008d8ef1ce91b1", x"1456e9eef9bcdb0b", x"0f33c27a8cae9f7e", x"ec69f6aa3663d7aa", x"3287bbee275399ec");
            when 6703686 => data <= (x"47ae2fb590de0588", x"23ce40c5526bc4b3", x"2e4e9dc652dd93ac", x"38373f06938461a7", x"6ecdc55181b203cb", x"233e46de09c2e361", x"14b0d67771b501ff", x"ce5fcdff54986aa6");
            when 12014051 => data <= (x"8e553ff858013ee3", x"ee7cb9da681d8afd", x"db84535b6dc16581", x"d03906ce8fe108a2", x"4b7f5558fed168f8", x"a7f6433876b7da59", x"de386dc417aec0f4", x"7a7e9d84aa7cb12b");
            when 31412467 => data <= (x"c71bbeed2ffd66fc", x"1b08b12d490db259", x"355b9871e11c2453", x"425b1cb31b65acca", x"53d6a1ccb0f286c0", x"1f1f5c95bd5cf863", x"dd7e6c7a3947b072", x"864e17df4d48418e");
            when 8329343 => data <= (x"e0031e4af63f3c01", x"f2d4162726b87505", x"199e7df0e8234c6f", x"f98921af984b7316", x"c1149c000b5cfc90", x"e50256e09bb68139", x"a4abefb0816e06be", x"561b07da3b68e03a");
            when 31142405 => data <= (x"f98ea7c8717e135c", x"5df735ca12e9c8fa", x"6b6f37b6ee051891", x"0cf431c31c94f659", x"f68ecd3585644926", x"2a29ca735ca58921", x"4cb4b2559ebfad48", x"317e9751d1a02892");
            when 8711650 => data <= (x"621f163a67a2196e", x"3fb1732a4f031a3a", x"b4a4984e0f384cd7", x"07b0bd4130d2ad9c", x"320323a8967f8fb2", x"aaa805c4562964f0", x"c1738c1ac6ea8e8f", x"d6f406b72881ca9f");
            when 11473096 => data <= (x"df206257ca0e7e56", x"4610a60ead76756d", x"afccf3bec404fb9a", x"dc3073a641daf8f5", x"05397f34adf8b3a5", x"579f0e6a390a6824", x"7990b9c5e3db6cda", x"7661cee8340b5061");
            when 806015 => data <= (x"08a3f4e66a4c7688", x"064647558f4b7301", x"a46b66c0e4a54091", x"0f34a31a90a43fb4", x"0ff728f130fd3f89", x"5fb56f76e8b87b4b", x"de2d8ee387516ee9", x"c925563b3bb100a9");
            when 22680745 => data <= (x"a71140753867bb04", x"b17ec55aa4bb4d75", x"262a723b7b7b9c9c", x"4518173887db5c19", x"be0832daa1cc0009", x"06582bd83570d3ef", x"4c43af108f6321da", x"4b135fd2e1a297fa");
            when 32982854 => data <= (x"e363fb0e6f2b4dd4", x"495bf295352150fd", x"0a28784c94070e8e", x"ca45a309b0a4f5e3", x"c82e79ac03820945", x"f563932e9babc933", x"9866c08149b4db6e", x"0529fef0d1bf17dd");
            when 31317398 => data <= (x"c16b00daac9ef70b", x"f519fc5481854fb4", x"36f3dba7e2bac187", x"90e61ee917c31479", x"daab5bfc955ce818", x"905e1d9b1b4cab10", x"f20cd52d946ff31b", x"95c252d79145f89b");
            when 25197214 => data <= (x"045daf4ec1a7ff08", x"9725b2404acacfe9", x"c0b54893c619cde0", x"1e34c4582ac3e17b", x"e3ca36c09e370aa0", x"e093be3a53fd79f8", x"7eed0faff046055d", x"36fe97e48c1179dc");
            when 25999014 => data <= (x"bf438ffd90fe7144", x"b632823306ceb136", x"328bd44397fe6b75", x"4fe17d8618ee3413", x"4558109448d8aacc", x"bc6e0bbf81911aa2", x"6c8e17a33ef53d5e", x"938cafcbfc606fd9");
            when 7111557 => data <= (x"acd56da253a1876b", x"661458a09e4fa1b0", x"e0c276db484606a7", x"97eda78be2aad9c3", x"b091f9acf1dace5e", x"899968eb9386bfd1", x"defe9c5f04f28fff", x"1265d50276224dd6");
            when 32746845 => data <= (x"af8306baeac3f6b0", x"6a360df53fffc838", x"ddec38a70833ee23", x"819b0384f75e5c7f", x"a11fdfe824051e97", x"de55cdae60d6e372", x"6811bc9a7111bf8d", x"a3fa47e8e86b528e");
            when 2717559 => data <= (x"957563848cdca36a", x"278269adaae2b4ec", x"1292ce0f8f1e45d2", x"e9b211b3d54922d0", x"2e4ddf6819b0105b", x"f1b7ff95f1fc24bc", x"e68f6205b8b67070", x"faa4ce6ae7af4f98");
            when 28653343 => data <= (x"97e139fd09a9620e", x"6ff24e998c097a23", x"9e998cd53e15d6ce", x"712da3cf1f687a7a", x"277b12d679bd5fdc", x"45eb0eee4e09ed92", x"86998089b2c49ab7", x"9a91ffb3e48a001a");
            when 18133568 => data <= (x"d517145bab2d04a7", x"324025065ee3c6e7", x"7897cfc8080e0afe", x"8501c805fdb28a79", x"5604ad409587c367", x"a7e893457fed0a1b", x"1f9406b7a65c5aa5", x"201230e0eca14527");
            when 6971464 => data <= (x"406395098f600873", x"6ffcf16b86b54350", x"de4dddfa535da6be", x"c11de5287670b049", x"a64ee74a2737e47c", x"44167b51dcd68042", x"77ce7690dd66d62a", x"3547e63c331b31dd");
            when 32185021 => data <= (x"f5159cbf755c181d", x"15552bd0bd171aa6", x"7299947dd61dfe9c", x"981de609b06e3e84", x"caa6579eecf73a96", x"2738a484bcf241a1", x"c3b094c242133bdd", x"482899b61937e614");
            when 28852301 => data <= (x"7112d4b2a47d8a69", x"6de3ed04bddf10e8", x"a945d0f104127458", x"47b002311fc32136", x"219e97b051d15cea", x"c9b936d2e595021d", x"4b5f74bc87561d62", x"4f263793662e5680");
            when 9925650 => data <= (x"274a464fa2c72afc", x"78ee3c605c0f8059", x"dea6712e8b583887", x"1e3a80f5168c99e3", x"27aae75e9ab3493e", x"c2623de5dfe9a9c6", x"aa37f2fe14ee05bf", x"5d7bf046142c68f3");
            when 3584789 => data <= (x"0ccfaa68ce4f396b", x"7de50594e7d690e8", x"179ffea62347a109", x"2007891bc4af2b3f", x"40d73c66996432db", x"d37ae6e68ed0bc2f", x"cc292d065e5fdbe5", x"a9949d21d50d87b4");
            when 9216323 => data <= (x"b8a9e12d192801b0", x"5523784dc7a53c74", x"a2c7869ef1649a36", x"913dd01ded2e78c4", x"dc164353121b9a49", x"b6b350ba57c3dd02", x"9a3373f818d0c0fd", x"4afe933a9acc2e55");
            when 4875168 => data <= (x"2cec1d545d7cd57b", x"63070f754a42ff95", x"e9968ce149e955df", x"c8f4b99d1dd92559", x"1a898f229f4f23d3", x"6ae4c8a4d505784a", x"d6edd26b0b4e9fdd", x"e528aaeef53b4c5e");
            when 13059786 => data <= (x"bc10b1fcf47f9ec8", x"01abc66cd114c2a5", x"ec3dd8ac7ff347bf", x"f1c6512ba4a8fa3e", x"f795598ee2ebb28c", x"7357ea5c7665c796", x"6d4137eebc76af48", x"a73214b6dc40c18e");
            when 30199068 => data <= (x"1e7386d207107f9c", x"1b88b263e787e8a7", x"621ac02b93c73bec", x"53ea067bee0a8908", x"23fee0e02cc3b66d", x"ea4ff44b692a71d2", x"10e3b2fe7c82c7cf", x"92b06b47bb9afeba");
            when 10408004 => data <= (x"65e1695c935537bf", x"94d81e405eede6da", x"b8fe9da7c2ea9cd2", x"1210d32d7938e96c", x"0b0bf662ddd8da9c", x"32e4e06852358d4b", x"99877b7c84eeb344", x"0761b0d5274d6959");
            when 9917082 => data <= (x"eea023cb7f45a7c6", x"964637698c64044d", x"e50325aa4a43dd80", x"d7c15209855e2e40", x"07af484b9420f3c7", x"4e5c5615dd7d0704", x"99e6a998dadcc621", x"e29565bc014637c2");
            when 19436043 => data <= (x"0aa58fa668811666", x"de7b2587e2b3074b", x"e3453b672b84ecf5", x"c68ec514ac71e095", x"b0d11167ee48586f", x"174b6a55de6dafc2", x"563a3dfcc42dc7f3", x"7f3859cfca4bfa03");
            when 30988109 => data <= (x"05834a19df4410cd", x"2bc3d8914d0b838b", x"ca95f621aa4e6f20", x"6f78f5dde74326ba", x"520d2bbd66d02a50", x"a50643e5ab590e49", x"a88396b86ec4fc4a", x"a1e4300563ddd7c2");
            when 14102508 => data <= (x"08addc404df05fb4", x"bfa8ee75c57f7007", x"837057e2e6142be0", x"2559421d67c9b6ff", x"4cd4bd9eb8d6edd4", x"38ba0cb7965c7326", x"a837b49719236a56", x"7935cfce6dadb470");
            when 23478484 => data <= (x"dbfd6898a2192d8b", x"e044a32e19f5eed7", x"26b10afb4e5e6d39", x"c7b466070e24386b", x"0b807b7d1aced072", x"1cad0199b3dcd12e", x"fd5f23775a99cff1", x"d15bcc05e331ae07");
            when 32780919 => data <= (x"e79818e5194e95b1", x"50d1d668e72a6af0", x"aee1aeb33b8da7db", x"de6a0051569ffbf5", x"809fa165bdf371fc", x"ebb98a29fcb9352f", x"44a4b858e1493c1e", x"bba22bb59fbc32cf");
            when 26657703 => data <= (x"79e5adae8bbb5987", x"336456b36e7fcf3e", x"a99b158e3b5896ae", x"5446b429a9ebe088", x"77c5048576bfe8d7", x"c40d477e97a80b21", x"9773683f44e55885", x"025a4646a3aa267b");
            when 16063107 => data <= (x"11d7a309bb298b13", x"3f4a9e7d63d34494", x"0cf72456e5cf7bb4", x"412a8371960de1ce", x"c16216739d23fc2f", x"e94d3c13884abb52", x"31f56d58ceccf3b2", x"96a6cc90324aa58e");
            when 6240094 => data <= (x"14bdf136b4b63922", x"5f589ae0e56598f6", x"f9a59ea3bf2fd1e2", x"b6c9bad37a1c41b7", x"fcf829910b17248c", x"93e29548f1e58d7b", x"ea91add864f694e3", x"4b6e45c33c277591");
            when 26611076 => data <= (x"ff0606123bd69dde", x"84ce672019a1eb21", x"c9e567af03987085", x"a0b36974ebd961a7", x"016e5e09c052a396", x"c7216ec690d10549", x"df70a30d0303b16c", x"6c15e4e74c01fbc1");
            when 23750485 => data <= (x"6d9ba0028457e1ea", x"708f0de0ddd39a50", x"39c8203ab856d703", x"99661cb6ad8d1a2d", x"a8e3eada0baa8cd6", x"c4b8f8913c9298ef", x"dd35e793b4df65dd", x"63b24b17a4c7ac44");
            when 13617129 => data <= (x"3a29e6b262dfb856", x"0c400fd0029a0992", x"39e8d0d91a40072c", x"337f6eee1be0ba9b", x"709a8889663978b8", x"9db4cdc7d70bb506", x"8550a0bc9347b44e", x"572c3f5e9cdb3e33");
            when 10766879 => data <= (x"6cc358bc2838c1e7", x"b26b667963ff029d", x"d3fd264901981d86", x"c44205b182f8b924", x"c80296536fa6d8f6", x"dd86552cb23f7ddc", x"0015af7db78eaa13", x"947e870d834c3cf4");
            when 7628450 => data <= (x"f7473ad8896e066d", x"8fc3fc4d6a086818", x"318b13be2b16678b", x"922e2b00e7f82503", x"b807a7613cd9bdae", x"36a694bb76eb7c80", x"3c1df78b08ab6f32", x"de8e7243f7551d7e");
            when 24211071 => data <= (x"dfb402808d9570d4", x"c39953e6f0ce62f1", x"d7480a68f38e4c41", x"9be6bf8a0c4cf1da", x"42efd96b2898821c", x"bfef0cdded608284", x"59b6fa6e41e92148", x"f90f8b983b2a8965");
            when 12812797 => data <= (x"4fc8df01cc425fbc", x"cc47945e0652fc87", x"38a11ae66c481873", x"4e0ab91deb6b8817", x"db12886b0672cb94", x"6f6a463a9f6a7f3d", x"d76e65d843e2b70f", x"e4079c56c252b2aa");
            when 5086656 => data <= (x"126814a98ac3423b", x"6ab5ae0e28492acf", x"daf22c800fd7dcf4", x"f6a382d8ec487d74", x"509cc99ef63adbb6", x"cf983f2f19baa756", x"f1b948c717b591e5", x"5fd0d3fc68d4089f");
            when 1786549 => data <= (x"3ec59c4e5faf9911", x"f0cbf8b9081d3bfa", x"ea6d477e8057d4c3", x"a347d9180766111b", x"c204d732996120d6", x"c00e1f3c0e5d0aac", x"9675e63d0b8a9f66", x"605bae88437c14b0");
            when 21332372 => data <= (x"c01eabbc6c11aea3", x"7d4762ff0cd4ca45", x"cddc4a7324809c0f", x"2d57088b4b350a0b", x"664e8aee728dd3a3", x"aa00d7c9c37a58c0", x"31165e46933e1701", x"4540aa4dac6a696e");
            when 26008043 => data <= (x"f83badb2a087b380", x"45c2e64c27b116b0", x"408371eac2f63991", x"3d0582d8a49946da", x"78cf24fe25011651", x"ec762830e4f1deec", x"5dbd94fb25674210", x"f96cb191188cc48f");
            when 9943952 => data <= (x"98c7c9bf5e233573", x"3af7d73e37f224f9", x"1157804b2c6e828b", x"351e09e777d2068f", x"537c028256d2bda3", x"53d39378a8c6b70f", x"4d341620effc43ae", x"75d3baf09dac9618");
            when 6338705 => data <= (x"045fba1dd65f2ec3", x"a9549efabde70215", x"b1a3c05d23caa527", x"f85ae89cde88bee8", x"fe33d109d6c85b20", x"a3228ebd583344ce", x"159a8f72fd545551", x"9950e4eb90f587b5");
            when 769238 => data <= (x"756db86da87b7e1a", x"3bb2e6842b7189c6", x"f55dd8e7c6b62e81", x"4a040a831cb24c87", x"e00b207160689fd8", x"85ade50750b877fc", x"3b1992432a8706ea", x"e5bc36b021c8a02e");
            when 7992429 => data <= (x"29a06b5a86665b72", x"929ea31674266c70", x"85a8dba0074ab0ab", x"f4ec3091bfcc74ec", x"d3ce7974181d131f", x"1471445d10cb3f45", x"a23d8aafb9cf9324", x"4b66f2ed1de5b0b6");
            when 5301970 => data <= (x"f751e3551bc04797", x"de5fe9ea0cee38c3", x"956ff2797efc6ebb", x"a20b2e2697c2bb48", x"66aa54ef1493e439", x"de148b3cd1ea3e9a", x"3317aee78b0926dd", x"64134513f2d8fe46");
            when 3053834 => data <= (x"1bf39039b8f15278", x"6d582088e915ef37", x"7806ba81da5ac2eb", x"cfdc436bed34aa35", x"45d3f9495f175432", x"15104b3c0a9f779f", x"3d9e7ce43a3827a7", x"18a5a987816c9741");
            when 11559110 => data <= (x"11358a4a9ebebc88", x"c898e78f383422ba", x"fc22e6b3b6c2381d", x"9345f30ec6c328b3", x"98d169bede441cb4", x"394f0a78def3bbe8", x"df6a01467ea4b17c", x"a7b201bfa128004a");
            when 31541314 => data <= (x"1ff09cb9f7bc1f6a", x"a39ec7dfce073b4f", x"24b132a30552f6b3", x"ff710350d508e84b", x"6704848ddf66f1e6", x"2314c77c56828038", x"9f3175b8f8471c8c", x"0cb1269d6f43b5d8");
            when 28390225 => data <= (x"ad08d5c143dd8e7d", x"d5808ef60fa2a819", x"6bae0d40a8fc220b", x"ae9caf3d3ef07887", x"a4cc31f1bea96ac4", x"6fd4ed641b32dd48", x"f3910b50ee10442c", x"fee9d9d3b6ee371e");
            when 16242989 => data <= (x"07ec76b707118e35", x"b3d4308057cda6c2", x"463ac469c04b7875", x"40c2d99039d966de", x"720a6c2f50010064", x"b959bb9551dc9465", x"458504a297cd4c4b", x"296fb0e2195acfdb");
            when 21123850 => data <= (x"4f6110a39e2b0989", x"2c3f20864bdcc8c2", x"96aef86821c32c7f", x"fe7e559ac87e562f", x"9e21e5487771f54d", x"6582b16232380553", x"263320ada36584e7", x"f6785556542f902d");
            when 4537681 => data <= (x"e8b07cb65e82c623", x"6a2c9023a78663de", x"190a0b0ffbb99f8e", x"80ab1f97c85fb28a", x"18c2c24827b3381b", x"8d95e15e207be36c", x"006f1caa3e07919e", x"90f443945b756c97");
            when 6549696 => data <= (x"efc35894f9210304", x"d14f64b1e13eb703", x"298a82d3a0b65613", x"7e1537279d8b3212", x"4b78a84265a97cf2", x"7c933db92e5e5efd", x"58fc9c023c437799", x"4e5cda47af279429");
            when 7853424 => data <= (x"05383591ee47dfe1", x"4474a93a0c9aba89", x"4a90fbe4c0ce4fcc", x"da7c60b7bcc1099a", x"fb732f8a43667cba", x"aae4138f32d7e51c", x"c77e4a54179db1d4", x"af6754e438c13ba3");
            when 10687550 => data <= (x"b5a5fa33d28f5ed8", x"f79abdffefc52fc1", x"8dad9617e16d51ed", x"17cae78195621591", x"0103ff20798c2e99", x"9ad73a06bea33cf2", x"a59c8bfa5ec5a781", x"d6d7f5cddf7b53c2");
            when 5427142 => data <= (x"2a0594a59d2909d2", x"fafd91d1c0aef437", x"91d1afd56b19b738", x"4773222c75f497aa", x"83069e3f4e952278", x"ff0ec42d22df6f02", x"d44bc0368f969876", x"28c913cd121f3c03");
            when 23905903 => data <= (x"cc60336fc088af59", x"be1c61f008909100", x"742592955ce323be", x"cd8d291b9723da47", x"78e2e3c5bab5dc81", x"b3d4c639db145af5", x"35b9720ade3ecf0c", x"01610f0c4f108deb");
            when 19990644 => data <= (x"86253cbf00838244", x"fae6dd7bd7e66766", x"e7c5de1a8c2d5497", x"db2f7f1c7a601594", x"ef6f5badeebb2d57", x"604850fba1bc9bbb", x"449b24324c2da27d", x"4aa2f7011806ebce");
            when 15162742 => data <= (x"34ed85efce9bbe8e", x"7b4f9c62d4d772c8", x"7ae7498a9a202f87", x"173e952b07b8059a", x"bca15a8653b55e55", x"e5ed567bd46d0d90", x"9ff3deb6e7be1460", x"44fde10117ea780e");
            when 29277341 => data <= (x"56933f8613356a67", x"22b829aec3e614f3", x"fa19ec103ed5d16c", x"7dfee23ace4aa54a", x"0c2ec6e583a6b532", x"a13b0c1f0608e453", x"6dceee93f59d2d94", x"d6b2619b8fe95800");
            when 1713877 => data <= (x"300ccabd0adc009f", x"834fbfe85ac88283", x"c8917270945f54b6", x"2d851bddbb1925f3", x"99b8a6400d977bbe", x"64774bf7217a5197", x"6fa98eaec4b8d35c", x"f484d25c3f2f772c");
            when 15657609 => data <= (x"b60c490d76370abe", x"a27357151b0de7a4", x"a27b01d95e732863", x"b35b915cfc694956", x"e0dfaa3e9bc31968", x"f63505bc09b5398f", x"4b05f344ab43c7f0", x"9ce9e98b09293fea");
            when 5592305 => data <= (x"ba1804dbc3f42379", x"d264cb13eab05e69", x"5104fa9f203cfaa0", x"ef9e58709f5bac6a", x"062468e549754b54", x"2c6b14b1baf75cc4", x"31cc8da060bb9c1c", x"6f4d4fac92432ea5");
            when 24127074 => data <= (x"9fd7d599f9fced61", x"3fc7c90b130479b4", x"e367ab70d98cdaa5", x"9ada9aad2d2a9789", x"bbe3422855a0865e", x"bfa99546d0c4bea6", x"b9f99b8877bea6e2", x"8650bdedca23e41b");
            when 15936338 => data <= (x"0bdfe2e81573658d", x"2fe7297617872c48", x"dc19aff63f98f3b7", x"4f42b95a98a978cd", x"e9f0d1c46a0c760c", x"a5568245e8da44b4", x"4b8f86fe9ff178be", x"bf5d223bf7b11186");
            when 12442453 => data <= (x"da254ce9acb6722d", x"476339e82d6fa42f", x"fe095875fa0bcdb1", x"0ee0561bd96fd8d2", x"44f056b3e2e1f0ad", x"6312cf48d6e913fc", x"fad8ed5ea44d839a", x"394ce4c58326d9ea");
            when 13406772 => data <= (x"f2e7bbf0538a3e81", x"0d53640235db5899", x"f39a61879327a3ba", x"15316b3c6373315e", x"91b02322abce7e2b", x"8d6a9ebbe1f7c0b0", x"f3550e70229b24f0", x"3725fac6b1a601ae");
            when 6902960 => data <= (x"ab4595588415273a", x"d8d471ebea585358", x"ebb4846dc0337363", x"56279d36d6a1a2df", x"83968969a835bc0d", x"1695a2cc606e9c24", x"694b00a62fae7a78", x"5dee3db58861b3b6");
            when 28421318 => data <= (x"73fa45117c3b0b3a", x"26c0185caf143c07", x"00bd395c7e7c7ea1", x"c99f149676a019bb", x"2fcc5d2852f9d91e", x"25dde851834cd293", x"56a863a58de819d3", x"d9b36dea1c9107cc");
            when 27704891 => data <= (x"30da277b6111dfb4", x"0ab91db5fe1c25a4", x"e84a28bdaa160ca8", x"bdbee04438cd6928", x"fd788826ce3b5a3f", x"f2444f093148701a", x"b35c1bbfd201084a", x"3425aa456886a3ef");
            when 2420592 => data <= (x"ecceb9a02511a6a0", x"eb3937d51072da5a", x"255dc4ac8f408079", x"09320ee413c69106", x"c6d5779cf5519a03", x"293139ed3f39fbf9", x"47176b94c623111b", x"f8f781d41920c1c9");
            when 33062844 => data <= (x"c4f54a82882e2dab", x"e891cdbab9e99ee2", x"2c07842b31c5b5d9", x"4839677af88d8a5e", x"14412f07268a670d", x"c8631396e8767ba6", x"23261b02ba980968", x"8f0bb2d4098fa1fe");
            when 30362628 => data <= (x"c1373bc7476c090f", x"99dc713e304f5e4f", x"5c73e35b6d7a19f6", x"3f6f35fecc99113b", x"1b6455a9556811a9", x"2c27308a40f808f1", x"8dd4ee6ec8623442", x"50deb42089bd1d31");
            when 24389225 => data <= (x"c6aea1e7d09af252", x"f342cb11a1309b29", x"77dc653d1feaf16a", x"a48f6dd0b27d310d", x"e74d2d054e512f4f", x"d18099d872621048", x"03f982e0ac3664d6", x"e6c6287a69f5e7cc");
            when 11213064 => data <= (x"2101956c58dbbb76", x"b7358b4682eee96d", x"8a52e771de69ca47", x"983dc9a7ba612edd", x"21698d83e36a6777", x"6ab0d0123e5fa2db", x"6763c1cecc54da16", x"9373953f06bd8309");
            when 32400044 => data <= (x"0e4b929ad3743a0f", x"9534db13d5b2cf81", x"293d97054b4b3b38", x"d2296ef1de053402", x"ea552c73105d0e66", x"f70b953e6beff55c", x"b8cb57343cecfa98", x"302fe454a7090d39");
            when 22800037 => data <= (x"39ecf7f0aeb7146c", x"a2bc0b05c5e48fba", x"a438e56a7aead631", x"d4702dc82c8500e5", x"47989b7f4067c504", x"562180c4a9b6123d", x"515378fc3bcc0642", x"4ae424083a16b7c7");
            when 24747655 => data <= (x"1e7dac62411200a2", x"4478aa07b6a178ea", x"47d6eaac36fe543d", x"546a06bad5c345fc", x"d9bd667acf7c8006", x"3e438a9c72846937", x"1285a34b514ac247", x"3c595739a61a655c");
            when 12291403 => data <= (x"68add477d1c02392", x"b0d86177e259b639", x"7e6a0b7575f1d197", x"16763ebaad96575b", x"a68db89f75d5bd72", x"ddbd58795e171678", x"224a23b4e1a2b6f4", x"ca9e48108b446077");
            when 22309521 => data <= (x"d1d055612a6d893f", x"17f76a77862bc554", x"1bd663530ead5abf", x"8c5278af32f5ae56", x"39040a7f8d43b278", x"ef04e7b37be1ebcd", x"8da237d8badb66d1", x"a692c08d912f3709");
            when 5192669 => data <= (x"b9c98faee8a20150", x"27f5ce633bc72438", x"04f7bc85b806d724", x"5a64b9d07cb49a94", x"db5a59fc8be7d97b", x"439323497f7c423a", x"509f0b2286c500d0", x"bc0208fe99a3b7aa");
            when 12341499 => data <= (x"a287c408f2a46f46", x"8bb22db81df1b986", x"e21e2b46d879b4fe", x"6278ee6f64e99a06", x"adbf859811e33ff0", x"a9e12bef2c103590", x"f203faf4dd69350d", x"c3de103b4c54c5bb");
            when 32041386 => data <= (x"07e598fc371c5aa8", x"7f0f2d857c3e10ae", x"4cd65b3c0f525774", x"2b0cdff62b77cac2", x"6780815129ae69f8", x"12d313c8db8f348d", x"4a301b81b9174de8", x"b6bbede744b3b0e1");
            when 20407659 => data <= (x"60c63e03523404df", x"8fcfe81930a60838", x"79d15f109f7090d2", x"712d096703a9af15", x"ed8df61c9b2624e1", x"fb9a6379c6514f36", x"6a0387d3930b16a5", x"4ffa7dcf397e30c7");
            when 17003018 => data <= (x"f9f00d072eae7ee4", x"46753d49fe8406af", x"da16f9f875febdcc", x"b50889560a03fa4e", x"af29339bee691b76", x"2393b3ae8bcd66b3", x"442bdf0c6a420171", x"9f8245bf68c88492");
            when 13559454 => data <= (x"db36d2e3002af5b3", x"5a4071c35d0a8c58", x"5f9c47028235f2e6", x"8de4bf9ab079117e", x"c40a014518511306", x"06a20098ab7a9ae8", x"1056aa78251bf766", x"55baa397925ccc97");
            when 23908512 => data <= (x"4403234bcedfa546", x"1ee3fed46e7909ea", x"87fdb084f69d3fd2", x"909a37eb12bd0024", x"6b76badb7b22247d", x"309a8038e2996673", x"6a0f9a5a2707cf09", x"b0c924c9cd2fbecf");
            when 24932369 => data <= (x"cda9055acaf45b16", x"0f338d8ef5980c6a", x"bc0f06bbf71d6021", x"5651b5ffaa9935b0", x"667438cb4e92627f", x"7ee6953426a686f6", x"469f04df5c1f50ce", x"b676f898e8ef4c6b");
            when 8588967 => data <= (x"75576d0752b704db", x"664731445a5e4dbf", x"f20b851d9f0b021a", x"b10896a4b417c6cc", x"5a098a994a0e1c86", x"95584c67ae37e38b", x"2cb5aa704eafdabf", x"4bed6721d03200f8");
            when 30213717 => data <= (x"2a63b7d3ff323b1f", x"f859209d0f44be41", x"988969aa4af41216", x"5be2dd618b0406dd", x"2327b36bb8b49edc", x"8b3059694aba083d", x"3a232afe89b90308", x"7191bcb6152d81ef");
            when 2744313 => data <= (x"7b8f1e18377464d8", x"3c73cc4920d64b04", x"ade953d1fc0a2e29", x"990c83807fcf7f62", x"2f3b148cb24f8558", x"6928ed13d728130f", x"a614e719ca45c371", x"f563cdb046685b19");
            when 13449420 => data <= (x"4d7cfa1ed54ae52a", x"017d406a674b3585", x"697d0ba5fc013115", x"c0babbcd20d2f383", x"8ba7a2eb7235349e", x"4ef2127081376054", x"3c29f0364623cda6", x"cc7a9a2f36432ffb");
            when 28780445 => data <= (x"e829aeab376c8b71", x"c341523fcd25bdfe", x"9c4701653af57146", x"d428902300524422", x"864a8a6ada8889a0", x"8c4f3306132f3554", x"c80860b88b60e5bd", x"8914ea3292bf4cb9");
            when 22260855 => data <= (x"2cff1abe50189f2c", x"d679a647f0038348", x"a2154eef96668735", x"c34f7cd51bb238a8", x"074e2782e6cb7591", x"7e43000204fa3ae7", x"2855a177f43eccfc", x"7cee621555630bb6");
            when 16369252 => data <= (x"76045d2da164cd78", x"ede7d716fd76254c", x"d1a8561e5a275e57", x"e5254e5111eb6b18", x"0cc52ec64a157b6e", x"97872afa9e649005", x"c6671b896ee1d037", x"04378e6497c0e505");
            when 2325893 => data <= (x"ef1e5ec830b664c7", x"8847ee676e0b1427", x"7bd8d42dbf069dc5", x"6b748aaa147694dc", x"8d9a2387f5b06223", x"2d643af2f19e887b", x"a275aa0951da268f", x"4ad50c5c73e9d8cf");
            when 21335534 => data <= (x"17ad2eeb38fe50af", x"2d4eebe415d5688b", x"7d86b721c956b389", x"c817dde65bf11170", x"f6500dd1c5aed4c0", x"7f7b380faa9dae03", x"01f5571163080211", x"14593508418f4436");
            when 17231279 => data <= (x"3299ff1b91ec2dc3", x"9ceb9b509c575a77", x"284bf35db83f42fb", x"cf28eb0960e65830", x"a2a05ba2def99a33", x"338aa1f79085ad58", x"39aaaaf89748cfb9", x"0ad4257f1ca6ba22");
            when 28089950 => data <= (x"d0ee730fd74be162", x"3a40c0274a04033f", x"60b6d5173ff3ba58", x"4424e96c44b7c0ab", x"fc4a387763b1e9ec", x"91e0d4e2e22d6e6e", x"8382667769c83d40", x"e8d4214e0867b033");
            when 28116793 => data <= (x"1d581f14b93e1a8d", x"8bdf8b30ea3f70c5", x"801265d6aee14924", x"64c0f336b34eed86", x"d7da068bcac9bc9d", x"8dcf3e1a2a16db5b", x"56f468da84c5730d", x"fc0347b60aa03106");
            when 26211598 => data <= (x"f5cbf83aa5390a65", x"421af1f4ed256e32", x"5fe4fd80592fadab", x"4df3c1a9e907bcfa", x"a3ad8643b2cb613b", x"ae1d9a9da985924d", x"d07837b6cde54abb", x"64dbf52a8b7f2b88");
            when 20103202 => data <= (x"722c81803d0b5a37", x"49938ebcb9849ee2", x"24c019f2e954018b", x"eddf117df078db15", x"4fa9980777b602e6", x"f462b4d07f676810", x"9fd528e6e8f98c11", x"0ea0602bbd79b397");
            when 12771984 => data <= (x"ecb8744b389c48a1", x"a3382025f4a5d7ee", x"60dd989535fd606e", x"0510ef528bde43de", x"48008475a6922c5c", x"1e3d0ebee149b64a", x"f9d169b14e3121db", x"c7fd9bc91081a214");
            when 6353993 => data <= (x"405bbd1beee08357", x"4f3f5508f77135d1", x"b509b1bb8fc2b82c", x"f363821007bfd4bd", x"3379a4394a076d1e", x"1f799d320e45a495", x"0c40cf5fac2136f8", x"631581635e1bce0e");
            when 2349861 => data <= (x"4277354a51e1115d", x"527c41ac417438a5", x"04dd7468dc2b3633", x"b6e81ce370f67df6", x"29d414a51bcf0af3", x"2dc4caeac50bb124", x"0462e26e202e806a", x"b461f7086d44d30c");
            when 26136964 => data <= (x"964d693afc834ccf", x"31184f5e9ab6a8e6", x"753edf6aacd08a90", x"b4b1550209f6dfc2", x"737b1999222793f0", x"36a0a11db9fe3076", x"9a4f4a68cfe25775", x"e4d799ad9c963f3f");
            when 31444642 => data <= (x"a8d7a6ae33f6c0c6", x"73c81914163152d4", x"b3a280377a52fcd8", x"2535502dfb15ca23", x"6436f0500ebc7a68", x"b9bf1d8b643a5fd9", x"7312b3d950862454", x"d2408af10d94f4bf");
            when 10280910 => data <= (x"4fcf1bc2473d3168", x"4780a7c36c5124bb", x"1ece973507ce6a92", x"bc159eb5e8da5505", x"a98a07e5fb14f982", x"a050b11b750aa249", x"c31867cfcefaecaa", x"1b37619132261272");
            when 10552981 => data <= (x"cc13ec8f54183956", x"9feb1ca69ad19b23", x"d8d62d1889864fab", x"847783b1fa631e92", x"3e54c3a61497367c", x"e0b7d907fcc3321e", x"21a8288067ebeffb", x"77841ea98c955f84");
            when 25125356 => data <= (x"7cc59c8a0060c920", x"c912ad93538abcad", x"94e0b559f95be692", x"18161993634cee2a", x"dd6e0746e018e0ef", x"f657899caa7b3cc2", x"1cd8cab7ffb8fe01", x"fad0ddfc7549db7c");
            when 32298488 => data <= (x"b024a54968baf27b", x"43626d3361ea829b", x"8ede7652f891a0f4", x"b3c21361fafa46ec", x"8d16fad1261e0f07", x"4ec1e57faad499c0", x"cb8cb5d2bb007dd4", x"c7a3f422d04c3e44");
            when 10923501 => data <= (x"e1fbf2cb5c81834e", x"ff5c149fd6dfb0f1", x"1e49e0f57558fd70", x"95c2532ce979291f", x"5eef9f881776653c", x"db75d77706099b15", x"5e6a7f5e3c6dfa9f", x"72e6ed292e9915a1");
            when 24270383 => data <= (x"2414b89b5a2dd4a5", x"23ab43863c666b85", x"322a042b74a20966", x"9b6d399c5108b91e", x"8003f1de01822aad", x"9232a3f2057a647a", x"1c0ed911a3ffb0b5", x"cc92ea54fd1beb50");
            when 23947027 => data <= (x"c323d4e9d31e6e31", x"172993452d7e9050", x"29514df79c18aa40", x"f0d48d8f934e5de7", x"52170fb0cf547f42", x"c1215fc98bf56662", x"99ad8c898c9380fa", x"0531b804803d8fb0");
            when 2405915 => data <= (x"430daf5c8f7324f8", x"564d26c4e91b6a37", x"eaee366370afbac5", x"8eb33c186a59e2f5", x"fcf543d0618bc87e", x"1d138ea909eed6c2", x"27a3dcf8c7344e94", x"ed7d3897e63c7611");
            when 26346489 => data <= (x"751cb9d4b62ba730", x"116b9c1e42e8eb8b", x"65646029f150cac5", x"26f89a154489b98a", x"012216c63e8f39ec", x"0d66769511c9860e", x"e9a3479cded2c744", x"850697cf50406b10");
            when 33331147 => data <= (x"05e3c12e454cd524", x"fab25c93d3efa7f5", x"c9cd6d2a7b1eba19", x"671638d81197f84e", x"7a5bf65bfabd295a", x"e07755c2d7a2b240", x"2f2f00ab986f17a3", x"9c1ca69a3cf5417e");
            when 30507597 => data <= (x"2d7dddba41526f0a", x"37b1c7710b96e1de", x"ce906fbbca42e100", x"d89c04d74e424f02", x"791c5eb527e4f404", x"f4fc7e534a69d930", x"0e3785613452a1f6", x"6e4926d784020a52");
            when 19112472 => data <= (x"08cb9b09e28844ad", x"122628efae8aedbd", x"62896fcbbf67b73b", x"e1653a8a479e9e31", x"c22ded6938667608", x"1ba494794ba92be9", x"3b7367844b0f4e17", x"7ce61dde9abc4cdc");
            when 22295889 => data <= (x"0172a1287330a1c1", x"493315931a31b819", x"239233d3b9cdaa84", x"983a9c535176cafa", x"b5c7667a503f9a23", x"5b1b47a07f594dcc", x"eb55e39dc6719937", x"18ee6832367239b7");
            when 11720607 => data <= (x"1372ded84f39c74e", x"2a5be82467f33077", x"888756f94921b4c7", x"1b314a710d43bd77", x"8165d2e8479b7bec", x"30c3b12a6a9f8132", x"3d23b43a32e525e0", x"e656972f59a4e62a");
            when 21055175 => data <= (x"3a797ad659123f39", x"51298dff07186c58", x"14a07836bdb4126f", x"dd9307d194230219", x"eedbbf14121c7201", x"297e58a77ef5dfc4", x"98306dcf9ff2f903", x"a83c47c961d58585");
            when 506854 => data <= (x"31701e15c888a6e5", x"4e49b9e88d1afb57", x"4b59bc5ba9bac378", x"077038555ea770c8", x"947a73eb1afa271b", x"f49074793ae1b55e", x"33dea45f6b0c9abb", x"d46085abec3b1899");
            when 408123 => data <= (x"d408a58b7784cf5c", x"fc75c86bb414b281", x"03e4269126175689", x"5a8479a1c443fcca", x"f83c5b7be1081961", x"4f17e533317b0375", x"1043c0ea60893125", x"0d32af4f1addbcd4");
            when 13427768 => data <= (x"d12ea4a947b01a50", x"36563a80085d7041", x"68b2a422d949be9e", x"f44427d8df043226", x"f315cc9794b1cec7", x"c7fa78775f4f5ea7", x"18543c4f6d44eb5f", x"6f457850b372984e");
            when 30490596 => data <= (x"9e08c669e2c90db3", x"348b7e82069f44a2", x"702b751ac7c26e73", x"98d2db3a03548a3f", x"06ed354eb9a64e09", x"63ade835b31a0e03", x"5389089dffd121a1", x"aea32ff593facc64");
            when 2624662 => data <= (x"32cc2d8a399cfbf1", x"476c6782eaa8382b", x"d3846baa58d7a0ec", x"281f19b2baa9fc06", x"ec62a921687e29f6", x"0ccdf66f7c0b6140", x"0b785e49e80c5e16", x"e4aedb9a3a7f9c3f");
            when 22217333 => data <= (x"d45f1f71d64aaf2c", x"bb87cda32e72df93", x"5e91a75a55facb79", x"ed722c20c8921cef", x"5d8af51e762c2815", x"2d9b6cee77d35367", x"8e54db141fbb6d93", x"e04d6b1cc8ecb679");
            when 16622719 => data <= (x"e979e7fcd8902ed3", x"3d703324744d6046", x"632b0b0c27cddb21", x"4a8d5878a359b291", x"e2f60ddb0d7a08a6", x"55c185e6d05eaabd", x"59c05cbadf89ce78", x"2a00e36a4e822f37");
            when 17025526 => data <= (x"762d21edf5a48b7e", x"13fbabd20fcfd497", x"9d4307b8cb9a0585", x"2a56036c0288d2d0", x"739fcecdd70545db", x"cc457081b5b54211", x"05e27d2435434c44", x"a2cbc5ab03bed786");
            when 23149953 => data <= (x"5ee4564016f83afe", x"6cbefdff130c98fb", x"b0a3a87a45b7b199", x"61fdf1f109391d82", x"4ee9fa2896a3ce9b", x"d27bfd43b4ca909b", x"17251ba1b48c381f", x"2799327c2a8c12fe");
            when 17411779 => data <= (x"cf453ee366e0406e", x"5c385ab51d3e00df", x"1d55fd5a81c3fc73", x"bd1b4dfb56c4986f", x"41b269e9e8d74a73", x"5c3b4cc7bcfce531", x"7a3f0c2677ca2297", x"30309d132d01b5f3");
            when 9021307 => data <= (x"bb706aaa556e0a0c", x"8f1bd91ee050431e", x"95b191b12bb55c80", x"25c25864064c1e82", x"5b6eaa093e25a9d5", x"434f300ce9778cc2", x"191f945a41f4967a", x"f217712f6181425f");
            when 3791294 => data <= (x"351fe00ebabf193e", x"6563cc114e915a2f", x"f756106304249eb1", x"82cb9685bccf4666", x"3611b62a95ccad9f", x"9ee294bb683338c2", x"895a2735773f5aec", x"649c710cf14292a7");
            when 25041824 => data <= (x"f5e216c683d48a78", x"5daaad05bfd14d4d", x"68c149ddf63a43d3", x"b100360836319243", x"6440363d1dad5c5b", x"5b22134f4c16252e", x"12a2b42690b11142", x"b42fdb0270f4d036");
            when 32576561 => data <= (x"426b85d66bc548b7", x"e2f0df84a29bc5ff", x"2d0a2b84ed231c7f", x"86ea6992a52d9684", x"61b2ad96ca1d67c6", x"0e576b30bcb43ab9", x"c094f36646508525", x"45c088dbeb1937dc");
            when 5025906 => data <= (x"f1f7e7798115771a", x"a91e4bf73956e3d7", x"0039d299ee44fb55", x"8ed08f15e4758d90", x"c1a8a7ca59a7dc08", x"c140c18f0bb41896", x"d57075fe890947a1", x"7c85585539306f7b");
            when 10138253 => data <= (x"5ccaa8bd905157b7", x"ef6be3dea6f2fac0", x"f26c1fb677560023", x"17ce479b60a7df9e", x"95bf66d056f81324", x"606c625b22eae4d9", x"0c7132002cd70fd6", x"c8899699bbab20aa");
            when 20659442 => data <= (x"3d479b5afa38d950", x"1d019846411ec723", x"efd50bf9f1e15d13", x"02e9c4e6cc6eea64", x"4abd81733dd0b9fd", x"6c6316aafa1d4868", x"2cdb7636815da5e2", x"ed7a521f890af300");
            when 24269753 => data <= (x"0a0b4fb45e04ee1b", x"628960998b692ee4", x"7a584b5a96900930", x"60ac7b460934ccd9", x"44deabb0898b7b9d", x"735bd8b4a161df61", x"5426dcbcc9b5832f", x"7c8ee5c81ed9a72c");
            when 19394850 => data <= (x"9d837f73c43cda89", x"b82e19bfd58d7fc1", x"2381a0376016e482", x"a5a72dc5743820b0", x"62f3c92f4dde8d45", x"edb3fb209fe5c47b", x"4fef8892a8cf9bfc", x"b9d7d429ed365d27");
            when 16296318 => data <= (x"a037025271f3d7f1", x"c07bdfde26b097ee", x"e1ecc0d9f55fd5c4", x"ba593f565ce63c1a", x"d2310330f0610e72", x"b46d2b7d3f9306cd", x"3e227ed7e4350ab8", x"4738ab6063e8acad");
            when 11495020 => data <= (x"54e2489ac51b81df", x"2287d9bc50bb75df", x"660da30950e0f8b8", x"f2279f4dd5125652", x"a7ba10d52b766c40", x"4f9fa64e451991b9", x"1beb7a4217b5b6d0", x"083637f062f12c61");
            when 9724769 => data <= (x"e19e4c2725afd029", x"9a03ca7d9c50de18", x"f43db48cf55dbfef", x"87363f963ff1b276", x"1c434818fb520026", x"c6e5014f560929d4", x"7e0e1fc9b6f79b0b", x"953ab52322daf4cd");
            when 5213105 => data <= (x"8996cec0d14994a3", x"f5ca738e2da760f3", x"cbfbb9f7ba4a6919", x"d715c5f33cc4bace", x"413c762adae1d593", x"acf6627a08305cc6", x"3b46ec121c7948a8", x"7baa14ea69659b04");
            when 22501077 => data <= (x"80b36d77e09972ad", x"51da8aa20c715a47", x"b764a215e9ceba18", x"512f862bd9ffea41", x"e2789586af84e2c9", x"cd55927814d8ae43", x"bace1d6b9edc070f", x"10b9b3eaca8fcc90");
            when 28790434 => data <= (x"0b727f575e983b4b", x"b5f09cd2ed9fca2c", x"944d544338bd38be", x"6bc073fa13f09b43", x"ab540548f4d88a10", x"f0c092521a82a3fd", x"3037bc6226a3bc20", x"d940eb9ce690a059");
            when 33423090 => data <= (x"67ba7eae1234c101", x"ae50fb0e6a92801e", x"12e1dc7d33bc2acf", x"51c11a17bc50d80a", x"ba6f3ddd5af7f1c1", x"7960eb37de26988d", x"df8ad985242a334d", x"1051834ac85b5728");
            when 7385108 => data <= (x"c4e37f067861fd8f", x"159f062d2588e270", x"454c17e00513c3eb", x"08dea4774c732db7", x"921a06bf6a935742", x"2f132e30f2c7698a", x"f27a96674293259a", x"794579e9c40e545d");
            when 26942197 => data <= (x"4dce7bd7df02f1f0", x"cc5a8a7838bdb049", x"ca5f480de59b8b9a", x"236ba2e2eea84f82", x"8b7b3b564f097922", x"3e0e38188bd5a678", x"33622d9182ed7e6f", x"f989b9c7f7ac3dfc");
            when 19310008 => data <= (x"116d84abf43e3239", x"c0518e544fa7d6d7", x"a0a1ddc348281e73", x"71eba158e10b9482", x"a0deaf5784858a37", x"49838b4a271ddff0", x"6b1bfc2811c0b80d", x"45ffa47830fcbacf");
            when 32652282 => data <= (x"ca2b9e44c4e36972", x"1d329bbca44e7c92", x"43f6494aca2a54d7", x"50adce333faa0ebf", x"be72692ea22aa912", x"9fdf55a4c5000b6b", x"c43ceeac97c51177", x"53580ea1469d9680");
            when 11111559 => data <= (x"83461440942b3fc9", x"1699d2d80c75b9da", x"4984f2c553c66320", x"40a91aac0bf85abd", x"b621826e4986f773", x"f207daafa24d4752", x"76c0da397d1c2e44", x"a93d636b77798633");
            when 23258086 => data <= (x"79c8d931f17237d3", x"f0fd0e3bc3d60191", x"5587ddc067b1bcf7", x"fc7753105025ab15", x"c278c0eaf1755ca1", x"6151c6ce999e51b3", x"6fcaa890d8dba5c9", x"a2b365d2bf03f9d8");
            when 26201624 => data <= (x"59e1689fa88f2b85", x"7d56c4a034e79457", x"4221f15d56236136", x"7b464940ac924119", x"ff1a497a65de5366", x"6f92d6d0a1b9c6a5", x"8172d1bf14daae7f", x"5f8f6fa281129c7d");
            when 1859086 => data <= (x"5fcbcbb4ace279b7", x"f81f68c1dcee844f", x"85d15cb80e293064", x"56baa1fee31ff400", x"27f59d1210401a9d", x"9c2abc3e28ba8adb", x"ec1f8bffb2eb01d1", x"4d2b497b055f1dc8");
            when 17962477 => data <= (x"8f724098a7fe1bae", x"296bb586f9bc03f8", x"2bd029398ac2a60a", x"5ebc6c0c5074ab22", x"ec0ae7bae5b8b464", x"4aba3f062ad15302", x"53a4899c55064f12", x"e2cbcd51730fb0bc");
            when 17846159 => data <= (x"1705778a770854ee", x"a080affdf9815ae0", x"3d26ccbb3db3d31a", x"5a527880c2412a11", x"9b4a58a6e7a3e8cf", x"e0ea2384e547fb15", x"cd51b1dcadb1eb55", x"d30cc56337e1702d");
            when 9654495 => data <= (x"8125f2bbc9bd7ccb", x"8d07c5bc2e1360c1", x"b7af94e8367b0d6a", x"d58b9c51877cf53a", x"7f821aa249cc80db", x"dd3715855e434332", x"362e20dc2f6188d9", x"d85dbea66aae17f4");
            when 15431996 => data <= (x"d9841907fdc2099e", x"1f44b3df24cbb40f", x"5bb2ce8c4a9a2d95", x"5d42e0f33e09a8d5", x"90832dd6f61f4893", x"c60c6945e908e683", x"6e110acfec07fd3b", x"c46f766c8a5537d1");
            when 31895448 => data <= (x"11cfdfc0a89890ae", x"c02826f0d310a78d", x"d6d2410653009cd9", x"8371190754ee8aaf", x"026acb213dd5979b", x"b39609dbffc2ca30", x"78d0f4cc3b1df017", x"9a711337e44a80e5");
            when 18332189 => data <= (x"adc8e5632178e03f", x"f4e31e04d972d55e", x"ce05ff633075a8d6", x"b5a47de316543cd1", x"f60413efc468ccab", x"80361a5e7ffb0d07", x"0694cba6460dbdc2", x"e0cbd403d165baf2");
            when 15840373 => data <= (x"de36926317f12660", x"0d93dde4f08cf395", x"09e7ac2392fb0c11", x"f1fea7506de9c145", x"6e5320e730078831", x"5e0f8b49f6332abc", x"20b8326a0fffef78", x"f4e9167a585e941b");
            when 26277941 => data <= (x"9dcf04592847c6a2", x"d04c63cde604f42e", x"a637d333822408a7", x"3920b53427752669", x"e2c57feb61f3cc8f", x"4983127e9942f4ab", x"33fa9f7f912b0be2", x"40372460048e79b3");
            when 24591198 => data <= (x"a72c8432353d3d2a", x"00b656276abb16d2", x"13f2b7d1bdd8724a", x"cd855fee19e65332", x"c71c179ba30ce92f", x"3b3b325e3aa7c4b1", x"956d636cac52acc4", x"a8685001eed75442");
            when 17940746 => data <= (x"dec707262fed91d2", x"d249d71989fd16a0", x"14c8ea716ac62c04", x"032c22963005ecaf", x"092469829dae4c80", x"fd7ac08108968222", x"ef72eccb2883ec25", x"f1da22af29d101b9");
            when 25415233 => data <= (x"4ef696df56c0049b", x"1d100adc73ed5679", x"e681a7565b261c98", x"ecc99892581ee2c2", x"0190044f57728ae3", x"25d491aba6bf3c06", x"a2d9db1e3551d358", x"8475503853a32a99");
            when 24058945 => data <= (x"c8f4e4c555527b38", x"78dc3654098ce67e", x"7a5dff2f78f28f83", x"7d8af51a9b626f50", x"8c1ee9ec4513bec2", x"e1e8896a7c175996", x"a0c169295b7df02f", x"06330dd95ea1eadc");
            when 20702455 => data <= (x"9433304c7a2efe92", x"c7dcea02f9414cb7", x"c160cb9375354259", x"3703e63f19897669", x"e3e5ea0a3eb091e5", x"955ca379d6cd703a", x"09a9a9fcc2d97753", x"3997e2c11fd109c6");
            when 21575882 => data <= (x"23360577239228bd", x"c1e3552f18a245aa", x"ca06994fcb934381", x"8f45230c7bf06b49", x"f2e3b1da4666a7fe", x"ea7f11ea9feca2e1", x"f2883afa759c51dd", x"f5ce518b18ec9f1f");
            when 25701852 => data <= (x"b3d3ec95cb8ca281", x"a209147ddc0999cc", x"7a4e84c5a34363d2", x"3cb7d27006162178", x"633261782ce312d7", x"5e864a08497e318e", x"1a9ae477185b19f4", x"5544fc6c2c7b8301");
            when 10185519 => data <= (x"bd90dd226649f29d", x"87786c82eae06ede", x"4da61e6b8befb6b8", x"26522166ef0bd616", x"bf36ce06682b2563", x"edeaf006db9e40f8", x"ca3f47bcfc8d0bdf", x"da7cdb6d778a4e03");
            when 30480763 => data <= (x"753a9f9db4dd51ab", x"07ace10eba41749d", x"e0532efc32ff9c10", x"a6d6a5d0f1e04143", x"dd16cbf1dbbe2f3c", x"cfcfb1f0480499cb", x"17dba3c965ef0c2f", x"32cb720ae4fd532f");
            when 17277775 => data <= (x"614e8ba6e0bc595f", x"57697c87fd5a0b08", x"7a48de2958b1bcb1", x"3a184963530f4a8e", x"a301184f13a9762a", x"1fcf4e36dd742d3f", x"1383479ee22c5eaa", x"d8d15f8fd2eb3aaf");
            when 18258055 => data <= (x"ad13f5e4d60fa9d0", x"03d384798113832e", x"2940cb5aa16fc757", x"63cf3b5fa8ad402c", x"ffcdee201b25149e", x"598f8f69e6994383", x"05b96dd47c723fab", x"ba2c5fbb8d44950c");
            when 11142110 => data <= (x"1005c0a7723d15b6", x"5365b7072174d33b", x"fd452ff9af5c6ef7", x"d2ed407348c9a398", x"8ff553759d06e95f", x"6e6eb61c1b1bf7ff", x"f93782180db62623", x"59ee3f7acdd9a1d5");
            when 5074760 => data <= (x"72dd60816b110708", x"fa46d171721bf3e7", x"fb52809cb2ccd3cb", x"f473c1eaaa44a898", x"28f5d55012099937", x"15f355c0b075e7b8", x"7a1032a8cc4c4837", x"6df6e0c5338fb308");
            when 22046929 => data <= (x"7dcb4b19a96e2fc8", x"d693643ab855b8b7", x"a91b2e317fc01132", x"def7b3451a64743e", x"2ef549de019de34c", x"be063f3c4b22bd50", x"14b602a00f2c5b6b", x"108e0bc85794f359");
            when 28590569 => data <= (x"3ec2918fd8772c4e", x"e3bf1181ba7dddab", x"4bce0822dd4d86a8", x"f87f1455f012fb6d", x"11b4852cdf64e741", x"62528e839f985150", x"28319a9dc5028d61", x"025cc44f0a54bb57");
            when 23685039 => data <= (x"a0f8451c0b04cbb2", x"70b5f0a799954c24", x"ab3757c5b6028c6a", x"8611e7a9db9d1dd1", x"4c2af1aa23166914", x"18bfd04052b3dad5", x"a50fe0bedb4fd1cd", x"eaeeaa2615528023");
            when 27600004 => data <= (x"38f16ec66848e49f", x"2a5cb62185e54364", x"59cbb3bd9b84a6e0", x"13f274782ef75cb2", x"39379a8d25279343", x"0063e400f1e8c9fc", x"fac7b66632a3c5c4", x"34dd0eddee0551a0");
            when 2148708 => data <= (x"1821ee45adfcd6cf", x"148ca9e2fd7ea7fc", x"e70eea5c891ff319", x"23613bce509bfe8b", x"a0ab0ea5235c0dfd", x"a0df914dd9020478", x"cc4a1f96546ba3ca", x"4c0f65e230b01489");
            when 3402941 => data <= (x"c222b7f7d6615838", x"338f7bd7487d19e1", x"7ffcd9c1e0fba321", x"70901d477e8107fe", x"9fa18a6ca06f4228", x"a2ea0e82d076cc05", x"52cf29a503e76f40", x"96aacebb49a85c78");
            when 8667693 => data <= (x"dc60113c3030f5d5", x"51493007dcb2eaab", x"9d59893ee2ffcdfa", x"6d8fc6ae465bf544", x"6b2357c1dac0f4f7", x"ee57d9101d65f7bd", x"2e63faf7d158ca3c", x"ecc8acd595b912ed");
            when 2200905 => data <= (x"69df05c4664c178e", x"fc07baf3e23e147e", x"532cb6381f0544c0", x"0468962395178fb4", x"3d32a57fc5aaac1f", x"a6a47cf0d2b03e7b", x"585234c3ee3fc2e7", x"1b1d4ab8a5ad0280");
            when 29863357 => data <= (x"75470cf4088201be", x"3c1a88df4b9fdc5b", x"d9beab755993f8d0", x"c206eba83196dfb1", x"7e2d9499c390c5c3", x"623eedbd2fb0714a", x"9529eed9600f71d6", x"8a1dfd99e1669e93");
            when 32919616 => data <= (x"d799b08b29352f2a", x"0ad0c03da1f26d67", x"c92a66aa6e40100b", x"e4e74f2c0f5d6121", x"eb7a427dc53a2043", x"cafa9110b23ef34b", x"635e7a04f51519ed", x"98751e6877fee058");
            when 1178462 => data <= (x"abf7feb1b6f992ca", x"d231f62d2444d38f", x"e2bc5f09b4bc0ab7", x"380d4e15ec15af7b", x"7f76622e889e820e", x"d7ca0916ca510f18", x"128b160a8f710bdd", x"0ffd725c6a091a1c");
            when 29876451 => data <= (x"35cb6752429df7ec", x"d70bf8fcfeaa742e", x"9e83c054098e7d63", x"4a6f208f6a58e430", x"fd9dc5f38b47067b", x"cb1a8ac532c6548c", x"fffd5505116476db", x"fd3efdd4c849781e");
            when 9404776 => data <= (x"3cdcff243bfd7d3b", x"0b77faf22f79e4db", x"7b024f1aa70499ab", x"f1e307d56a9ecb25", x"e76f4bc59a028989", x"71c03a930b91a6c3", x"7de229299120cf4c", x"4dd1ea586aaca40f");
            when 5644509 => data <= (x"a3291a7de886793e", x"c9d2b43ad4da9f69", x"4031dcbb30a43234", x"e6b22953da34259d", x"ecab67968cd58cc0", x"072d62f3ec2cc22b", x"ccf65b307abb3914", x"acc6400e634cb93e");
            when 1146690 => data <= (x"41a474b3484bbf75", x"7eee55ff00cd73ca", x"fcff76ad83b6dfc9", x"92a3d14535a12457", x"ee2a1c14092af808", x"b5c493ccaa82c721", x"314f5536838d38fc", x"67eb3a3073bdac23");
            when 29123161 => data <= (x"101697d4c7015839", x"5187049c809b2246", x"d03ee85396a3b8a4", x"78ba24324a363f23", x"ec7641bfdb7189a1", x"b49c0555f6400552", x"ac2ab55d3ec038bc", x"70d765f4ecf04cf9");
            when 19552008 => data <= (x"4af3e5906b2e715c", x"fc73b44c1f85b3f2", x"c51b0b4e98a2a7cf", x"fb884b2597634c78", x"a63d3c7ef6c3e7a1", x"ea4b7977950b07c6", x"72fef41f5c7713bf", x"e8bdb66dc9962171");
            when 6814654 => data <= (x"55821d65fd4e0a5c", x"587643f7b7ae4ff6", x"6841302963d62093", x"67537ebb56e7c821", x"4aa8605f005855e5", x"33f35b7062603efd", x"bbaa2d5a3e121b1a", x"812d8db0762b9126");
            when 16064523 => data <= (x"f36316a82702e241", x"e3a612c4cd749a8d", x"4f921d81dad7e166", x"3c71295a6373c3f5", x"0ac4b37c8877a426", x"52ddac31b978ee8c", x"f0469131025e315f", x"614bc32d2dd7bf1d");
            when 29413160 => data <= (x"d982dd2c37b768cd", x"d7cec4e7fd602f1a", x"2bb7841d998c5863", x"0c3ba55e9822189d", x"691ae2889d8b01de", x"92a9a0a25dc7979b", x"66ada642b65df3ed", x"21431cc2126180ba");
            when 32802705 => data <= (x"cd3544cd06bd1621", x"bea178c88c08ce1c", x"f8d41f179260bdb1", x"0749c811c4bc6ad9", x"43ebff21412a62ca", x"c203b5ac7b0208a0", x"1be8bb12dd5e56c1", x"0905f2257784795d");
            when 598246 => data <= (x"71838c36a3a47a3c", x"c80b58b01d63769e", x"c9de283cc27ad69a", x"56f415cc7fcfe4b4", x"bcecb322de636ec0", x"72d2724c23e3bd54", x"d8f4c43bb1958942", x"5d45ca7083e54159");
            when 12285306 => data <= (x"df1abb2f5d8f3618", x"58fafb2c9a0b92bb", x"5b3b058379caeea5", x"98ee3ea1490d2254", x"8a3d1a47e66b1b47", x"babecc5cc9dd6a73", x"1d5aaaa635d1ea6f", x"9dac0fd9c68034fb");
            when 4167612 => data <= (x"f71143c8d8086da6", x"d7b4931dd89d4ac9", x"413ae75679d2771d", x"9c37f2f83ed834d8", x"4e7f5ad6b8d7cced", x"6d395e48072c98a2", x"6170fc3a6cdc2ef6", x"a4fc167b13fe23f9");
            when 30583111 => data <= (x"8aed840225727693", x"c34424f329d1e2d9", x"27b3d54ef6b0af3d", x"3066895df3701d42", x"58601c5838755c1d", x"6b1c62b0bd96e0e5", x"56927bb383a4f413", x"1937202a4d4b6536");
            when 22493096 => data <= (x"3cb072e398943a32", x"91bed8dc0bcb28cc", x"710841a6dbcc4a6f", x"1e21c3d8e9ec5c85", x"b06f0a73cb01f082", x"d3618c692ebf96f1", x"4c30a510da06dd6a", x"588da84be41bda41");
            when 11093130 => data <= (x"a9dae4891ca6625b", x"fbb9f9add6d8d679", x"2a9e49eebdffe6da", x"c4f470f35069949b", x"31f5af6ace0c97f7", x"30f771b2a0c85426", x"f427da5700b437b4", x"0eef50e45658dc4e");
            when 12714851 => data <= (x"c18c8fc95751b132", x"fe773c65bc7ac81b", x"885a5d9a09c7cd0b", x"6c5f12510ba8a917", x"862dbe84431ac8c9", x"269b1ddc2b9fe5c8", x"297f7074b8032f46", x"63373133ad194a42");
            when 6785985 => data <= (x"0af43cd601190b6b", x"0a445ef419031e18", x"5d2251b1d6856573", x"d70c6ffa529c860b", x"6875b8458ef0a659", x"fbd54ebab5793ce3", x"1a65cb8493f8869c", x"9cda0bb7f20d0642");
            when 26828676 => data <= (x"5bd2789b1dd66959", x"733ffbc78665c8d9", x"c219b87a94b1211e", x"528f5aa72d62da4d", x"5309c2a62783bfa9", x"9975463891049ae7", x"5c18e1ef5c4b956c", x"6bf6d3849d789f7a");
            when 30389326 => data <= (x"a34155fe76474aa7", x"f2bf98222fe9723f", x"58880c0bc24c6f86", x"09eaf2cb1cc041a2", x"7e638458a5336636", x"3191eaacbc1950cf", x"439241bd71fa10b2", x"556fcaeae27e2b9d");
            when 9198892 => data <= (x"6a1f3824a2bee1cf", x"a7f747627cca8463", x"ce40f6b242ccae38", x"9954a5a80b50caa9", x"ceabae6ae7e06b86", x"6ef1eccce4e3e0e5", x"10e6a5b2173319fe", x"b8e546db3b97b9d5");
            when 3499417 => data <= (x"1e986724f2b27148", x"cb828ed6bab21d1b", x"f031eed54f39be7e", x"b65c05f9731440dc", x"c4558111d2408300", x"99038f3ab9cae7ba", x"88d4aec86b707edc", x"7eff7636aff41401");
            when 8650697 => data <= (x"b0b57ffa59219c18", x"461b0686651cb3c6", x"19da0ab994e34ae7", x"9be0434bf19065e9", x"4499ebb638506b0e", x"a8d50724e12e8443", x"2c1704c638a2ff4a", x"71f6cc236c58d29b");
            when 14701326 => data <= (x"b7bc300f9c34b47b", x"c65d1f1b4f4fa71f", x"1e57b293d03a4902", x"5b4e66cc844826a6", x"537d1430b800a6ea", x"866bc2fe8b8aaf5f", x"99b808bef0ce8e34", x"019ccfb49c71f528");
            when 27844105 => data <= (x"af39e47bff3829a2", x"4f3bf265034d54b1", x"f16098c774884418", x"98fbd3641b96fbaf", x"e6eadeb2bcf9fb35", x"4e7a977a88d8bf87", x"8ef9fd5e9d4e5dbd", x"e915cb52afa28c80");
            when 14378501 => data <= (x"d08baae22b8672eb", x"71258c77c9a3d30f", x"3fa0790fb2fec863", x"b82f56aa1e681537", x"c9469950071a2d74", x"0a0c026d5800d7e2", x"ec28ee6d048de4f0", x"e11199fa0858ee4a");
            when 7180695 => data <= (x"e7b7a9ef1f0b8ad4", x"c78e09d73079e21e", x"b41d2b90ed10bb53", x"4d741685faea827c", x"8d84c8d6347b9cfe", x"a661819d56c86b1c", x"efa301c66d26ab52", x"8442040f31b89043");
            when 20970486 => data <= (x"0f47809f4ca6007c", x"3256a3b11a67072c", x"8a34c8952c8871fb", x"32eac6b5c0a98006", x"45a57cf3823676b3", x"5f80c36750225373", x"0e0ee0751234e1d6", x"67d2b436637ce9bf");
            when 22450945 => data <= (x"d68ad9b20c302ee9", x"b6a696359de92426", x"6f548634677cd1ad", x"11b7f63360934b0f", x"7e7d4e27aaa8c3d1", x"a488349a172f1da6", x"dfa166a9f3c62a23", x"9130069408d94c15");
            when 30761414 => data <= (x"c5ef11bb3b7ed1f9", x"d6554e2b074b805d", x"8f1227036890f738", x"00e349485b7c776b", x"1f63f94a5cb74b4d", x"814000dd51af58c1", x"960b8333462644cd", x"22645243a7db0114");
            when 12195806 => data <= (x"d47e13951b77f1d0", x"4a43c4ae5aacd509", x"2d6b8b800f878003", x"6dd691ad097729e4", x"4868628f3b19da98", x"acf5e56b4f3a46c2", x"e009e6e53bb52ce3", x"448bb3623a05da6f");
            when 31741288 => data <= (x"a48641d28d60f3cc", x"e6c7ff4fcfe07c4e", x"6aa3c74f5deeec7f", x"cd11025fa6493c1c", x"bf224045c9c0ae63", x"66526bb293333784", x"5d6fa69492e9db37", x"41dcd93b25a4efaf");
            when 13660795 => data <= (x"1fd6d676fa6a2fd0", x"edc67fe2d3f3ed58", x"582d1d918acfcf3e", x"7b78d6288af52a22", x"47d39646c3796484", x"f86fbe71c2f00678", x"bcf099103154d840", x"cb59408d82824087");
            when 27629105 => data <= (x"cbdc26c4c876733c", x"227c76a6977385dc", x"52189c23b9c589a7", x"7253148e7ab9b01c", x"c63786924e76b72f", x"2332a83b75d975db", x"4c9e92649212f17f", x"342d11747586ef78");
            when 25955062 => data <= (x"55b4b478d3be043a", x"e0d8686ec463864f", x"615c20cd94c37304", x"7df620fffb4a4073", x"349555eb261eb426", x"d08fd96cffe043e7", x"afa41e27a059e68c", x"a91d7f139ce8d309");
            when 6885595 => data <= (x"fb717e92a011bf42", x"66059e6c03b5837e", x"128edd60f44706f9", x"712ae3230c269596", x"b5e65fb4cc937897", x"60b81e8393b0c7e4", x"e0874db002571b5c", x"4cd9459034c2e64e");
            when 24624149 => data <= (x"a9fa5e299f2eefd1", x"cc8db61f0d8d96f6", x"06fb73a3f77f630d", x"eeac361a8c6f9fb3", x"c16c351eb0de689e", x"fc31433439516b01", x"1f0980ec14223528", x"8dedfd3f52b6a4c7");
            when 25454185 => data <= (x"4d860a4c09a6a536", x"b727cdcd909746b8", x"e65f47a1e4d48089", x"ae68c973056ff51e", x"1411d5bfdc53cda8", x"87fb6e8ba29845c2", x"bcb075ef84374fe4", x"0ca7f3281348ad7a");
            when 33747567 => data <= (x"5a3452272172a955", x"a651d4d9c4782ac2", x"ca0985c9b3eeb64a", x"496f2308e7cad6b7", x"52014514730118f4", x"b801929ff4485926", x"b8e9d8359ea473c4", x"5801745550b02f1d");
            when 2872797 => data <= (x"d37c6934b80df4b1", x"9af01adf94122561", x"429518c0892253be", x"4c22d07da5d79903", x"f805cb16a291d329", x"f219661acc1bf3c1", x"19bdff0c92a3cab8", x"946a3f61929b8b43");
            when 31815887 => data <= (x"78c8a5ca865ab044", x"65a70169ecf35498", x"0bbf2d44041ea1a5", x"2382729819a6f8bf", x"8381e27b6b64b489", x"a5684025269a4d8e", x"77eb43770836614c", x"f27d3899228ba22c");
            when 31561375 => data <= (x"46c6c20a10bffc7b", x"01600b96fe114129", x"f01bb06c09cbf463", x"0029264abdb84a47", x"3b725b0f2406db2e", x"408b3e31f91c7b35", x"b7051648880ef733", x"701dc2468ea0e585");
            when 15517377 => data <= (x"82bf4908faf59d11", x"51df7480c0aff395", x"fa220fa7aa2c8caf", x"ecca017287cebab3", x"97631d4ee9540a58", x"c11edf46c37460d4", x"23ce2ced114f805c", x"c5274911ade591dc");
            when 12728583 => data <= (x"69cb0bee73b84d95", x"0271b6afe89a3cd2", x"8d466cbc45e62e6c", x"2fec75f27b93d247", x"fce701f26324a369", x"e81ecf3bd76f611d", x"e4d2aab971253426", x"f0164190a0571825");
            when 12803139 => data <= (x"91a1147c96930829", x"e2931886b45846fe", x"675fbcb3a59deb9f", x"f1a98a6454ae16fb", x"12c8d2f39bf20bc7", x"221de9d7dfb71039", x"18d35242e09bac52", x"938fe512a2572c58");
            when 13566148 => data <= (x"70b62105b9f1b11d", x"a44c04998b233c31", x"f5fa7b6a8565f122", x"1e62dc4ffe91ecde", x"53782a81016f11b1", x"2b9856612747ad45", x"d7826514bd7dd630", x"b8de8f370d6bbf28");
            when 33859427 => data <= (x"747a14f31ecc3f66", x"f21fcc33181adda7", x"3604ee078622ff9c", x"7c71ac6e18c0b1ad", x"d155271a8165ed3f", x"ff45045c9d7db214", x"969140d0dd10077d", x"0a770777e74b4321");
            when 11662147 => data <= (x"881f9a46305aa753", x"91a7e1f13a5fb310", x"fcad07dcddf230d7", x"1592087b144e09a3", x"33396065460dd6a9", x"7b5f06ee637230cc", x"84f344236247b054", x"085695bb0c2d7a76");
            when 4105591 => data <= (x"494d2946366fd369", x"27dff94b52851721", x"62a05c5dc9227f2a", x"408bf7075afb019e", x"4cc9d61baa0e44d0", x"7757d82ee7c29deb", x"edd6659bf802ae2e", x"ef7f5ae7a815a4b7");
            when 14632142 => data <= (x"3627318cfc39bc01", x"94576a853f7dd453", x"94b547ba788355c3", x"b55e519987a57bd0", x"b7f67269a338a154", x"93cca9753c898ff2", x"f797d286a2572f50", x"d5911616dd2bced8");
            when 4160988 => data <= (x"b8c6a907796547b8", x"be4d45f0e0bd2e41", x"41731ac39e77211e", x"ac5f786675f7cd96", x"9f16924db6b0f409", x"4e485c3a48610893", x"7ffdab041a83f222", x"4d59e5a8ca3f4e9c");
            when 14084468 => data <= (x"2aba039defb96250", x"65ab908c5cb60de3", x"583bffc35f5fd92a", x"d7009e9d3fa981bc", x"25be96d1defd9e33", x"b7e615f23e470445", x"5bb8c8f78645ce4e", x"75766c86ea47eb2e");
            when 31912464 => data <= (x"d7e4073a678d6526", x"f6820efa8eb10b07", x"8decda292700b4f6", x"5edbcb6ea97ef593", x"a6c2c45f2926bad4", x"1f28c1cc4fc6b994", x"af73a2493d1cc980", x"34d5d4daf5838f70");
            when 16091801 => data <= (x"a8990c30ae87dece", x"10e279284fd92fc2", x"bc12e979d8d1ee78", x"e1cdc16151f6cacd", x"57e30d21eb0468f0", x"b65bc3e977d99502", x"7c1dbeebae573f4e", x"b8a7cec0e3d1614d");
            when 11080851 => data <= (x"f16a0dcc282392d0", x"accb785d309dbbf4", x"818e4c100dab4622", x"adbf0534e58ab198", x"c9ba926658d60a97", x"1476c0d5d3df1a6a", x"c2c9dd9abdaaa7ef", x"c2a1ff8cd065b9fe");
            when 16065431 => data <= (x"05481d88f3bdd5df", x"74535537e65af3e1", x"85c9cb47e54247cc", x"4190ba896015a58e", x"a3d7a64b854098af", x"3709b0eb3d9a859f", x"1c2cdda176923b21", x"6ee26fac30a3f599");
            when 1179270 => data <= (x"9b0154f83a12524f", x"c133f8f799f1977f", x"efe6acf90114f60a", x"646f112f4b7d7ff5", x"cdfe00e8c59965d4", x"f9e9f6d0f2b5e382", x"813a154d709399bc", x"9610d4f33f6fd0b3");
            when 15068265 => data <= (x"44bba904c498828d", x"b19c9e466c423ad3", x"3032dc744283daee", x"197aab3e1b209fbd", x"ff5fc8532ace6ce1", x"50473436b136eec2", x"58cac19dd520d570", x"1689b0862fb1b4d3");
            when 31313350 => data <= (x"5f4c0087fcacbea6", x"9841359803fb33c7", x"edc6123043432a41", x"e699b12375772a3e", x"885a59cf9bf2d2e9", x"50781aa042fe41a4", x"f1d027b16e6b677c", x"1ef2350303827aa7");
            when 12801161 => data <= (x"416a56f450b39563", x"61f7aa7c5f1ddc24", x"564e478955b802e2", x"a64a75101a4adde3", x"ef3a571712a350d1", x"ef19386eda8bf169", x"cc92b9782e6cdcf6", x"138cbf2fa9e555b4");
            when 25487551 => data <= (x"d91da2738f21b799", x"e2101e3433020937", x"c977096c6f4dc02d", x"e68cc993b55c1765", x"f81d75d8e270ae7b", x"383c299f6be6dc9a", x"37596b9569022159", x"ee2e9ec3edf3f4e0");
            when 28476695 => data <= (x"0bc5b71e569452c4", x"4eac7901e237e30b", x"e750b84740f945e2", x"8653e02168535d7f", x"2847efba1f7f229c", x"85e0ed2228f3ff36", x"d146f7087be8d801", x"4e3db645463f6fbe");
            when 32298271 => data <= (x"a6d6122e2233d0d3", x"0a9d31f61754899c", x"9209a0cbb62b279e", x"08c2553ececee108", x"69ea39909cf9af88", x"0fcc10122b47b141", x"eec76df1be6f8499", x"a1fe2a1aca69f7bc");
            when 3911887 => data <= (x"02c46abfab9be66a", x"ffb6b9fd0b4a57c6", x"b26a2a2d08a00701", x"3aa0e0b7fff87c00", x"ba93e262e26a2882", x"ec88e58eefbb045b", x"1d16d89e249ae1ed", x"f15b70f8df83965e");
            when 31619330 => data <= (x"23b4b1b958393332", x"8d235a72fbf407c4", x"2579548221a5472a", x"1bdc337484ea6c98", x"502bde2b45d50253", x"9e783220ee737f42", x"a40ca739317bcdae", x"7fe26e30bbe4b05e");
            when 29964605 => data <= (x"e45ca0f391ef42da", x"658a18409469ff19", x"10d287ec315abb2e", x"8ded7cddef3b4437", x"8434ddf8b6031a3f", x"5c139bd67e934463", x"4babb225cee6ea77", x"2050078fcdcd2ce2");
            when 3354244 => data <= (x"ce3b8a43b7593285", x"e81f4097bf52051f", x"80bbe5036d02fc3e", x"3b27228db0cd6793", x"d854205031cdcab2", x"237a6a7965a0033a", x"5431bb170a1f139d", x"4d55ac073b8aef31");
            when 32271129 => data <= (x"9a52bf0ccf175e90", x"558c3ccef8f2b50b", x"20ddece7b611ea79", x"4292c69bc80fa6a2", x"3f62f350b7a407dd", x"5d4bf477e9e1fcf8", x"5148711c151f1251", x"a078b0cab55c916f");
            when 3295826 => data <= (x"52cbe82ebb1c87f0", x"d09b0e7a8cf5b6bb", x"777a20a0cd6304e7", x"dcfadc772c08c7e8", x"8a36d180f755b99e", x"03d4ecc432998340", x"6aab692b00674505", x"542ef005ec618cc4");
            when 3787550 => data <= (x"0a24466958440671", x"b9348818a86c065b", x"8cdc8b21772641b9", x"a5e3a0541b568892", x"360823028d723bbd", x"9faff8c98e21e8aa", x"d3174f86e10d3571", x"22a3e54cbb35b8c3");
            when 21788674 => data <= (x"1a0287b89412e572", x"2959cff54b86c770", x"c98dd79875eab3ee", x"f491fdc541b2be2f", x"a37443bd0283c344", x"b02a3d1f8954935a", x"0aee4f0bbccbb8fd", x"8a874a3e971df81f");
            when 15208951 => data <= (x"4d3c69a53fd729af", x"e5bb4233a8bbb656", x"4dcfde0698d2f74f", x"5edd3989c111c407", x"9735a031612fd011", x"cd7bf16c4bce9139", x"4a8ad72def95ee8c", x"2e1e13b09bc0ebd3");
            when 6719055 => data <= (x"8923ef66d4157f30", x"2be1e33df7118123", x"ab955b57c595f94c", x"0db68069d9c345e8", x"dca0e33434dd0f54", x"20a9aa7081701d35", x"9dcbefd575fa440f", x"d44dc9a0b9f85ad8");
            when 24174422 => data <= (x"0eb240d30d5b55e1", x"ebfa877bb2dd9e4f", x"2446b05ebf08c133", x"36fec3d158a4d63a", x"502bcb67f5d4d1ff", x"2a57490d305e3820", x"c5dd33f51cfaacb4", x"61b6fa2837e2a90c");
            when 17889007 => data <= (x"67affb0e55d46bb6", x"bc3f6487709b1204", x"c27da8fb46c8ebb0", x"ebd8b52a738822b2", x"e4c36272b0964cc0", x"51568fe26d70d85b", x"2d8526ee2aa25c6a", x"2543bf96d3e092b8");
            when 12044983 => data <= (x"7f661e3756178a56", x"4a28e19eb89e4d8b", x"20ffebf9270f4552", x"6a1c2c268bc9dbac", x"73ecdf1d1d33a46a", x"965647a2e0481299", x"8fdcbd3141ca76e9", x"0037dfb821c5bcd4");
            when 11428975 => data <= (x"4d0b496cad2fcacb", x"bdbdded2c43245ce", x"03d8b47cd9e60356", x"15366a524b64bbc2", x"5c4eaba0c04aafa6", x"5ea2e42b8cad7fc8", x"05fe867bb8853c58", x"6c5d4c61c4ab4c06");
            when 24503280 => data <= (x"d5fecaaa19d9dfde", x"a9803791a9e5cd6e", x"1f998ca5bf4224ad", x"cb648f6d982ea34c", x"7a1ae2bdacdccae9", x"df466020780e00f5", x"59cb2957249d3e9e", x"c44db866f4671a7e");
            when 32284142 => data <= (x"de38272cca1a07f6", x"c537dbee812e7d5f", x"4be11ad7331084b6", x"5f40878bbd5d807e", x"9d7f5cf7cb423a69", x"65427175ee61cd3c", x"abfd58402663714d", x"d2198a7709d54fe4");
            when 3752726 => data <= (x"31eecf5827ae3caf", x"169bd509944b200b", x"0ee3196141d9e97f", x"d6b76b9f5f51f99b", x"3cbd2e7f8c73b322", x"aa6eac246f467a7f", x"4d5db1c400be6da1", x"307a85b92fb0a4e3");
            when 29550405 => data <= (x"29aeced1315d7ca0", x"7e4cd32a778a235b", x"1058fc873646f4c2", x"66ea25630ee1c06b", x"8845c0c34995ab3e", x"12db73f96104d4e7", x"18bed66cc74d677e", x"f420f2479f4ddd3d");
            when 23823240 => data <= (x"1b46bdc2a2227fc6", x"b47cda222adc4c4a", x"d70752d67fa5448e", x"311f799039eb1068", x"e9606fd32336dd71", x"eeb46a65a939a576", x"64a9d05601b2df95", x"785bd9961d3065c2");
            when 18410739 => data <= (x"597543ff3fb5ed69", x"1fc4d901088ffffe", x"7fe50877b24cfbbe", x"1933d639bac5ded9", x"ba62874ebbbaf97f", x"c5e1afa90639838b", x"c7f09a76d9e8dbe0", x"3145a45b3b436659");
            when 31406174 => data <= (x"af00149189b4f0a8", x"5cb1c49bcde4e452", x"5ccc672687159875", x"87d31ae02033e302", x"a4124d578abb2d55", x"829b73141fefe392", x"e4723a5016d630a8", x"1269146fb679f46c");
            when 24239836 => data <= (x"48bf5b7f927870b1", x"1e55085de8fbdc6d", x"733e1172ddcda61c", x"97d2e70597020c9c", x"acc4976471c75474", x"3f0fa57dc74be719", x"30b4a885920ca0d5", x"424712be891f87ba");
            when 12948765 => data <= (x"c4d7bc98f1a3a86f", x"826625f0f18ae320", x"055fb57b46e84bbc", x"bfd51e7fb676b733", x"f99bbd211fde5da2", x"4f75d5f3ef4df23e", x"3573f7b4f2b48e6c", x"22956d72aaa7faec");
            when 31956129 => data <= (x"03bbfa6cfb09e1e0", x"60334569093cf29b", x"e53de13c60fae1a0", x"6f2aaf7e7d6e4614", x"1e09552f9ced25c3", x"28346e00802673de", x"5dcdadc67f1b35a9", x"9ead9ee670c7d901");
            when 17329779 => data <= (x"065f94d904a4cbdd", x"72953aab93c5e0ba", x"80ced607d9506f82", x"d589e8fd9212fef0", x"ad702d415d5a7127", x"b1ceffa63b15eadc", x"411dd275a88012f0", x"7cb6f65e977fe526");
            when 15846774 => data <= (x"4d75a0f6bffabb3b", x"956bd480e0265218", x"72708ea28637b0bc", x"399d57754bfb662d", x"5df84482c392e287", x"3380c5e047de9c0d", x"a1efa7336e788d5b", x"8f8710a63bc11ea7");
            when 7237744 => data <= (x"0a3bc8d4a7bb7152", x"c4572572754d04d9", x"7abc381f7392e811", x"31f87ce70d4ae05b", x"07c646ca1e60f43a", x"6cbf7019fb9a77f4", x"47a90e915ff55336", x"fe53c2ccb2285e94");
            when 19460670 => data <= (x"5511d68dae5c2652", x"918f2dc2a9eff20b", x"556c35a0a44cc2cc", x"30cd5200ffdd588a", x"9853f1b98de24dfd", x"3f34be1d4ef72fed", x"5f95aac832aa3662", x"f2e2cae4979e5c52");
            when 21438161 => data <= (x"e70a904a8f0663fe", x"b9d25c261a641ac7", x"a6ce03def2e9e10a", x"7442668488eb23ab", x"adddebe8eb790fb5", x"1c6914d3749d13db", x"e4fed21f121ccdf0", x"8c873e661f0f94f1");
            when 11194397 => data <= (x"2a9b13c8327a8cbd", x"578781beabcb801b", x"e9f13fff95de2c24", x"7aa24872f54e3314", x"1d3f62a7c9dd11d6", x"2bfc78f0dfd44535", x"b3b3629f0c735b6d", x"347bd326801fea54");
            when 24998285 => data <= (x"87a9c842a67a41d2", x"6a61411154762141", x"58839973bb0ce4ea", x"1e67d32821508312", x"b14255eb4ab534f0", x"da86accd5b44680e", x"ce85b8a63b468c1f", x"8fd4e262bce7357f");
            when 4125328 => data <= (x"b3e08a06e26cd11d", x"199af18fc8bef9f9", x"5142a16e7cf05cfb", x"31943b8e9a336059", x"6484cd3f398d1a94", x"16306e133f1cd231", x"838d13bec001f802", x"0716fbbacbd0ef9a");
            when 16521601 => data <= (x"6d2280819cf5e025", x"2b4b4a395b9c41ab", x"b445ac08cbef7825", x"cf62d3bcb963de6c", x"a247299312d415c8", x"658837a2fafd2def", x"d2e27eeabb8e91d3", x"372784e93ec42472");
            when 19221037 => data <= (x"9f76d0e936161c8f", x"223a03f19481a366", x"a2a136bf3414ed1a", x"201c92eb2f13c6ad", x"efbab1131ae9f319", x"3154612611df8cf0", x"df962dcd3abf8937", x"e62d9b6a5ade2a04");
            when 29862856 => data <= (x"cd918c84cdb25351", x"6a0b5da9465e8058", x"5510eec718dec7f3", x"3ec10da8fde7718c", x"fd5070105f0a2a7c", x"73ce749bac272caf", x"4508422b9323b69f", x"2720dd12eb83daf9");
            when 1680266 => data <= (x"40369dd0cd912fc4", x"cd3bb8d63fa1b192", x"2ad8d48842c15820", x"f98b27dc525d3374", x"8c58e8675503fb63", x"f04417f1b96d9919", x"29eb307f51a495fb", x"8f20bdbca9673c31");
            when 14435042 => data <= (x"22152fb6803aef4c", x"949582ddd52a07cc", x"84ef0a2bd5c6eede", x"3a2589a475ec1c3f", x"32f12e9a29b9f9a1", x"5a96a0b904e95090", x"a70aa341f57337f8", x"035db1d0ca205efc");
            when 17174877 => data <= (x"0439321d3c15fac8", x"ffae6553ee479077", x"606f0798e9bc0d72", x"0337a1ed1f5a94fe", x"9bd0c5973188667c", x"408d237907f2c9af", x"21a4b0491447ba57", x"1ce9858576a12274");
            when 31344765 => data <= (x"e11a44cbbfce9a59", x"e04d07511d2fb33b", x"0e80529803840121", x"e4be32e4b3f0051f", x"4ecdb2632e1efd4f", x"397561ab7c192445", x"53b163eb77f07c35", x"f5b8342a85c640bd");
            when 16975901 => data <= (x"fe2f31e3ecb341de", x"200ead73148f41f8", x"fa0f182d4b0b7d5d", x"87b1d79d7ad1830a", x"a2e0ed98b436a0f4", x"9da1fd33c3ad7a8c", x"420c2adf9689e459", x"d14b80e514619036");
            when 28751717 => data <= (x"8d292d2f1766a746", x"132b958ff57efefd", x"dda26d9264de30a4", x"e5d62f051f37ed83", x"573334cde3eb2faa", x"594293744bee227d", x"38e444d2aa0c22aa", x"28cea14c1f4dd2f7");
            when 20596276 => data <= (x"9695f6796642784f", x"48db440d30b84f67", x"012fe713fdb63c53", x"8ea395e8ac2dfead", x"8e2314cf3fb244f4", x"f4309afae21d4784", x"45f9ab0544cc4539", x"307922deed3cd7b0");
            when 4172520 => data <= (x"5db6b6e935367ecb", x"0cb9e3fb4f27218d", x"6176ce5e45dff3d6", x"a149a289143c6b3a", x"15ee0c09008bbf0f", x"a97e591533261892", x"d4ad33bad0f01221", x"2d1d86db402b25c5");
            when 17623961 => data <= (x"3dc5d6a5866d59ce", x"9302fc76a1e9d051", x"095fe3dd92a5ccea", x"d91ba193c3de7b43", x"b513eb04c051c7c0", x"f8082e371b6dab84", x"f26e08768f6e358a", x"c06bae18dd35e52c");
            when 26486945 => data <= (x"733317dbeae3737f", x"21c4006fab127d95", x"7e4ab64bb9a67176", x"fdcbd3db13997b60", x"10f1b29ac976fac2", x"16a81ef5fdc08476", x"e0fa980d8b6bd3b3", x"c101c0a21a1d4e50");
            when 27698486 => data <= (x"86a1fcdc50012e21", x"85662f675df23766", x"260eebc35c449109", x"86df550f6c64c5e3", x"cd20215d2e8fc136", x"8c3beed9660cd75b", x"4146b537405fb7ad", x"cd5e16b033bf1e0e");
            when 22437539 => data <= (x"baebeaf5bd42bf48", x"c178215448a9ac1d", x"146892c02444524c", x"dd5c3ebb43f412dd", x"258be24d39f6c833", x"affc65622af6344c", x"e3be64c2666af827", x"2ae66eea7a815acc");
            when 25837728 => data <= (x"acb8736bef078c75", x"ede3510eb3877b2e", x"6ce27b6cec6075d8", x"4185e473fa5386f3", x"b2c55e670eedd340", x"96364890b405cfb6", x"98fd3a69ef6d9a71", x"bd5a71d90f4f2ffa");
            when 31009651 => data <= (x"b55556bb38fd3c00", x"5d9cc2cdf557590c", x"ecfa8062206126a9", x"d47855d035d594d3", x"e99bc5f91e7838d8", x"483a09991b1f8d33", x"efd6ca676c2c07ba", x"4e07346756512dfc");
            when 23897163 => data <= (x"37a1de71fa4655ac", x"7d769716fc2fe599", x"0882398ae2a9e93f", x"3ba913a727e14d3a", x"52be379fd66d148e", x"1f7f814bb37902eb", x"b4d0d279cc3d41fd", x"d0530b75708f962d");
            when 28509684 => data <= (x"8456bffe7327e549", x"55139e232dd11478", x"487ada318210e15f", x"0c553cedead74612", x"4280430eb2542806", x"283cbfa25183843e", x"82c24defa3b276e6", x"f8b51c11c334fbb8");
            when 18581442 => data <= (x"7f10ad46e0876c61", x"5cb9690a2778d934", x"0143ce72f6286a66", x"7df608c765cb23e5", x"079b4e76a7f404b6", x"252e46bc6ee53e5f", x"eb2dd2991b282a91", x"79746aeea23141f9");
            when 407609 => data <= (x"0f689e2e62f2e698", x"23ec208b47ee35aa", x"02d1f994b71e0079", x"7a1c2d03e6b77450", x"8e953cd593f37fd3", x"025ff424d393c644", x"31f3004f8d7e84f8", x"4ec0283d9b99e175");
            when 12967849 => data <= (x"2001578bf2ef7119", x"e43e6acd58c0f268", x"9ba759cb061f4a35", x"da02bb193d1e0b1b", x"3c7958a677dec1ff", x"6c37d30a53788db7", x"8043bccc53a68039", x"954b04688eb2fe8a");
            when 4729745 => data <= (x"194b35f0315b10d3", x"d73b653e84d09f43", x"cd575cb1dfbf3208", x"84a2ff1d07fd0e0d", x"f75f823d513f6e5a", x"e3e3bae202748a14", x"e430a560ab77ed63", x"3ff427f6ecc05860");
            when 12997213 => data <= (x"ac7579c269761d2a", x"f0fe9a8134ad06b9", x"12d51e49a622d9c6", x"0d76c2d668309708", x"e9d64310e112b2f9", x"98a63d91559f2b59", x"824f748e6739f94d", x"d1c9e6e55b3c6d11");
            when 31698531 => data <= (x"76950cc3d4f4d644", x"a63e81d070358564", x"0f8790cc26ecc1c2", x"2e6b8b137221df41", x"f429a4af8253bf2b", x"c73d80ad6eefc96a", x"cb9fca2a9282efad", x"742fcfeea666d8a5");
            when 26613977 => data <= (x"1f108a414dce5959", x"bde1f345290754e4", x"9164dfeb1b68f461", x"904bf3f0f9158f07", x"54d9119c301ce080", x"495b439e63f7956d", x"1e57eb27d7356187", x"8b73bab267f29b5d");
            when 32528885 => data <= (x"ec2cac0ac006cb1e", x"6367c19ed7660b4c", x"4ea189df99b24c75", x"dbc938879bb70d2d", x"22891dc373f7a745", x"96c5018f9d34c39b", x"3309bd9846b4008e", x"1641570d6895c983");
            when 21752754 => data <= (x"785ba1b9e0be9b35", x"a2ecc40ad5914da9", x"37bcf3869d007d50", x"989dbb69a76ce9f2", x"c2795cad2aebed61", x"d99e2f5aca0bf99c", x"72fb1368ca10f4e5", x"6ede6cd269e1dd9c");
            when 21265305 => data <= (x"2b73b106720628c2", x"61b32f3add2073e8", x"f684834b84093566", x"e2953371f5b25f4c", x"e9afb984dc16f16e", x"49ad108b1c9254aa", x"0ecfaa1f85fc8739", x"fad4003f40b66fb6");
            when 18539768 => data <= (x"180b66011e80e59c", x"da409a7606e866df", x"993fc0a3d9380219", x"fa98c6af1d530c49", x"a84d1840373d8377", x"157aeb5b4eae0c64", x"a2e39b8cffb2d641", x"297bf2ddf97b747d");
            when 22970020 => data <= (x"33db0db0e0fc45f7", x"662d70a78998fe2b", x"ebafa360e880f7b1", x"b247d963a83474b2", x"1968bfc10236ba4a", x"f249727ae441972c", x"ba9793803351b703", x"0737cfa0b6cfbc9a");
            when 13341603 => data <= (x"3daa8d159da31b3d", x"27ee77a724b5cdfa", x"4093f884e5137405", x"53a69f3bb8096978", x"95b59b4053446434", x"a3a96436b6ffe361", x"b1a62f2a5e171339", x"f4406fe66c9ac51f");
            when 3341614 => data <= (x"72d2ce43f6684b87", x"31468f29968daa0d", x"96178256d12f8fc3", x"1498d7b58b06a450", x"40173334e75421c4", x"bd540d0c2162ed12", x"273a37a4bc34b1d6", x"86238aaab8b9a7c4");
            when 15356774 => data <= (x"aabe21eeac2862f4", x"13d316faa67e1997", x"8094dc6115de1d10", x"414ad517b0843ce2", x"3a63ae597871f905", x"3580ada74626b32f", x"16fb1c87b368147a", x"25bc999e8fe5283f");
            when 10143216 => data <= (x"c5b9c4444a2f97d2", x"38241b4cff5eeb2e", x"c8a04b321f72aa47", x"c5c20a32b26e67c7", x"0c7683feee8c2c2c", x"b83e5da91e3ede82", x"9ba405ac04bff3fc", x"7d4081db5b1cc2a0");
            when 13458140 => data <= (x"aa29d3af0cc7677a", x"67708623cfbcde78", x"8dfc02b845fb8c2a", x"0ac4744b88c42ce2", x"37d455cb838dda6c", x"3412e0d1b3f7d54d", x"a501ac6ce40c6ca7", x"2fc2b30406e50407");
            when 5923678 => data <= (x"ee71019fe6b50838", x"c71faa18f7df5416", x"0f859a14781b7060", x"57237e55b94e6710", x"b87b43411e90a0b1", x"c2d89b9209dd9109", x"5967f1e3163b0ea0", x"db28f5d30c6054eb");
            when 9563446 => data <= (x"c9b94d866b8a14c4", x"e8152210fa2d2d62", x"a325563cfbf4df09", x"3bae04ac7996fb2c", x"d01572261412e439", x"bedab869cc398973", x"7f89e061da57825e", x"aeaff8d9dbd72755");
            when 11253423 => data <= (x"f757102a9b0d0484", x"3cd699d6774c55fd", x"cd7fedfd6b17eaa1", x"24690b2f7441759f", x"dcb1fc272c32e897", x"57c1dd0ceac012a4", x"cf8eea42a13d79dd", x"7b9881e572d37aeb");
            when 20696761 => data <= (x"6e72c68c57f85c40", x"824914780fa267cb", x"000af4c32ebcd284", x"7a685efb1b2dbb12", x"b739b32ca6c1fcb9", x"aefb182a304f3be7", x"a16cace7b2d30e23", x"a7e21d3a47029f81");
            when 31996591 => data <= (x"f021116aee9b134b", x"9615aaf92c865729", x"c6d8e0043519451e", x"54f0066224ba70d7", x"7455d0906e96e4cf", x"db9f0490af4264fd", x"af4ee9758fe9b39a", x"7bc8c4d10f7e13c7");
            when 17989326 => data <= (x"551e0bade0b2d2af", x"8b35c0bf2c5c17d0", x"db4e813d69cafc69", x"ab8df3fb4bc4babc", x"8f66f5db6e6687ed", x"2aa80a8345a1eefe", x"2f49213ca0b10447", x"d350add77ea656f6");
            when 5299102 => data <= (x"c680ef65041130ac", x"b3a423cf4576877d", x"ee3923d386396886", x"c57ea9e91b8b8343", x"821a1c2bc20d57bf", x"92b0d8669a7015a6", x"70ce4f529848ed0d", x"9f4cdf1678a4a273");
            when 29414829 => data <= (x"f2f8f9cca1355709", x"29da982a2f60acf9", x"860795dd00d56327", x"660039351c3666c9", x"a02cc9008c559e82", x"4f17df64330ca9dc", x"b82c321b629575ba", x"88e18ca7ffa121c9");
            when 9099218 => data <= (x"3fea61727a8f20b5", x"f3bbb161b7c63bfe", x"7d63d6263418c202", x"fc472d66625f1e1e", x"ad7fbc1ea25989d7", x"340fb5de622729e0", x"92cce40161ce29bf", x"671fc4bafd836e46");
            when 8061468 => data <= (x"d1f3ea0110bd337f", x"f1aa2bf494f6e1ee", x"0a90e427153ddedd", x"72eb84727c41a14e", x"b2d36bc91823604d", x"61063e585a309f28", x"95fb634859aad1bf", x"8c9fc3e4e3db37de");
            when 30820021 => data <= (x"3a73ff1e6391a1b6", x"23be7a30111c769c", x"241e595ed1b290cf", x"bcffd178d10efa06", x"44c9837bb7c70e8a", x"53647e31811f530b", x"b7f3d1c82f8336e4", x"3a6de87170d0c592");
            when 33107324 => data <= (x"95520a3244c0df40", x"6b1e2d51c04f24af", x"3bf2ef1dd47a57ca", x"15ddc40b8b093185", x"6f3407f2a45a6412", x"8c022c8671835503", x"0cd7bd47c48fae51", x"e593952c9ee8b60b");
            when 9716929 => data <= (x"7b91cf79cbe8ffe4", x"d1360de786183d42", x"47be3484b2796c04", x"f18300e5991a3d44", x"24d549b625de37f3", x"33b2a148f9b54a43", x"ada0b70229d370e0", x"58327a71decf63fd");
            when 21291180 => data <= (x"4afae97517390d01", x"f5a322051ef02339", x"74f58fe0559ff5c3", x"8e45e0c62ec2cc45", x"6db59b67ecdff247", x"1362b29e7c4b9388", x"c7c936e8ecdb78c7", x"34de064a07baceb8");
            when 9726800 => data <= (x"6dfabbd72b244f00", x"a2f6c64b6323654e", x"d8e1255f8fd8ede8", x"496e9af5f014414a", x"c986dd83174b910f", x"c4921321fbfe1375", x"3e828690705d9bde", x"61c5e1f565c75580");
            when 23713036 => data <= (x"a3f6d4920a5aa39a", x"0e52d918a041aedc", x"39b896fb6833b681", x"223e3d2a6c71b558", x"674dc65e4ebd6e7f", x"76c6944d22309d8a", x"c552b96fa742656e", x"b7e9c04602497fc8");
            when 21616220 => data <= (x"2908fb329b1e50a1", x"8b0997d3139b5b18", x"5f8fd18f044e4c04", x"80530b112b04acdf", x"1afdc228a5a9f660", x"a0bb7ea640c08bd2", x"5e8ff32fdb292c71", x"f4f2c70ed896caec");
            when 24561371 => data <= (x"9907771833983b51", x"7ef397fa667da139", x"b1ddc0f859380462", x"f462bb429e9e3db7", x"14078a574093b069", x"93f85d8c4019a2ac", x"00d6d3e62eb5b1a9", x"7271eca431ba4c36");
            when 24832064 => data <= (x"24223fd3f8cfd111", x"7c98ad769e9ad957", x"9579cd8fbd1d34b0", x"e5870e9dbf4396be", x"abb6c1922a64305e", x"567abe0bbc8d1f0a", x"b1376bb6ebaeb323", x"c85f3d83deb1684f");
            when 24481586 => data <= (x"1eb1d4567dd2d62d", x"f3f26e48cc3edc94", x"77c263d283581317", x"c8d920c2b1f91676", x"99bb6e5e28e8f74a", x"cb2f5bc7fc6a2c57", x"128e2e2680c32cec", x"fcf1d6e8e744ce0f");
            when 16890697 => data <= (x"09266d3e648f990e", x"428a677d92b4a94d", x"58cd90c92f275502", x"c598e702374e0dd2", x"4a54764aa450a760", x"f3a8c2319db130e2", x"e9fbd7bb19e27986", x"320476228ad949f6");
            when 18689760 => data <= (x"073400d5f8deb713", x"d4b2cbb9031d1190", x"fb3c2e761744c501", x"2dcf58e4d92b673d", x"afe09777dae6cc75", x"43460d9a240feea9", x"4f1911c8b42e67ad", x"38d8527a8ba45914");
            when 26184024 => data <= (x"812a00c5e34e908e", x"4573bf99798d3d97", x"ac1fca0cfdd08e4c", x"4c486f4896c467d4", x"54240cd1586bb683", x"7b0174bb6e2397d4", x"e9b35bff19f68ddf", x"2d1dcf435d06c668");
            when 15439899 => data <= (x"90c91cbc7d827756", x"5f431f21967c944c", x"abf3ad8c79976255", x"c33d8f98d0486dcf", x"a120a49acd824ac4", x"437d48c1eaa4ace2", x"d3a62f88549b7828", x"3e0f6c60782a1ba7");
            when 4939926 => data <= (x"28d3f03315915b92", x"437b0b3559c4da03", x"116f16f282dcb3f9", x"0f8c0e6f33646a39", x"30819661b188c2ea", x"d3556b5ce5f6467e", x"37ad5f3a328916f3", x"055a39564770b4b4");
            when 11409327 => data <= (x"c22e0a0cf09fd756", x"ff96208ddf8d492f", x"7ac58070f6500c2f", x"7e10cb794cea3fcf", x"547b2bbe3e8b98dc", x"7143efff6b7b278a", x"0ae27b1424c8e95b", x"45e2bc245715db29");
            when 29394202 => data <= (x"0199af5c7a5cfdc6", x"989d8bfecfcb93c0", x"cc27af9c2076047f", x"62e0dc0a5c036807", x"e95bb67803128a1a", x"d2fbfffa394d958f", x"285034e6704d9a1b", x"570f125f1a1caf93");
            when 21895400 => data <= (x"9a6584a46cea14fa", x"ecad5389f9fb935c", x"7d567a700c8e25e7", x"dc4af9cd48ed62db", x"808c507ed887de22", x"66f746aebe73b7e8", x"faefc12981043fad", x"640d08cef9ae0341");
            when 5310181 => data <= (x"3581dfd09ae22572", x"491c7266377d8c57", x"b106d4b0b3a526a5", x"35209258dbe37d0b", x"bee4c36577737fe8", x"4e74363396486b7b", x"9e60ffdf05bce759", x"20c7b0d9484e5d90");
            when 16869328 => data <= (x"e5d13785d4193e9e", x"287bcf0a9dda4ef8", x"f586210139abb49c", x"abd03c3dd6223edd", x"a3bb51bc59ec67d7", x"776bb547a9020309", x"4f119e7150c92600", x"99474894f6c61ac4");
            when 29444593 => data <= (x"bc7303c8b6b10585", x"3ff9f8124b52ef2c", x"57dbf62c216bc327", x"ea3dc31e940a170c", x"890da5a3f779fe11", x"bce0cf76630cc0dc", x"9de38b7ee9b6586e", x"4e33d0543afbc392");
            when 29960082 => data <= (x"f30f0b34c6f261be", x"4e9e04e3df7b8f9b", x"9f9898217bb6eb1a", x"d7e40d0ff0c703b1", x"812352b72fba06ed", x"210a4efa407c87de", x"1afc5066f50dfea7", x"1eae37ab30caefe9");
            when 21817427 => data <= (x"e3e83d4ab3b51763", x"423935d258066ee3", x"434af1dc0693ea64", x"bfa0294d86912e73", x"f6fa53480fc960fe", x"6a57bc5a2e5791c3", x"0a65c6526d4f0096", x"b4394ad670c9ec1e");
            when 4951030 => data <= (x"3a14e16a3b5693eb", x"37cdb6c8543ac91d", x"1abe665295c591fb", x"1c49ac18a553dcb9", x"f9c6d99533831334", x"0e08aa856059ab70", x"2ceb92eda9020d8d", x"9f6fbe4cfefe700b");
            when 11960532 => data <= (x"19e6b14acbaa6c61", x"f6a22b3b61c33bc5", x"cefd66141c4edc7c", x"ef7c66a44c2c7f3e", x"a5bd3624d8850572", x"6f4c318f847909db", x"54a84c0fea4ea63b", x"c5da7858ce129a40");
            when 25388155 => data <= (x"6359b79c506e95f8", x"19994e0b00d41b75", x"48ea9018e9ee32c9", x"917c5ec56f3eb6b9", x"d4d513ec2b497a83", x"a4ae80eed9c5ee77", x"21e36a341b9774a3", x"5e4dcfdf9651c27f");
            when 24729208 => data <= (x"31c45df762d8ff2a", x"de869d02c357f436", x"3b7ad43ef1734057", x"f5cd27fd346f4015", x"ca7c28bb90c9e39c", x"e1cc98a89213fcbf", x"a636b24410d1b8a4", x"aeaf4714332015f3");
            when 15312035 => data <= (x"b7e89c2a0be8254c", x"69a97dab8445f4dd", x"468a69f05d9aac39", x"53cd36402e814b52", x"299007c6541dbc11", x"98d8f542fdc2d5d2", x"0be6eca70efa18db", x"0fc0dec073c29d9f");
            when 26287513 => data <= (x"da03c0430f8c7402", x"ee16508813d877e8", x"0fdd0b6500eefada", x"9e3185eb1237f282", x"16ce78d28a4c094e", x"086bb4705da87851", x"dbfb26bab236069c", x"dc46b504de5f1ca1");
            when 27347179 => data <= (x"3a5414cc80b92c40", x"9704a3744088dfab", x"8a5d5f9726fd37ee", x"5c6f85157e5ae4ee", x"789782511b2a5cd6", x"4255caaccf4a5824", x"17df90f7d855296a", x"ed4f7faf9237c468");
            when 3628505 => data <= (x"5e63b96a120cd271", x"44b05d4043766cdf", x"0111b84d08f2cf13", x"ef49adcd3ab3ea1c", x"8e5f7d6e22420920", x"f44403cb09d6a599", x"8f6e3948c9cdbf30", x"094ce83f85aa7611");
            when 6886444 => data <= (x"d2cca66cdf0887dd", x"3eb5ebc7c3777044", x"8dca044f70442f99", x"318c8e1ceafe4bf6", x"a2c821790fd020b9", x"cee42dc61b51138f", x"e106e11a3e8b792a", x"3d72a88265dd1164");
            when 16267347 => data <= (x"ccc7ac427bce0e55", x"d18a6fe7a757f53a", x"c2f068f4b7ecc926", x"f0afe23323089edc", x"db9eb40a90c43430", x"30a7edd2a8bc144e", x"03f376e0d156c1ba", x"01739035cdde3a79");
            when 23096557 => data <= (x"398a420079a5cddf", x"a60451c1450fc768", x"0ce537cecb69ae00", x"782e2bb0a5abf267", x"e9c1f66e2ab74421", x"3b9455138efcc028", x"af67a3c1856c4776", x"0193e14a8db27674");
            when 29754214 => data <= (x"72e8f87950552e5e", x"75045246a9a23ec9", x"6d7f97337ded90bf", x"493ed0cd1a5f84f8", x"38e9b02e20142523", x"39db90e0df78bae1", x"450f51887690989e", x"8e53488ca84816ef");
            when 27608629 => data <= (x"1d5053916e369ed3", x"01381695bfc8ecb6", x"9327cc57f5f5e90b", x"3288785f7c025fc9", x"7c89779d76ab3b1d", x"ec7cc817051ca8b0", x"f08ae3ea2e09f058", x"a9db66c4a9d62b26");
            when 31997640 => data <= (x"3c70d865f678bd4e", x"5a748dddf9d10690", x"69bf6e2547cc65ac", x"9cea063bbfaed162", x"97a135767170368e", x"9ea462283cb3e779", x"3a96daf937ddf6cc", x"76fcc2fc46fd3237");
            when 32174918 => data <= (x"f62acfd087a48001", x"5634fefaa805cf1d", x"8de5673da6d3d27e", x"7ba819e26ec4b9b6", x"64cde7633fb5846e", x"5e7f593ac1054765", x"a136701831e885ec", x"cdb14f85d9a4ec64");
            when 17911106 => data <= (x"6846acb36b590036", x"c15462bf3839e5ad", x"69e2c2311e5c9ba3", x"0e534fe27ed3a9b6", x"b9ec03ddfad46c55", x"dbd8a458d379a58b", x"f36109ff58deb923", x"a4ae817240c256b5");
            when 1229157 => data <= (x"00cfccb506aafb18", x"62b7c19287d60b7c", x"d0a07b35f7f66407", x"ea8ef7bcbf8d9b5b", x"26b3d0d12c7b7db2", x"4922639a8d4c4028", x"cc90d5a39d9ffb68", x"12d5ec23a7359f66");
            when 29529106 => data <= (x"d6376bdd700d1af5", x"f705f5d0b7a83610", x"04087f2d1e2f9837", x"dd91d736958e9b18", x"a726e2c8e2ea8d25", x"327160d119641321", x"de8eb801080f8248", x"fc2ae5c04cad0018");
            when 22118490 => data <= (x"067da27505fb0079", x"48426d078127594a", x"23f047131ea8f9e5", x"e526cf33cc0ea17c", x"2091ce8ca435db35", x"65e70eedea892ed1", x"c98bb317cb7b5e25", x"200caa252ba414f3");
            when 10042289 => data <= (x"39f1650f5c1f25d6", x"8167f02aa1e3a88a", x"cd30ce1a0f4b367e", x"3f34faa00d2b0b26", x"05633d20a5343d5f", x"847b9955fa27f38b", x"700d8ef8bb454bb6", x"22d3ec302fe07c50");
            when 28837622 => data <= (x"64a8e8f9c259869a", x"d7ad33d588b9a96f", x"d803270e7f7b8523", x"479bc37d9c3c2c0f", x"12bb8633d6c1163f", x"46b9cba876a31eaf", x"6aefe37c7e24731d", x"21b77d27d6d0fbc2");
            when 21587204 => data <= (x"254db3201e723d3f", x"2ef3ca75f89f60fc", x"5dc25128d2928bec", x"644d810b8f6081dc", x"3c9f7f66bf45d932", x"cc41604cdf529b01", x"480d5aa3e9e525d2", x"e76db3abfa748152");
            when 14421853 => data <= (x"352f38aad695376b", x"4539cb9e5de1f813", x"9b9bb29490efa21c", x"d8fc7b5dbfcd8811", x"632ca74f63b4d2e2", x"90c6a83ba25db3f6", x"7f5d51c0bf99edbe", x"87bf853ef7495cff");
            when 24280168 => data <= (x"cf4732d62c770cb5", x"9a9fb82568813cf4", x"15b0e591098b6396", x"c5834fd5af86d35d", x"ad44ae67daec5032", x"2f65ff0da21123f9", x"95381ce498dad513", x"1d5318f0a3bf8a0d");
            when 7085632 => data <= (x"c2e13465992ff2b4", x"6a11f3cd9202fa6c", x"ae796ecc1cbaa72f", x"44cc58e9c62da3d4", x"b752955b79545e49", x"a83d1fc9ab8274b2", x"8f7b36a02acb6865", x"48777925f33fd71b");
            when 717563 => data <= (x"29ef977014d9372c", x"b4a5b608cc62f551", x"030183ca44f71288", x"d9c33177d6db078a", x"ef823ed7be2caabe", x"fa23efb1783693cf", x"879588514a4ed430", x"d1c1ef8bf330dfc2");
            when 32695796 => data <= (x"2168a2975820a5b8", x"e2273654d302a4cf", x"f20163387c6fac18", x"869ce1bcab412108", x"c45ee8164f229739", x"eb55333e4274e923", x"20f93e185b8b76b0", x"da432f73576aa13b");
            when 23757795 => data <= (x"aa81949ee216320d", x"ec0d3c9c3dfaff9f", x"62e96b1e1c272f32", x"c3fbee807e751247", x"fe5c179ac413b015", x"763e56f63089d945", x"c4fd4e51a9faed8c", x"040eebe18145abf6");
            when 33061844 => data <= (x"214fa2fb81dc76f2", x"ecbba77d89fd593c", x"5fac2e484a4ecbfd", x"ba19750744492c26", x"5af7ae6c492f71ad", x"68b2e604a4350d3e", x"fb2dadd92aceeef4", x"7d6fe59a3ad3b836");
            when 29421468 => data <= (x"7bee9298f09b6303", x"24928a20603f71aa", x"b6111ac0b406df9f", x"a1d52e9d45225670", x"555a69440b0315ef", x"41806facf32cf3a0", x"ec4218d083dd2c09", x"35967b66accde1b5");
            when 9419593 => data <= (x"2001e230e7498488", x"f89e0d9b934c82a6", x"6bc528977b6c73eb", x"d0db1f64663e10e4", x"25e2ea1ea6e08ef5", x"98e61d324c8af2d8", x"f7816134947f2300", x"74603458b13c72f5");
            when 22664435 => data <= (x"a7f1f1d8c28e1dbd", x"0ac5dff4a79fc1e6", x"c9ddaf0f55e77127", x"098fc8cc51bca05a", x"afa15f5aa2a8ab45", x"a165bb849d4e694a", x"d52e1c5210c57876", x"8a0dbd953490fba2");
            when 23980171 => data <= (x"042a405f46a56f99", x"a5d351c86991208b", x"d597604a4a4e4f52", x"11fbb32fb44d5a56", x"c4435dd8242c296b", x"7f18d5e7535549ec", x"7071fc3bdd90ab60", x"bb0ede0774598ea7");
            when 2483401 => data <= (x"f5bd0ffe5f5e803d", x"43b2c2d3c78e119e", x"52c6632f68f49c88", x"c0130a52ea6615dc", x"62ad4de9b1ff2b74", x"3e977ed16fe4a22f", x"f7c363271c942a14", x"2e59d5f8f587489e");
            when 33707604 => data <= (x"f48f00182ee7ed44", x"4ee8ea5b2d0859fa", x"b3ed4ce3de2d624b", x"37b6cb20a5ec4cfe", x"d3c6c8dfc502f19d", x"a5998c7b2e98c034", x"46cbed14f28f3cfd", x"00ef1db422212a89");
            when 2570036 => data <= (x"cb420e38c48a2827", x"065b1677fda6f043", x"00016bcb6cb7793e", x"e001978a2e6d985e", x"52a53f3f9e70be8b", x"5d44665a50f6d5dd", x"55e1472fd430337d", x"d8232ab4bd023bf0");
            when 9899935 => data <= (x"9e88e867470a4cc3", x"14b13d4fb883114b", x"64b593624716206d", x"6d3b03656c3e7504", x"06a5205fa7850cf0", x"a9825b86148e94f7", x"89186db8fcc3d95e", x"d6ae75219e042537");
            when 29144439 => data <= (x"9b5a557a2179ca98", x"6b4252bab23cfcdb", x"ad665975b824b68b", x"eb2545f17f7fccc0", x"2ef616f50eaccf1b", x"cbcf4897d243b103", x"1d94fb29f847af1b", x"c132e2eeecd38d40");
            when 33329211 => data <= (x"8e7f569c99699433", x"68d982a57ed71e4c", x"2bad79a1482243c9", x"6150b17aabe484ae", x"fd15027c920d2957", x"d988d8e574e367e8", x"a144a0ec6ba620d5", x"4250a70224459340");
            when 17195371 => data <= (x"c00f6916c66fbcb9", x"07cf93473ad94047", x"227f332ce97643f2", x"f43fee3095738ea7", x"8bb65dcd472ec6fb", x"77cc89a5d4eb15e3", x"666cda3803bb800a", x"7d0e022f51768433");
            when 19075186 => data <= (x"83ddc9d4a42e5c43", x"529059956e9e2906", x"fec46379a6e4d8a6", x"2fa3d5053d3245f1", x"4424b225d897caeb", x"23c66ac5fb078fd7", x"84cda611094260c1", x"30acf7efd4790aae");
            when 519639 => data <= (x"f6ca76cd259255f9", x"3b372a007880efca", x"4b0078c643f598c2", x"1a8619db94462484", x"4219bcc2a7f57333", x"984e445002f2602a", x"bc22a221ffd62ec8", x"32487bef4fe68099");
            when 31299260 => data <= (x"41f399de4eba3886", x"3398b60abdbe809d", x"1d56ccff8a38b92a", x"58169e9c09fa63a2", x"eeeaba54999dce12", x"c9ca55d9c8a29467", x"8fa74d252cab04b5", x"2bff3775f85dfa72");
            when 22876413 => data <= (x"80ac4dc9421d861a", x"c42ae9a0b3f604ce", x"d99b259020a09a4a", x"7243cb8c5470da94", x"eefb7af7d08c2965", x"b20fb01003f37a82", x"d6c632b3edc91ba7", x"703ed74db48fbc81");
            when 10941728 => data <= (x"fb4077d4f9bdcffe", x"217e901d3b6eb259", x"f6026b1714631195", x"dd04308e542cdb2d", x"de3e193de676386b", x"124420be1b5f44e7", x"2268030a111081f8", x"051c312a3ae09d82");
            when 2312866 => data <= (x"2e95aadfc11df26a", x"c7828ce5946f4ea3", x"c32ef11484b71474", x"4a57d67f426b040d", x"f56b8853f623110b", x"aef6110999f75d86", x"c6b2c0190e030f98", x"8eac83643806e4d3");
            when 20655277 => data <= (x"a4d415777c2a83d3", x"d8b356f2eca65ee8", x"0da2388419430cd6", x"ae25fd8250ea6211", x"ab27e03548d7d0d4", x"a63a1e36673d0777", x"1375522ac2175de8", x"5d6411cef9ab6d54");
            when 14448994 => data <= (x"325bf7aad22a6d3a", x"618a3beedfafb038", x"037e8041a413176c", x"09031a788469e338", x"5afd1ff0f8f4b7ba", x"f28604bd40c09dda", x"5efb5bd934ad5e6d", x"212a6946183af76c");
            when 30608377 => data <= (x"625e2ae55d2eb7db", x"9852a90ab1a59c5a", x"2f295d66a53bc7aa", x"f550cd6dcf8fc712", x"1d5934d06bbfeff3", x"3a30dbdca5b6670f", x"bab1e6a1ca925918", x"a2b312736d68a0da");
            when 17527421 => data <= (x"c82bffa23c84fa53", x"de0de6c66d428c2b", x"12e0c325160d76bd", x"94ab1e7a62228a4f", x"8780ae0b60d9d8b9", x"7e14992523350307", x"116eab37b93936c3", x"d8b3e44e3e1dd3e9");
            when 19925040 => data <= (x"71af762d0358353c", x"c3e53a10295eb663", x"77707030d8ffd83a", x"fdae6c93926505c9", x"e5734102376fef6f", x"7db2f52e248b0c30", x"d75513ef01ad0341", x"5dbd82cd5c7d127f");
            when 20146673 => data <= (x"d95f1c2c888b3eaf", x"3cbb3c3ef627b9a3", x"1dea590733731860", x"2d66bb1885943dbf", x"cd20ac9fe9111d8b", x"2d998930a4ebbddf", x"428b1a550a33d6d4", x"32383c9d407c6bde");
            when 18196647 => data <= (x"27f9a1d1e041917c", x"1e4a322a85b3703a", x"7bc3e07d51e30bf1", x"ed6abe830a5d4936", x"3fa8b8a7ac73dc82", x"629adfed73960926", x"78a66719b0384e2a", x"eacf5f5b212955dc");
            when 32166519 => data <= (x"53adef354bb045e9", x"3e03ef8d70320500", x"bf9fafc624d912c9", x"b8f4063c502cbf27", x"ea62fde7c634c6b4", x"a1564b1d3e58da4c", x"310dc1e5dd0d0808", x"aac0b543525c9cdd");
            when 15504270 => data <= (x"c1ebbd9b9cce15e2", x"db8624aec48a1822", x"e67adc0c0020e7cf", x"345fbdd6415642d9", x"16683f1fd65a7449", x"5f12680be472345f", x"cb146bf3f085d333", x"520981e83b592346");
            when 7888527 => data <= (x"3fe0f8e84289d380", x"fb6cb4dd5ec0893c", x"861731665efbd52f", x"2b6f289e075883d0", x"ba1ba0e1eb267ea9", x"2910f71048c4a138", x"df5fe0c3ee54bd67", x"06503ad8ba7aab19");
            when 32160550 => data <= (x"501f997a2921ffd2", x"3bb70a104b225785", x"f6122a44945066b8", x"462691cce32be93b", x"9a8e60690737b551", x"bf10d1ad70f79fce", x"dba9a232940f3421", x"07692bddd861857c");
            when 30603281 => data <= (x"e25ae7199d69c602", x"6ce6c9668b419f92", x"4c4b69faa9050139", x"3fe6dd823e1252fc", x"5a072d70857cfc92", x"9e532c2f7c5e1cac", x"292ea785bb96e6e0", x"f3955d0d35ca6f37");
            when 30902014 => data <= (x"a958302a1a79a907", x"e3709cc802131050", x"407cd508588b9fae", x"98c277afaa0b710e", x"d9f2195112f0b059", x"62ef85e5f0af5667", x"917a23837c78db9f", x"8cd9f358c336aa22");
            when 10140801 => data <= (x"427a9e62c29a9351", x"f9a119ee5e720993", x"ef6551b9b52b5bb5", x"d9ec767aceb2e8d0", x"d4457f52b439f57d", x"94eefa87f6dd7301", x"a1271754300b2442", x"3682ca51f5384d1c");
            when 22161632 => data <= (x"38e4c01d93e92a3c", x"025761aef26fb942", x"b56eb9aae7eddc58", x"83a4414946a095bf", x"f8aefb8c7ef9d33c", x"85097985eb67992a", x"d5eab691af5ddd3c", x"43a2763a7773d519");
            when 30627240 => data <= (x"643225c3b4e00ee9", x"d15d726d39964dea", x"6a9b086e2f3db720", x"8333f06bc8ef3260", x"916256bd23c39894", x"87ef81647f953a4d", x"b7060d1c6faf3ba9", x"cdb9f83a8ef53290");
            when 5328274 => data <= (x"26e418b8c4a90974", x"738a70aa0e1b6f72", x"012b6c9f731bd780", x"f3c2da2694c1092e", x"239b73259d3d8437", x"1a1fbb8665567e8b", x"a9107a7dd6a56a60", x"fc9eded8cef047c9");
            when 2893830 => data <= (x"f9aa649d73dfa95d", x"7abe54d106b11763", x"f6835e8c9b6cf510", x"eee6dd4a78eac855", x"1cdcb9b6f43c9c52", x"6af93763aac56885", x"aaac331f89a96b34", x"404bb033fbd10056");
            when 13047770 => data <= (x"ea31a7f96ffec100", x"e3a67cf50aaf2528", x"7f3caa8ca2f8b06a", x"87099c73451845ed", x"0be8f601e53c914f", x"9973540d8fbb1d84", x"92ee70accf85a3ef", x"4d86ce0c6d7ada8a");
            when 11964642 => data <= (x"0099404f2f3115d3", x"b30618c2b65547cb", x"97c67bb611b1ab9f", x"ffcbff894ab13ef4", x"4e7cf47356a1eaf8", x"98079ef95001edf4", x"1f6fdc8d0dbe6a2a", x"ed6456e5cd035c08");
            when 25547650 => data <= (x"677c8fab2552d10b", x"1562bdd60178f874", x"26f73ca1d7193d1e", x"ca0d91cd827c4427", x"3502212460378d6b", x"8f39f53bd35ff11b", x"6ec393268b8f4e14", x"6c97584f36fc70c8");
            when 15211303 => data <= (x"a3aa3cc90e4b2765", x"4242fb799d45d424", x"5d0119b62826b9a5", x"e302be139bd5588f", x"a498e7f785554af9", x"281dece8c8e7ac58", x"759c52e797380d2e", x"6a69dcf49ef6ae33");
            when 8037214 => data <= (x"ef45525d10b9ce68", x"c415a1cf3f955d31", x"a64b04bbb664fc0e", x"f198fc63d317120b", x"8fc7bfb0992f089f", x"b89e6bcb431909d3", x"3b438e3b57ffb025", x"5e7df4f3531db97c");
            when 29498433 => data <= (x"51ae08f2e933282e", x"b14b5a6e87e88598", x"3310c9b00cda2201", x"e318f40f500e7756", x"3647138cc2ab1793", x"fcbd32835aa978ef", x"310a54d7128e8906", x"8e80271f89521419");
            when 33426100 => data <= (x"50b96061c1241399", x"a4517ad66a37511e", x"3432eeeaf7bc4ffc", x"a52d44ccd66d1983", x"bbc48cc76d0932b2", x"e7602dd359ac3ad3", x"7029bc1137e4ec38", x"5c54c31bd2156ea3");
            when 29328716 => data <= (x"042fe698eac63a36", x"f1f3bc7d433885e9", x"d7c87b4dc4ae60d4", x"f081c453648e45a0", x"ec12cf2c77186a55", x"f3cd30702d723619", x"b69cb603e260b881", x"316b9a1574e8493b");
            when 32377179 => data <= (x"b27b64cf93085879", x"3e4404376a4f7f27", x"cd2fefe202546768", x"10fdcffae8cb6b56", x"ea3f94a96a0e0ec7", x"5c3245cf9e8e1909", x"9dda3735a6a26f81", x"082c1305a27fc457");
            when 27458088 => data <= (x"1dbd60396ebfcaf0", x"34c3f49d2eccbc68", x"63629ca3bd216500", x"f7bf722ab6b4bb83", x"592056d49682f3c1", x"cd6479e059543317", x"c8305b46bd1345b0", x"6e269a2ee79a7e6c");
            when 6732512 => data <= (x"02ec6d34eac4ad0f", x"6385ccdd183d0515", x"eceff9af77ca4bda", x"9aa1837d6f1b105a", x"a53a1eb491748337", x"29147fbe71c7b175", x"bbe8f6aea8f11a3b", x"12a7ad6cfd5bac0b");
            when 16803223 => data <= (x"e31767004c263a6d", x"d3386dcecd51d7d6", x"2ff714b089530120", x"cf77bcd68656dcb4", x"faa7ad9a99cfd66a", x"1d5aa6b70e9a078a", x"ae6b55d195274e2d", x"75d088ba6c4615b5");
            when 22110926 => data <= (x"46e3bd73f1738ec8", x"7cf2f05f562123c6", x"897c6a98e7335a59", x"c86812ecc26fed1d", x"a6f65f833c25d318", x"7cc5aaabcb3a524d", x"432358358d4a7549", x"ac5fb267382319ad");
            when 3635590 => data <= (x"c092095d1591e67a", x"b5bb9011662a6a61", x"a2ca9859f949eb3c", x"0c2286c8bde12fe2", x"510d16c9b8bffd77", x"bf2ab32314be5ce0", x"25a8323645b63fff", x"85463ddd57940f72");
            when 16148773 => data <= (x"6b96b3e5766d2255", x"1eb50acc2d23edb3", x"8284725e972533e1", x"aebb13eb4343683b", x"d0cf3b5a01df0d66", x"511ca42a4cc32425", x"1a1f50530ddaf4f0", x"dfa06f89cead75c5");
            when 31648315 => data <= (x"29d7ee148d83061d", x"3259811d370ff741", x"9abf30eb2607d454", x"03a69309fd98fdb4", x"2d5d05e41f36909c", x"f7f3f0f269ac2372", x"b5713198cad0466b", x"69e297b46b6fb38e");
            when 27613709 => data <= (x"31dc6597518c8ac5", x"f78e6a62f508c435", x"6c095914586dead1", x"43be891e3903131b", x"8e5a839381c03a07", x"532e29b6207a9aa8", x"4c3270f5bd1ef439", x"8b277d74de35482b");
            when 15200820 => data <= (x"b3595ec88f288c1f", x"97a1432d959c653b", x"935e76084ce0b352", x"14e4468f16ddac88", x"e2ea237b2c8e06ff", x"4cda41260c738537", x"39c6a62f4f3d84ed", x"b24ee2923b4149a4");
            when 32296094 => data <= (x"b9b14813c1d1202c", x"bb9226a41625d100", x"487b7f468cb4095c", x"89c3fc7f4cfbdf10", x"fd853fc4cc41290e", x"f048a3ebfa2ee328", x"9d4cda6b50e63d0d", x"cb02783564175f14");
            when 20967992 => data <= (x"e14008b62255a39f", x"9d7990d08bbe95a0", x"7d52250285ebba6f", x"80841ba496d843d5", x"d1ae7d78f06dbd09", x"f0b98308a0e05318", x"6b6ed02df7663850", x"e5ddf8c92439ed01");
            when 3813164 => data <= (x"092ffcb730cf4ee3", x"b09eb8212286ecd1", x"aed9a61b1ba6cd05", x"a668463b9dc6b6fd", x"11595b1e13b9edf9", x"289a7747543f8f9a", x"24d6f63cc1c8d4fd", x"2cc133afd04d96fa");
            when 19097589 => data <= (x"c4a67740cfb4f2f9", x"3aaac87c86ae8f79", x"b936f9fbb7fbcbb9", x"bc8ab8eb0d24dd00", x"de9f519d72e7991a", x"08b737c1148ec13b", x"73379461ea308144", x"742b655e2c6a1ae8");
            when 2450870 => data <= (x"35d403c015e26c12", x"a57a5d6b95ac8fd6", x"ae2cbcec22f5aa35", x"78c830a87c5b6039", x"937a069a6585dc46", x"c5fbec236c098e97", x"9e6c826e2db52daf", x"9dbf2bf187c4cc76");
            when 13661565 => data <= (x"cbb41681ac67c6ca", x"eb59bc89cecb0f52", x"983057a9130fdf89", x"d9d0a4cc0d4506c5", x"ad77ee61150cefa1", x"f4d267cbb8eb3b14", x"f901042bc667c276", x"d06a42289a264c6f");
            when 8018559 => data <= (x"6f904d0a04041951", x"64f9e8eae59a7eba", x"c8f42f1fe4e39694", x"b67bf0ccf61366cc", x"4123f23ea08341ee", x"0e24dd303027850e", x"e75bd6ce164e5c2b", x"6d2c25e1428a1b92");
            when 32739964 => data <= (x"df2a8e0b6c688f9e", x"9f2318aa1016e59d", x"931777c9b9097648", x"76d54748e9298f13", x"bbd924ea19da2661", x"36ce1a0bf0a9a789", x"6fb761392d8a84e8", x"a3cefd4bd5590519");
            when 29128242 => data <= (x"f37c213b98e7b726", x"5f8a37940a3155b7", x"0185a2c95ab9b807", x"d49feeea10fa36c9", x"9cabb255e5973b04", x"cd31aa8be74f6147", x"5eed0e473cbab68c", x"27c42e932effc13c");
            when 23291443 => data <= (x"fa970f75a222696e", x"8cd35b5519ec1a39", x"473ae1115913379c", x"f98cc34e91d69778", x"967e094088da01fd", x"7d0cc6ecdd9c4424", x"bb5974d55bdac457", x"7b3d46ebdcf58e09");
            when 26696886 => data <= (x"d46dbbd43aaa0d3f", x"2591dbdda9eafa59", x"06d4bb48597ded9d", x"a35877c0f7644deb", x"859fc97cbb5c8b5b", x"e3094fde6d43b237", x"76c71ec737bd3ae1", x"e705779130a983b3");
            when 33473241 => data <= (x"aef2718fe7d7064f", x"01926a75c9233235", x"6d2946eafa49580c", x"5c7a3248b453256d", x"7075c725e9e4416d", x"1d708814dd1ff599", x"9f84b27137be2ea1", x"34801761e6a7b9cd");
            when 21605763 => data <= (x"f36bf0d0ee8b96a3", x"043fb7d550bee62f", x"d336b1e24d6ef798", x"c09f63bb4d1ffd35", x"aedd0a84115b6f8f", x"d6e23d85c061aea6", x"044bb0e358d4d78c", x"ba93de6ec27fcd33");
            when 10064942 => data <= (x"60c54aff7c7da255", x"8c862bfac04c425a", x"06bdfd394f100c98", x"8c4dc544f5697648", x"5b35d286a739be3f", x"fe5277d30afad859", x"b2bb7acfdfd804cc", x"9b4cf4dfb31a77e7");
            when 27881675 => data <= (x"2cce6e54ae151873", x"4026108cf6cf67ec", x"06de33befc0ac683", x"36dd7152521c0f31", x"16812afbce6fe407", x"04e0bbc46d22a01c", x"5f08bda01b72bec9", x"6006dec55770217e");
            when 24456372 => data <= (x"862d3bd079a1b46d", x"cdb3aec28b04c0da", x"0bea29cc1d86b552", x"84b9d8f609f5f16e", x"aa1db7d318807ce8", x"bdc8c3cec14b3545", x"ac0be94fa5073aea", x"3a8855795356ce63");
            when 2534972 => data <= (x"9258443a92eae7af", x"1f033ed2ff3a7229", x"5218e7e912401d9f", x"f5691f642b4db42e", x"00ccc777c83b2257", x"3969bfdd1da0611c", x"892bc78fd10d1707", x"6ddd7bf607c8bf94");
            when 28773501 => data <= (x"5a38baf004a45e74", x"feaf6b93f02abb97", x"3e91d28f4689852e", x"b74fc7a661a8ba91", x"9bcdaf3a808ad98f", x"725862e6347c9b73", x"ca0132bd3ba41979", x"54e47cacca68576b");
            when 5763009 => data <= (x"610021a986effe7b", x"2df764a68391631e", x"25d1f1efa50a428e", x"3bc882211f7d723f", x"75d46a096f421eca", x"6f8b941c14f5a626", x"0559fd521cbf5719", x"059d630d24cbb212");
            when 18682330 => data <= (x"5283dbf57752b932", x"6ff15b12f7debea0", x"3a813004cc8aa587", x"4cdb7eca48e9cb89", x"fe1c375376378898", x"9fa484d8f9fabcd9", x"b7429a772b16fb34", x"ece69d68ae1ca465");
            when 14787388 => data <= (x"d1373dde42d9de7e", x"2985ed2a7e42b318", x"e90ef0dac48e7423", x"2defcbe62fdc8f94", x"9c58c3a80cd3345b", x"e563d5d025e24e0b", x"83167f141ef41f2d", x"43ae0fb0a43ed13f");
            when 10394075 => data <= (x"f92993845405d037", x"9517e5ff30c7fdc1", x"ce003e0d3f66745b", x"0494c35f51bc02e4", x"c5c048e7dff3cf0c", x"20147d56b7368dbe", x"aab078b7ee3a60f2", x"caf6b0b4fa7dd323");
            when 18899652 => data <= (x"fe59c50cc0465ce3", x"dd6a80cee561b593", x"bd96be3cd2685ac7", x"2db73aa8c839ecd1", x"304c82941b62f2f3", x"70a120a3a125e5a7", x"507b9ac2a7c7ba65", x"c1346129cdab1038");
            when 28746923 => data <= (x"2433d08ca4713813", x"7a60cdf055c4a56a", x"ea86e48c15b54808", x"4c5788924d1e8bc9", x"35e5a760756c104c", x"5697703fac890779", x"f935021c3a261cc3", x"df7a47b7f32cc202");
            when 18979132 => data <= (x"4d78528900185f7a", x"33274a9605d1231f", x"7998c70b57596a04", x"0be457e0be0a5ded", x"43b9a71b32c15b2a", x"bb5fcf736a6450b0", x"c2d930d9d966efab", x"c2b53fceb0727dd6");
            when 15868340 => data <= (x"7265f74215716451", x"2fb2ca5618dfa0af", x"37661c1df88c1127", x"1ed77890bd31284e", x"1fa1dd530925247b", x"9904d690d1b40d63", x"6f45ada9884ed5d7", x"b12f29c77dcabe3c");
            when 12981386 => data <= (x"0ae8aa3fcd917a2f", x"65c3c79c67266add", x"e2cc34280c105081", x"8765e09536f64101", x"8a20e825ef754066", x"035d73acd0e9f41b", x"c60a3b435ceda162", x"011f04204663065e");
            when 23385859 => data <= (x"1192a200bf8ab7cc", x"71abdc95739813fa", x"055896fc3d7424e4", x"68f1d8e4718a2e56", x"7947561d4bb12672", x"43640f0a33f8f30b", x"746c1d0017929cf4", x"9349aa196802b749");
            when 2454985 => data <= (x"7b316f39d84a0851", x"c5989a20956bd214", x"a97c9e8f03382843", x"0731779f0a49957d", x"ff0de249394a2a64", x"60fd0c77b93ff7c1", x"15db4ef21a58d27b", x"d9036d6ee151cc6c");
            when 10507231 => data <= (x"cce91ffade67958e", x"86b190d0f2bbe6d8", x"e22f0349761ef474", x"4cde137bba29aed3", x"574cc7548b886b7a", x"1c9812fe82f2796e", x"14e453e86fc66374", x"99531127766dc552");
            when 16758652 => data <= (x"e6560385f2038ea3", x"d05400485e88ef31", x"e5e3d801611bf751", x"7e96ef4323b70ba8", x"829af32d8fa0eb7f", x"66548b575d1e006e", x"fd0034432d3152e0", x"716b398e7dc1f16b");
            when 4796384 => data <= (x"2d2e7e8b4b759697", x"817c6c9dc0922ba1", x"dab6517724d295be", x"804dabbcb2fd3864", x"13434665e76d9849", x"7a28155286c7346b", x"904ccd8b8a9c0d85", x"1921b337fbc5364f");
            when 18507060 => data <= (x"6cb9390088dd2241", x"90fb54f7ebb344b6", x"b648391b5a44f48b", x"8e07cf04f9f733e2", x"de37c2b238083677", x"b1fbb1614444469d", x"44193ac8254935c8", x"d879225064698603");
            when 25333588 => data <= (x"f0ad01781060a328", x"96af004195a4a3a8", x"bd8fb890c0f42a93", x"1e1bd461cbda03fd", x"0b120a701aed99b1", x"e2ce696d077c252b", x"fe05796e06853e5e", x"681385f5555cf845");
            when 9122099 => data <= (x"5bffabb28d9249c2", x"c871a23def9a1208", x"65c4a7c6e8006a3f", x"12c2a5f134e1c693", x"13d4746e6f44c35a", x"45f0ee8077f99f6d", x"a13a480b756e6821", x"5398f7148692744b");
            when 20690486 => data <= (x"f884a8b9a4e9ddd2", x"d63488bb96d9b1f3", x"aa9592b16f846b96", x"78d24e49388f9b04", x"a8ca7637f7945ea3", x"cd2783a5fdf2b7f0", x"aa8e672773f521fb", x"282ddbe0fa645ebb");
            when 20454979 => data <= (x"73abe29574564895", x"89068a8ca95b156f", x"3163f86c27420ab4", x"96d49d64ac501916", x"f53fc095b2077dac", x"c36a40d37dd9d3df", x"c19540c5dbe80519", x"324a17b403567423");
            when 6929022 => data <= (x"591223160460ffb9", x"990d4f7b85409153", x"ac151fc8e97286c1", x"4297d910af783cba", x"2cad831a53b6f118", x"93be55625badaf6d", x"1e213127b5203849", x"12602d5efd235825");
            when 27703851 => data <= (x"eb71759068052642", x"0e22ce987168cdb9", x"de39fd953f395187", x"ca975cd538f754e7", x"04555e4c7f3b9726", x"39d9163250878be0", x"537e3cdb6feeea1a", x"6ff2a625e38ecd78");
            when 23752311 => data <= (x"c47d1ec38b451742", x"4fb469262aff54e4", x"57f8ce12f84296ab", x"2ea7a9bbb248e7b3", x"9a1c894f18ee1ff2", x"9f5876e295f55119", x"153ecbffbd971369", x"4c32e293d2cb6778");
            when 5146065 => data <= (x"53eb521e6d9da5f8", x"716ea102ff27a848", x"fae840fe560871f1", x"744ca01ce580dbbe", x"72e793edd73bb9c0", x"df2408e4cd466b67", x"f84de38149990512", x"ae4c779fdea61d18");
            when 12470161 => data <= (x"c90deef7177e7c3d", x"01d2c3ba34573f48", x"0f4155b77b55b374", x"e509b9f4a889e851", x"44fd254e48d73514", x"09a39460e6d3462f", x"05923be2992baa28", x"b6e6204151c85077");
            when 22017170 => data <= (x"15b7297bdaf661fb", x"8efb9b14cddb982e", x"7c524ac9de21ca01", x"b6f7941532a178b5", x"ff17a10c97ef2080", x"483892105cbe6d89", x"9fe6eb71a8b824d6", x"ba5eec6d485bfef5");
            when 12400056 => data <= (x"be79b980503be838", x"111fc83aea6ebb1f", x"e2a24f15efd1fb7b", x"777d557126476afe", x"fc85f865ffef06df", x"f22b803c0ed0f380", x"2439eaec4df1ed59", x"634e5eefad88e9ba");
            when 33269769 => data <= (x"a45f2662466bd54c", x"7884fa10463303a7", x"69a06bb6e47b5b85", x"8500de8911a8d78a", x"26a4a603a49d2bad", x"58ad861333204b78", x"fab44a545dbc2fd5", x"7683ede6701995c1");
            when 29439094 => data <= (x"a16ceb4bc48a76a1", x"0d7174592aef9996", x"b5ec0f305c7241f3", x"d941a27a2840d8c2", x"9c77257caa261302", x"7676775d8a21d867", x"b2fd897e7ecf17bd", x"f5c047f2f1f22944");
            when 11767448 => data <= (x"669f164ad0054904", x"a79c62758829a7b7", x"cf8ab9cbb02221f5", x"b0de437eba340093", x"fb4b7bbdbd4a297c", x"fa7e231fc64936a0", x"28d496051ae4678b", x"187bfbe280583221");
            when 20775558 => data <= (x"d8b733b8fa588006", x"1c72c66c58e84295", x"b3daaf187ae5d801", x"e95d073ac43ce183", x"a6634f0b7e064b2c", x"722b8f07ffaab250", x"82f6beef798395e5", x"58b4c9ed1a5178b8");
            when 1597259 => data <= (x"8e72e61b1e655e60", x"74b22015949f7965", x"5556cd9de5417a95", x"396909f51bb8a658", x"e6902423334c9f87", x"ac8c0573be628cd8", x"8d357d12e9c48703", x"9b1a2b6061dc8e16");
            when 2844587 => data <= (x"28ec9fad288828a7", x"19da23371239f961", x"0a9700718fd5f3cf", x"5fa74183793d44fc", x"4bbf8fb347e6fb72", x"06e35d89cdab7476", x"d350205662b87332", x"1e123b0b7a691f59");
            when 12171755 => data <= (x"0f288d9056326841", x"28dc62b54c5d1e67", x"2a259dd757de75be", x"8c5bd3d0c43f75b8", x"c020f65356e4c490", x"73415c761d508d50", x"c3ecd22a2ef59cd6", x"e3844880b4b2503c");
            when 24987934 => data <= (x"e815f0495b25c320", x"b18acf1117481a46", x"d8b60c324614a616", x"e278183daa47d383", x"7fec19027a3a7643", x"b047d8ea4edbd546", x"7df67b07625070f4", x"81de7f7ec32ab936");
            when 7733448 => data <= (x"8f30d988bbb95a2e", x"3e3946703c3c72a7", x"79e7d0e3e92f809a", x"b467794b149c1d82", x"ad37106138c712e7", x"5459573eb96052a7", x"da486d8bed9600f8", x"eeaf61f8333e1d2c");
            when 18600798 => data <= (x"eb1790f2293a22c3", x"588cd1e7861c0eb0", x"98a26099d55617fc", x"340cec1207f77194", x"0ea03dc0c4cc6b4f", x"191040f47a1c5756", x"0f115ebdb79734af", x"2f0da1a73ea955eb");
            when 29799651 => data <= (x"495f756adaf2bbb8", x"dabae0bc5b087727", x"ad431410c72095bd", x"a7d396917d108572", x"4ec906423c85ee6c", x"6885070191e66dd9", x"0f29d4f3cc50507f", x"6f6221806558056a");
            when 26198724 => data <= (x"064ea48a5bae8a44", x"3dd9ef8dcb1053cc", x"37a3593e04cde5a9", x"2fa2960dde219364", x"63fedb15b16f5dfe", x"26d882866fffe8e2", x"3e8943289b9bfe47", x"9a229b31e48e5f9a");
            when 14721524 => data <= (x"e1754d318c02fb02", x"e27515d69c69f373", x"d8a801dab81270cd", x"b52115421cc4912d", x"4b8b1bb1d52de855", x"2972056b27bc5ff3", x"45dfdcaeef264a65", x"6af49e7729dd13d7");
            when 8427316 => data <= (x"c89e139ec0e34ee6", x"572c9f2888eac768", x"22f71c3be2b8c6e3", x"e94fc8377ad59f52", x"789f2b246c2d9568", x"ef4dfd8632d03d3f", x"bc6f36bac33519de", x"6dfac488ce80145d");
            when 18899576 => data <= (x"4051fb3cf4e69ec9", x"8248e9a46c2fc8cd", x"d65798aa52f8a840", x"a9fed80fd93438d6", x"5c1accd06053980a", x"3388317407dcbf7a", x"1b7cb5e71fbfdbef", x"cdd2f2dc22cf0301");
            when 15276517 => data <= (x"5e4658ac53042392", x"c30de13246a7d245", x"91e828ff29c006ac", x"28ca088a4e6ee8eb", x"c3636eede82e5e27", x"67f818fa73e10ca6", x"129eff3c7668a991", x"c0b9205c7fe9a066");
            when 3512738 => data <= (x"5500826148478c6c", x"123718704ecc133f", x"b0f96ae01ef47ba3", x"8c01aa613906960b", x"75180368059e13d0", x"4b070ebd447479e0", x"014a0ab924e53a94", x"1aaf8c71bc1f87ff");
            when 19302503 => data <= (x"fb5a46300fca60b2", x"a49f9e77296e2483", x"8cd7d7b7c51002b2", x"5460752733f94c47", x"ab1b64c52ae3429a", x"f1a6434ac30b160b", x"8cf09d18175cc9e1", x"22facfd8ae6416a1");
            when 16721402 => data <= (x"62dce85aeddf52ba", x"87a66a92d9772f4b", x"87b6206de41f9597", x"ac5006c32873dbcc", x"1a9c8dcb20c30046", x"737540e3c7b0c0e0", x"e949981648877909", x"23a17015748dd984");
            when 10881638 => data <= (x"24a3d768984ad011", x"427474e83cd26121", x"3bd778f6ea12d2db", x"645960c6052577e4", x"9a2e7819d01f6438", x"5ecfa5a7f6563633", x"a068061a4e34d894", x"72afdfbd97aa50f4");
            when 12732330 => data <= (x"215e01c765adef65", x"1f5c2fa5e9283c64", x"5d678652e986bdbc", x"6732ae656b0c6a08", x"6048aeac3f341bd0", x"b11621fc287d6258", x"487a464289eb674e", x"a9bb76ef416f80d9");
            when 11633745 => data <= (x"a78f26865b4bc8f1", x"8b29306734558ef0", x"7908506519783524", x"49ef1e09e45388c9", x"7a98e9ae290e6d58", x"b2ee53e9f880083d", x"f3514cf71d045f44", x"11835f937b2eb99b");
            when 14473385 => data <= (x"381ea851ede4dcc5", x"9a23ae7744312253", x"eadef161067b0224", x"3938cbbd5bbd5822", x"e85948d00e3683f8", x"86f7c1f30c963ff4", x"dbaa094c67dde653", x"8d211047b29b0ef2");
            when 3353676 => data <= (x"b1b48bd47e1b5e46", x"d4a72cb6004d0ea1", x"d643ea4ed0f96afa", x"c8417280f593175b", x"07ee5eef3cb1f617", x"659b3ca193382360", x"6524ec1d63079829", x"2fe72ecf29e017c8");
            when 19661117 => data <= (x"f701e935158a482e", x"ccd9199684bd5768", x"59102c28028f19bf", x"f2ce690aa09fb89f", x"6c918923089fa582", x"e4fff1511b3ee151", x"39ac8a40b7f77de3", x"9c084a4c96199670");
            when 3145930 => data <= (x"b1eecc81af6e38ae", x"fce3cfbc3c402c38", x"bd854cbf4cbeeaf1", x"4d712a6b36f13838", x"22d50d842aeff283", x"df27cc392d608ac1", x"d438b226eb5d9334", x"5c8d399f2ec83598");
            when 32415998 => data <= (x"15f3d71d84bac2e1", x"acfa7ffa062523db", x"bcf998d0281f921f", x"5f051eef07c0acf2", x"3e4ddcd4ec5b8961", x"e624a14f0fd241c5", x"967180567ad43101", x"2b5b90a4ff7e0a7f");
            when 25586069 => data <= (x"31b4a00e3d21672a", x"f938d69b9ca82a90", x"46ca73df7cb82b9f", x"a77747ee3bdbd0b4", x"19d817b1220204f4", x"55d1cd604168c17b", x"8490de42a32412eb", x"e4f64c1b9ee0c5d8");
            when 22925393 => data <= (x"54ce9850b950a43e", x"0978fd8d6ef1f26f", x"54184923401388d1", x"7acb34dbfe61c008", x"d795c5927834d77e", x"5d29d45a7769ccac", x"5a471d6fa9570c3e", x"f572743356c65011");
            when 29501067 => data <= (x"866fabe416f8c33b", x"6a78fe93b3d9aa24", x"aa09b770b807f331", x"4821694900390eeb", x"72b2c9936186296e", x"f5380a5639c10580", x"e352fdc3eb67f57c", x"614037b1d3f5a41d");
            when 11242225 => data <= (x"12e787321243644e", x"6203032fd3956eda", x"9047e14256379cc8", x"2be621217df8cf65", x"7db286fb2cf9be48", x"d1762878f5184550", x"a54156eef97e6f5b", x"8107b5b69f1600c9");
            when 21666701 => data <= (x"ddcf8d84ada2b5ad", x"9af0fef795bbdb52", x"bbf8e83a075fdcc0", x"f6af8beb3acf7b13", x"e1e78babef9bc7e4", x"b047f1b91917ace8", x"3e5d8de87a3eba4b", x"eb48ca9453d2923c");
            when 3159974 => data <= (x"97a449f69c6d1717", x"32049313cf47531d", x"e2fd19b46e483343", x"1f5e662dedbd147b", x"b4adb831057ec365", x"45d564b8ea6bb147", x"527fdffd68095951", x"8633d46c830dc0f5");
            when 33633150 => data <= (x"26e060f3f3dd91e8", x"457aee38f9c16a2c", x"748b48f0872968c9", x"e66e369a217a3bd7", x"55c3d164cd8b0a8e", x"b31c3bdec773acae", x"f2f5c1bfa6e8fee8", x"8e89adf5fffad75a");
            when 29942303 => data <= (x"0efc36fbb2da1700", x"d09293d55b64a7a8", x"2596376f6d6481a3", x"f8a2223fbc62973c", x"ff239d61b9073b9d", x"c101f4e332a6a949", x"9a2646b6712cae57", x"6783c3a4ea1a0265");
            when 26375644 => data <= (x"fbf66ce622473f14", x"ae415e889625cf36", x"281462df2d8422d1", x"c2ff919f64f1c10b", x"73b3dca48241cd6e", x"f591192a859fed4d", x"5f76ef6299f3fdb0", x"09b815ee9eb488a8");
            when 32156485 => data <= (x"bade8d353a112713", x"13e064d9cab964ba", x"060a3dc9871083c4", x"b9174fd69cf74183", x"050d498fbe435927", x"b6726ae982ea1ef1", x"1221a0f537d83c40", x"ca7aecb7a4695e9c");
            when 18608235 => data <= (x"2372e9608635f2eb", x"2c30b5f29c5396f4", x"b92f9e47970cbdd7", x"3dcab5cd51e55c06", x"d6424e3fd465b1a4", x"7a16445e44626531", x"3e92d17b24cab221", x"beab020d587833e3");
            when 31203810 => data <= (x"423834bebc6c3652", x"0c1f577fb4332186", x"49fe9e54b43ef1ef", x"96a3c4c174d697fb", x"33390da8c204b99b", x"77f410d5dc5f749a", x"2b71a61c7447bde4", x"c4e698da39c145ae");
            when 18771781 => data <= (x"c4f54b6d11ed78a8", x"b51e42383217b463", x"777cdbbab47b9f93", x"c89ee056d4582918", x"b9b6095fd38f6839", x"a9e5fbb2827eff7c", x"d20e8a11e2700f90", x"8f8b34a5ada424c9");
            when 12489712 => data <= (x"ec1e02314d3960da", x"3eb19c2713496b46", x"e720cc9b04a0f145", x"966040d81c19fadb", x"a50d2dce995f3274", x"69c14e26d4288844", x"2909e9d42f4a18e8", x"ae6081a00b43dabd");
            when 3969945 => data <= (x"38c0eeb3d43caa0c", x"eee8684d0e588bfc", x"319312c2c85ca670", x"792b67d694e36b2c", x"596398c22fd70116", x"f94a9ab865f072a0", x"8657ab024251995e", x"e0a95fdd7c25802a");
            when 3738921 => data <= (x"088706e51ff631a5", x"fb850538133dbe2c", x"1f239c1593a092aa", x"4493555204ca84e7", x"ccebd1a1f3daff28", x"e9cc6339ebfa5d0c", x"846ee52fb797d45e", x"2406c12579fc7f38");
            when 29683207 => data <= (x"fecca611ce1b0606", x"44a78e6990d7899a", x"2df2f69ed1683a1c", x"e17d2199c81cc158", x"0e95d7e480364616", x"d769aa79e14dcd4c", x"94134d63f998ba7b", x"4c32e0522fa125e5");
            when 20596386 => data <= (x"e627c67f64714cf0", x"1acafa8956d6f023", x"fd3aaa555e772b6d", x"bd92b60b1cc3a1de", x"558947c286554777", x"ff91ce965bd0b0df", x"d439645c92eb63be", x"27c9cbf4cff28602");
            when 7999745 => data <= (x"c0acda29daab7a66", x"ecc557ca92ed74a3", x"336300710c0810c4", x"95b0121123b9306c", x"7ae9957cbd210f67", x"de202e6a7503bead", x"fffac2a29a37173d", x"35846a1ef6311d81");
            when 1468653 => data <= (x"24bf9089c5307e95", x"c76eb16d58387dc1", x"bf379e3775fd3a8f", x"b4fbdc25bcce7ec3", x"b6a0fbac96da8db8", x"375bd25dbaa510f5", x"4466d45d63e1fea4", x"bd5ced4cff9b4d26");
            when 30163183 => data <= (x"2525ad9d18e14f49", x"fe515f849dbe8240", x"333e9ccfa2855995", x"6badd4f28bd4f9fa", x"2e39fd4bf2c9fbfd", x"4aaf32518bdebe7e", x"24aeb4ff440a4d50", x"7db8737afbee7ca1");
            when 15659754 => data <= (x"7feb3e053507c190", x"add8ccbe74cc5e84", x"14bf514d8edcc460", x"e398e5738a7585f9", x"2a1fff85b231c24c", x"d01bb0ff09a1e02a", x"6239fe73c40c8956", x"ee4ab315d219d6d8");
            when 26279539 => data <= (x"c62af139e728db78", x"3fbbd2308b219401", x"92ec0b66f656b62f", x"ba3cc0e02d447320", x"266d2389ad31ccce", x"608684e35a5bc3bd", x"171905b5e4192dfb", x"3490e9ba4af93550");
            when 16154388 => data <= (x"4dc7faaf799b5051", x"82bb86b34b026e5e", x"44a2c1c16b25a57a", x"ae4d1575a60505df", x"1f9d212d2b904313", x"41f30b7f7e6e04fc", x"6b6881f4b800786f", x"449dbc9c4a6eacf9");
            when 17518759 => data <= (x"1248a2a2c92d19f4", x"1d470c6fcb186901", x"be59a6fe5d286b80", x"e7ada581cf4b5536", x"21407492c705ac56", x"06485d38fec5728a", x"18684a93eb06ce75", x"4f4aac162d9c9ca3");
            when 11115025 => data <= (x"1c38565e823eb5be", x"f9ffa1e117932dea", x"2709b03798a3214a", x"7f19de15767a9900", x"98d888ba70c49103", x"a3c98868d2026453", x"950d19616b765263", x"71b87a1fb0fff3db");
            when 30449358 => data <= (x"3e09230b13100c58", x"1da33e83798d0f8f", x"827f6516b01b4fa6", x"d42062d76a24586d", x"99ad1529fa3f572f", x"868cd0b8bb8eacad", x"e81c94dc0378506f", x"d76c6fe43c3cbae8");
            when 25807528 => data <= (x"892e17971ae21f7c", x"4d47dd880a2fb48f", x"ef46a2c583f25bbf", x"5d20d04a4a059fb1", x"f1fe479e0a03cd72", x"680d63ad56bc4870", x"100551dc0dd8b86d", x"9ca5ae9fbd085f7b");
            when 17495415 => data <= (x"c935ce4c44dbf44e", x"f644539cab12167d", x"bb7dba783e03778f", x"3a63c6d6e27a7b07", x"176b846451181659", x"dac39bf03640e2a3", x"2372d75dcba78aac", x"dd1ff4c481ad1fba");
            when 26587483 => data <= (x"f5e0b08c2adc371b", x"b08a90cc847d7323", x"b6cd61f23af2c54d", x"2e0e77ef55d99f5d", x"ec27543adad4e7da", x"7a0d33eb2510c2bb", x"cb5ed6a0d15480e7", x"94051914d305cd6e");
            when 23578879 => data <= (x"e29e91e6b7f85dbf", x"161fa44101086c89", x"9d8c4cfde056e261", x"f4e3d5edeea89636", x"ab651aad42179c8f", x"9df35944b9243ba0", x"0223dfc1c833dc1c", x"8b862aa10dc0447e");
            when 17923050 => data <= (x"a6165c944fdccd81", x"53f02e9b960127ef", x"0f1814b9c2b968d1", x"947ed974c6ae088f", x"55d7c6b76b83c016", x"8aeec67ddb76de12", x"f4d86005aa29f4c4", x"fe98450da58b7ac9");
            when 10257289 => data <= (x"fb4d4e9ae5927e8a", x"4b30560ed42e757c", x"51fbf9c2c21f249a", x"c39ec835ddb89375", x"e9aabc25c8e55ee6", x"516d5b21ec802b18", x"1dcc86580e91fa6b", x"822f0a0794f7a7e0");
            when 31448765 => data <= (x"1281855bfdc44e7e", x"8f752a5d1755dd19", x"00e5e36417cac2ae", x"d85b91f98ac26b37", x"8615e952468dfaa3", x"be53b2466035cdd1", x"42ee7a27cb323db4", x"c22a46ec02fc9f4b");
            when 11169364 => data <= (x"6d58cc72fd63ea02", x"bb0f95715ad025a6", x"570d1ee18008d19b", x"991f3f38e34cb1d5", x"f99fe8ddd808ad1f", x"c0779d9b5c2c278e", x"2247c3d9d7566c99", x"7ed2276488aaeb4c");
            when 20203978 => data <= (x"d1095a697f6ce5f9", x"fc72a5ff523e7bc6", x"b58ea5fb573e1f53", x"42cabdeb7fd17843", x"c5b17dd73341a9c3", x"e242d26c3720ab9e", x"f559c8d3822d3b0b", x"4ead2b34e62d7e08");
            when 4269662 => data <= (x"615b613a1dfc67d6", x"ef6c580705ffc902", x"ac11b7ad6da6214f", x"f99b1d296986beb9", x"b1344df9433bb7f8", x"8e6dc370657e40d5", x"6b0601e28afeb697", x"f67f52d6ebf8dd05");
            when 7995491 => data <= (x"184dbc43839a3e83", x"137e8f663597eef9", x"c237e81ca91867bf", x"89c24b72e67f0ffc", x"064dd37aac9a4ab3", x"cd676d441ed2d9e7", x"e290c28938f80552", x"3297195714389645");
            when 5747822 => data <= (x"9b3b1260fc442299", x"8aa00cc337ebd51c", x"dce38921e819d8f9", x"89857178544ad707", x"bcc9f566f0526c71", x"dd6357e29f562d2d", x"917aac7bb44ef4cb", x"b2fe8c4a6f059ebc");
            when 32363186 => data <= (x"16989d267f2581da", x"12b8c1f1b5779b5e", x"3777bbc109b43a0d", x"270f9d0db4b42122", x"cee7670feb513a29", x"7c828251c41b5fa2", x"95f4f1ad6ec155e9", x"2069bfab2540083b");
            when 4881939 => data <= (x"7e2396b150bc6eff", x"142537f7d71c1b7a", x"14d907be82c3c8b9", x"ffe0ee9f823f6ed2", x"42a0e12ae014af52", x"9ffaad23d74762c4", x"182a7683daafd004", x"7a75c494a5689819");
            when 29705205 => data <= (x"725598aa7d0e0214", x"53e8deb756de5f3e", x"1e458a09b872d830", x"847fa0790ce2c38e", x"5901793eb70060ef", x"56a2589fb2a530b3", x"e217c719906a1228", x"414b109bebec2f2a");
            when 6798267 => data <= (x"c464f712c470d00a", x"cf54228453def7fd", x"dc08e394d958c89e", x"7956065f4ad2086f", x"a1984ed76c707c89", x"c53fa9e39657d5c4", x"c39d25b0006fa3d1", x"d1378c7a5585880c");
            when 31014388 => data <= (x"674f65e2cd936bad", x"76aa96045b3cc8df", x"b1b42ee12909ca5e", x"39de3855d645693e", x"76a06fd82462eb48", x"4a344081686b355b", x"7c7d9ff2fc9270ec", x"b4ce262d37e80f7a");
            when 19390323 => data <= (x"49a6b62345e65eec", x"99eb442c4951c7d0", x"d9242628a57bd398", x"45cb1bda53b344a4", x"103a284e5507102b", x"18ffb0da75b30b04", x"f0f7593a463ad167", x"f65e0606fae04792");
            when 19307865 => data <= (x"18ba05b8706fc9cb", x"2be01c0b7f270eea", x"5f33b915c0e82dbd", x"6146fffbd251d47a", x"6a6bff74685dc7af", x"ec12faa10869309e", x"8a21890f01a9743b", x"6d37506ed60ce629");
            when 30533391 => data <= (x"b014aa64e8f9a64e", x"3eaa407528baabb3", x"db5a269439d84b6a", x"a5d2397ec743d304", x"f0fbf21dc79adb54", x"37977a4d256facf6", x"0391c31fcd42d9a9", x"22bc5fa4995989d5");
            when 25549937 => data <= (x"17f0c504b2b9a8fe", x"febfe845ade590e3", x"8b514d47485856d1", x"bcb19f43988cba91", x"6cd5a7c7d7a8f6c2", x"340a320c2e1bf6d1", x"b2bfc50f1eb71bce", x"e07fdbdca834ddf4");
            when 6543431 => data <= (x"01733d5ea4f5a61c", x"af0c8134f9c8f44d", x"861e1a926484e32c", x"2e9de8e2ced61591", x"95d2c996a7e93e97", x"eb75f04d3675b224", x"356050de555b0f92", x"976700b67decbd95");
            when 33524974 => data <= (x"5262b958f3fe1915", x"c906e0dc7fabce2e", x"e5ff43ae2c799d14", x"a099cd3757cfa049", x"645c6df1c899912b", x"0649ccfd19495be6", x"7c82d743a128d239", x"f84e48d983ad9d91");
            when 11068255 => data <= (x"f4a146c5daec196e", x"ef4a180c244d91d1", x"b918ab1e03ec5c9b", x"64d98416e42be4a2", x"0a628b99ba7692ac", x"8fc0efb6ab551c4c", x"cd14f759cc7788d9", x"cc15167f589d1419");
            when 26106089 => data <= (x"485f83d52d5c0b12", x"02203081342c4c4f", x"ddd9ff4326913596", x"6f1073a9d3824759", x"d1650ab2d582e222", x"fd3d94a3f8fe1e72", x"49cbab2d43a0bdb3", x"85e4e8cfeda96e15");
            when 4340311 => data <= (x"a3719c25d14066e4", x"b273b714a7a0ad76", x"2de770848fd6ab67", x"af0f6130ef0b8b7b", x"df0c3c547dd29a6a", x"cbf758cd5a8fdb4b", x"30ec3d4743aab38f", x"745fd86fb5582b8d");
            when 18974324 => data <= (x"d17817c72d8c5773", x"5669fe3296c3ed77", x"7b2357e20a004aac", x"53bf17a00f55b7c4", x"637b70f60313b125", x"ddf8d73c11800988", x"837e7ffe5954c1ab", x"25088c129a2489b8");
            when 19961112 => data <= (x"fb2465aaf31b3e37", x"86341d676df01bc1", x"f8cc33f3eb6786fc", x"bffcee309918f517", x"3fbf2855ad268792", x"eb2f3bf01c8a628c", x"3c328644bb4e982f", x"87887313b10bb73b");
            when 30472584 => data <= (x"b430146b67f6df63", x"a3d8a234e75df128", x"2a931c94236ba5db", x"45f8ef419df299fc", x"3ca617ea99c26285", x"6a4a3734ce9b19ca", x"e582ff9748efa8a7", x"70e7336cce03917e");
            when 16899714 => data <= (x"1ff9977057ef0f1b", x"962d9a20af9df88e", x"f5c4257968b6739b", x"7e5919e250c6bff7", x"89ff860a90a5241a", x"19817337fff79f60", x"e9c6d6edc0c2b59c", x"767f57e3c45b2a3d");
            when 3196421 => data <= (x"7c29ae143b6e2668", x"f4ba30fe1995591e", x"4ecb34a9d7edc4ee", x"c66a36986552f03f", x"dc0e125a2e050ccb", x"63911314738d4eb9", x"7fdb491099144792", x"bd432a179253cb0b");
            when 20772908 => data <= (x"a2e933c9b1a14dd9", x"0f2751155ed2f781", x"9a79a2103fd5070c", x"09d6d6c754473c0c", x"32c848ea858115d0", x"e4eae1f89157cf73", x"f6e32a8bb47efa96", x"7aa909b5397d2139");
            when 25494179 => data <= (x"b928c447ea1cb713", x"e0230ee3621b5bcf", x"badfacc303a398d7", x"851d914bb5590010", x"b31fc53d23a548ec", x"3e2a4c4959c2d1b1", x"aafbec2777839334", x"76428872357b9d6b");
            when 33299443 => data <= (x"c59aee8742cd47b8", x"ce5de0645ae3975d", x"ae157a66b1ebee1f", x"9d90b2b938e96d86", x"64a864fbfe9ec812", x"74be4e7c42385e48", x"b0ebec0a1fdfec46", x"0376010ef24677fd");
            when 4050154 => data <= (x"d63be90319d1895e", x"5b870d66e713e5fe", x"b2235fd58c04c4b1", x"a0df9e265778a0a9", x"4d467df32bd8370f", x"8e5fdf20e103b6cf", x"09b539b6d3e228b7", x"d4dc090af906ab2f");
            when 24568229 => data <= (x"49c2d4117afc6200", x"4ab7a22bd4775c83", x"06caf175447ae963", x"4a5303aa06d08149", x"529b41a54309b11c", x"937bd6c6f1c095c4", x"865f67b001565696", x"d5d193a8dcbc1b57");
            when 29702803 => data <= (x"01128e3b7fb2afd1", x"512b151e45b25eda", x"fff793399d6dc967", x"d233e682ba661247", x"94420aecc185a27a", x"8c9e3e0af3db2667", x"65c61dc1c8d4427d", x"284cbf3bb3b14a0f");
            when 554962 => data <= (x"f859bde4fc2a64b9", x"a93a39495aaabf6b", x"f8240e932c9edb33", x"685d259ed2b3ba73", x"1011dab6ba1bbbe6", x"a9a50ee48cd7d8d0", x"451d3c7d317f07aa", x"29227367a38aac4e");
            when 23455587 => data <= (x"fa970967417e491e", x"f93618c669d0efc2", x"40b699aab40a8d56", x"ba4057c4e5e587a4", x"f0b566c793cbac3d", x"6bf2ecb59970aec7", x"59eab809ed51d9a1", x"212c705ba27bae7d");
            when 31449953 => data <= (x"72689f7687327d6b", x"8512e68bd92b72f7", x"625a34bffb630736", x"37671d2c56f34821", x"1189b105f9b00a58", x"152dfa35d68727f0", x"5af52e03ea391fec", x"128bce502905a081");
            when 19630436 => data <= (x"f6db434f3f6ba9c9", x"09243f97531ad20f", x"040929da99534f13", x"161bcce69ceadc38", x"f046993c0eea5fc4", x"4958cee4691c5ea5", x"c1c9d59340a05760", x"005fedfe3aaa0a97");
            when 3827923 => data <= (x"b843a5d2fc14186d", x"07249c2827466f36", x"757bca8766dbf66e", x"a48e4e82d1b56d49", x"6844d77d94770dba", x"2ab97d113867723f", x"dcd13790248f823d", x"abef22913f076abd");
            when 28222242 => data <= (x"294655d36f8840d0", x"770676e943a438ff", x"a5e6d1ba97942779", x"27f7e1253a30588a", x"b71505390291847f", x"4b80ccd99ec4507a", x"473f62c454102347", x"20b3f94dd397694b");
            when 5998692 => data <= (x"05c3d07a606a5373", x"0fbe4c09614d8362", x"d180d940f87854d8", x"b2c0d0aa13da8712", x"69f2329573bbd86a", x"3755a6cfa6a9889b", x"bc57f7fdb99434c9", x"1653c19d183b0e70");
            when 27424279 => data <= (x"c6b95d230f8f9f71", x"ee81b08b89aeee96", x"224a9764c0acdd12", x"e10127ca3f5cc6d3", x"ef7748d07c15ca64", x"397e9748b98522b9", x"a9dd0fc3a1872386", x"6953052524266bc5");
            when 1772840 => data <= (x"dd413bee74b77689", x"a38bf39cd7bbbc00", x"e5cb5d2ce96a4c4f", x"8022b9923a44cd87", x"e9e32575a76ca404", x"c36a31d432aba787", x"7b027f8f17f7ca7c", x"4c3861203cb64a7f");
            when 21833795 => data <= (x"7e66d8005487e616", x"dc192184471c9591", x"54eaec33810946e2", x"afe67b6f308fb8e6", x"6b0e5582aeca97d4", x"38a7171c1f9496b2", x"9abc0a322307aace", x"95b3b8f421453b0a");
            when 33524167 => data <= (x"cec4a968ec6f6908", x"c272882e8d885b4a", x"5cb39ae22406dda9", x"6e314560e079b6fd", x"80431a86928bdf7d", x"a9fc0fa186ebe160", x"95b949f37c7612bb", x"e54e2e1943e54767");
            when 10874573 => data <= (x"245f2330cff71cfc", x"70116f219bf4ee74", x"e0df9eeab3779633", x"3f3077d8dca36f0f", x"f68977e7fafa38e4", x"0b381206f1d55d60", x"f3e5c10783141183", x"3d1694c95b960868");
            when 12905978 => data <= (x"b4cfe6ea2997fc7d", x"cce31c51de692772", x"bc2613cbd31d7796", x"a95ff4d23aa3369f", x"addea1ff5435f998", x"8a2bad2b1de15b86", x"e0cf26a44d6ed766", x"4a45eac0166ae995");
            when 10849783 => data <= (x"a434df876031f093", x"1cd04743fc6f3020", x"474aeaceafde733c", x"831309f4bf2eb012", x"3676a81fd566f996", x"a46e6de568e283f3", x"928ed8afba07e8f7", x"b3fd41f3841566d9");
            when 14397380 => data <= (x"8097b2afe285add8", x"b9b70fe79cd494ec", x"04f8a3d07c9f0565", x"59ff473140a76019", x"1db2953acd578f50", x"7755c71b51df17bf", x"bc4fa7e2593ebaeb", x"4b7454128137caf3");
            when 27464099 => data <= (x"a13a08bc6c30e935", x"b651d493ea548a69", x"ae3d77558b45de82", x"0e417e909e170a10", x"f6cdc36e6c736411", x"6e553707f37086d6", x"aa3fbfed275d3947", x"a16ea2e53cd75228");
            when 6912228 => data <= (x"0c1bcffeb46c9797", x"c89e0ab0610444b6", x"5831d7f2992c8b0c", x"e3a9cbed6ba894ae", x"1f0d26abe2e0a19d", x"9887070c832a5c51", x"6cbbfc282d5ac5c3", x"a1e94176f7223c07");
            when 33302071 => data <= (x"c798996827c84e59", x"e8d543f11f3e0ce8", x"6b40cd324fb94763", x"a85caa8848480520", x"034093d4b8f02522", x"4e3d2d47835aa413", x"1182b1296a595812", x"b4e0e88500c4af31");
            when 14217344 => data <= (x"cd4c231589357603", x"341c499f5405f0a1", x"3ce134ae10c9406d", x"76840100675d0f8e", x"e9a6053ec1cc5c74", x"763f3b9699daac1c", x"1fcd1bf98df1781f", x"dbaddaf1d86f8c87");
            when 32031751 => data <= (x"931a662c71b3949f", x"706f2b64efd0b1d8", x"dbed54df7c709900", x"bf09ce0f0dc7cab8", x"3393c8a5d4c5ac2a", x"70910aa0fc857be0", x"70b0a1d3a9ec89a9", x"886d7a1def79263d");
            when 23854971 => data <= (x"36fed332235ad8ca", x"2a5e8944c471937c", x"38e6d063a73d3af6", x"e98eedf058252b16", x"ccc7b6c9a471c18d", x"2f2bc2141942318c", x"e0b24f092fcc0830", x"f0d718c61ffa64c6");
            when 17106173 => data <= (x"a56e527b1a23a7f4", x"da4394873627ecf5", x"1a7437003b728784", x"8d6f7be23b623b05", x"de57c834f313d004", x"ca14bd959e7d8e77", x"06777e28e03d0f7c", x"dc5bcd6fb324558e");
            when 23324937 => data <= (x"51bea5afa6f4e7e4", x"10e7053fe183061d", x"f8ecb6b6fe06def2", x"dd61ae8c02dbaf5c", x"09163aa4aa02bff0", x"fc86c0c170919b68", x"60e9a745b6ee675a", x"f9fee97852fd8a19");
            when 17197905 => data <= (x"501d5c885c0e0d9f", x"0b87a97a41bdbcfe", x"026057f3247f75b0", x"f1333a52d71e9fbb", x"537292a8c4f8a2a7", x"58513750b78031f8", x"aaf2ae20117d81bd", x"add4483220b968a3");
            when 16359466 => data <= (x"c42a736585829a75", x"443079bf5eb46bcb", x"c066f7fda8541f3f", x"1fa9ed3e6368eeff", x"4cf32d9a5561c133", x"3ada7a7d6d132ac5", x"de1441df45b6a68e", x"7d0ce5cd93675e96");
            when 33513406 => data <= (x"c183f389b8ab49e9", x"5750629cb0548752", x"6ef065cced00ee1a", x"9ecb223e6ec474e3", x"3d4f449f98f1a15f", x"35b3eb1da7fc9c7a", x"1d09601b8b75b262", x"96c23fd17e93803c");
            when 10776867 => data <= (x"6af137260815e908", x"4e56a0d2dce49e56", x"5f9b17d14abc0814", x"4651ac570295d37f", x"a81410041af8592d", x"1b73e269fff8f445", x"567f317814cf03fe", x"785f97e0df1e9a33");
            when 32633290 => data <= (x"f3be50ce1707e856", x"f4f4cf79d5757792", x"f79eff0dace7fa24", x"68dd97bd8e36242d", x"8530a21085a780f3", x"7e9ad0b49b03723a", x"f431ce9eb86c3275", x"6858b4d48d501d15");
            when 15010107 => data <= (x"1357fc552efdb9e6", x"0b0889cd68c09731", x"9186f8b360c285d6", x"9ad510249055bc41", x"a620d5845a763fc1", x"d5266c9b3d165ba2", x"bbf0ebff203398a1", x"c7a4909306b8e5b0");
            when 10094106 => data <= (x"b72691dd1ca3e13b", x"6ed9f28a2773d94a", x"48d18afbf30cb01c", x"9aeeb1d778911610", x"e3447956e86052e9", x"f1ee9dad62086118", x"cdf9779bf0b786bb", x"2bfa8725b2ebb437");
            when 10970904 => data <= (x"b6e41920e4bc911a", x"8e2ee37e1019228b", x"b04de7c26cab8dac", x"e8c886ec3ce22938", x"13d3e51fee907557", x"0fe0b985a3193d81", x"ae178b89a9ca35cd", x"68759123376c831d");
            when 28172547 => data <= (x"843eef2421e3dc3e", x"5ab637f679499c7f", x"4a264330ffe3e930", x"28d6ed8cc031a781", x"8f378bf8b3e4254b", x"6635d8e57f56725f", x"e5a52304fc142220", x"9e3d49bcca86cf42");
            when 20719907 => data <= (x"74fa772aefa2aab0", x"59e720f2618e8a02", x"da3f6938cd2a6746", x"87530b1860cb7e45", x"9f03bee9d6de1743", x"6fab967cee2da6c6", x"154ae2e2f33a61fe", x"9593fe486e3ced5c");
            when 27226513 => data <= (x"901ca0cb4530b3eb", x"30330985da364896", x"11662f8ecc97ca18", x"15d6777f4f31e4f0", x"ddc6a8cbb947463b", x"5ece30c3a3069589", x"19ffd9ca7229a760", x"ea1a0e0cccb561bb");
            when 17580915 => data <= (x"1134e0fd27fa5b1a", x"57a751da990ececc", x"26f5c416a65f1b03", x"904f042058405228", x"54961ea2fd5d708b", x"75b43ef5f75b853b", x"edd88492a581d1e0", x"22776541498dcdf6");
            when 30301893 => data <= (x"5c7d02d0b3629ea9", x"b63c122563e4340f", x"79990b6db64c343f", x"91d3e14187ccfd60", x"0733daf101994ad9", x"294bc78b22d0996d", x"a4ef2a15864083ee", x"6f9b84354c0e57f9");
            when 27847640 => data <= (x"31aeadd2d24b9d6a", x"9b5c08862fb124e3", x"3482006689935219", x"63ffac6d8d6b2c32", x"fa56373adb9ebb3d", x"4d0eab94fc6826d8", x"a17dd745fae58e85", x"f90b9548939ff43c");
            when 22954242 => data <= (x"dca9764bcefed4a9", x"2e3a7cf88d089fd0", x"ac15469d32a575cb", x"bfa7a7a8fdc9a982", x"2018758487f93d1c", x"a660b1cb73e39b34", x"fe0e2a430f2e8e9f", x"50a41cc9a7957e98");
            when 10347882 => data <= (x"7cf13989ed7f376b", x"eef454b7e5d4de48", x"66e13883d038f276", x"df82be23e1af4386", x"8fcb9f9da46429b3", x"c6eb884516fef802", x"52b749be905f0ef1", x"d164fb898886047f");
            when 23091132 => data <= (x"baa6cba5eb6f86b3", x"7f841efb5fef48bd", x"4c56257899a74025", x"ba21906ae2264cfc", x"5d2117c9d0638b3c", x"af0dfb986469e4d6", x"1e9f451eb8baf338", x"6e9744dc1ba7bc9e");
            when 6194585 => data <= (x"435b2e52ee8382b3", x"844ec001197b0bf4", x"10416da767c54ced", x"e0a87efb6224242e", x"300a2ac75699ffad", x"a78e80ed189c8233", x"b5ab6d1f92fdfd73", x"8a22898ad2b3fc8c");
            when 26344232 => data <= (x"7d768cccb9fc6013", x"15b04aeda4f3f0c4", x"190d46a10f8af923", x"8f8e6b93b05ab475", x"1eea49ffe3e02ebf", x"6a8bf4a62f979a0b", x"56242167633e6736", x"85faf69549e2c7a4");
            when 12780113 => data <= (x"98d89285af4a9bf1", x"8a4ce06a7d74d84f", x"0048178e41d5cc5c", x"79c6e6e0e30614d4", x"6a1bbf0eea3a412e", x"8b1b9568c7e223d0", x"0bb66736fc9bd1e8", x"a632cead5afc4fdd");
            when 3754758 => data <= (x"d146dd249f7703bc", x"68ff368b1b97a9ab", x"078d08e6912565f2", x"64d83f152a3ae93f", x"efc5bcee4f402a58", x"4397f625adf77023", x"59fdd4853298e9c7", x"42dbf6501e24adfd");
            when 13470478 => data <= (x"da29da4efcea8867", x"5993afe38b6d8889", x"e59c569570cee5dd", x"0e1e2e0d6bec41f7", x"5825819149b7cf43", x"06322968d403f3ca", x"23de6c3fe3677149", x"0d2a5d195d11ded9");
            when 13336499 => data <= (x"15fd6fd90981d7d8", x"b167831db84d4ac0", x"99583c8995fdd847", x"50010da5436e63bb", x"9393e62eef9ffe84", x"c7098f0f9e49dde6", x"5de3a01d0d48ee00", x"a3ac742282dd2601");
            when 5746532 => data <= (x"1cfc8ac4f570f95d", x"9f8de9296d9300ea", x"61524c0307cbf9b0", x"d1b73d18b0db5204", x"57bbb0368a47ccf6", x"dd24b076d5037aae", x"cea9b1ad572fdd61", x"73c15b4b1156a1d8");
            when 20834223 => data <= (x"3f96f2b1442d2fe2", x"efea1f79b675c04b", x"4f1d89fb6f10a35b", x"cabfa370d2057ce7", x"add63616fcfa8cbb", x"3a5f97e58ada153a", x"16478d4e6c565f0c", x"d00a1395d78729ad");
            when 9445096 => data <= (x"e9d6fa1a92f6dddf", x"a948d7273fef8601", x"40dcd034be2d1afb", x"8b0df7723b1b1a5f", x"b45256a2ad4b3584", x"7ec9238182a60519", x"5a0c4b5bc15b31cc", x"8620ebef1b987d4b");
            when 21441445 => data <= (x"e5addd1dbe20d7df", x"eb0f924cb1afc0c3", x"dd9a4f3b82b51b59", x"882d8531ddb1c5f8", x"9914e924f681006d", x"7458672a828f6d97", x"db4a0877e46f8c6d", x"4eb8a4ce897653f1");
            when 4876890 => data <= (x"062019b0ab7b6d61", x"331776e62de38d4b", x"ae97d3c6f234c6d2", x"25a121c1dedc6d62", x"baf637e82d99a848", x"8957bf7f5582d644", x"d804bd991bb0ee31", x"0f1f2fb53e6f685e");
            when 20327868 => data <= (x"c6a6df87a161b14f", x"95083129928ed012", x"bc8e4e63997c9b2d", x"184694ec43cb7bba", x"3925a5cc372fb5b8", x"9e82950bf5f7d807", x"3477738425fc6ee5", x"b9b53efdbbcc6881");
            when 3610861 => data <= (x"a460b70f8cdd609a", x"1ee3ff7bc84aba33", x"5570cd9d9f335114", x"a74972dfa3d0affa", x"997b75ffc2ffadca", x"579518a0f6504b73", x"c133c5d428d08d91", x"944a8c3a574b1a7e");
            when 31544061 => data <= (x"b42b392f95896b4f", x"1d9756b301da2990", x"1ed8da04fc04f01b", x"cb09542890400633", x"2405d2757d15aa5c", x"0b2a37c9e57c36b1", x"8459d05928128c15", x"d6351750cf8cbfe1");
            when 33391751 => data <= (x"dc5aef7e2c0717e8", x"53debbb96458fb6d", x"3d054e76562762fc", x"137cd65085eae587", x"ffff5eb96724417a", x"a2f3f3f3c924e029", x"153c695c9be78c82", x"60e5137d3f475d49");
            when 7513493 => data <= (x"2d7043caf1541fea", x"642aefb8a4c3d01a", x"c94d4b243ca515e0", x"24d3539accb23e0c", x"140dacbf8d05893d", x"9a94e5ab84cd9223", x"3470897c614d705e", x"de6722d31b73243f");
            when 25784292 => data <= (x"0894acc2a2819c1d", x"a83b743ab99cb5c1", x"bdda25cfc3cf14ba", x"f884fef4619ea77f", x"242427ea31480367", x"3c380af471cbf4d2", x"55c2467dc8f7c06d", x"cec1dd21953cb7dd");
            when 12563951 => data <= (x"e15b92bca73d5cea", x"07f98b5d807bea0f", x"6eeeea0a974b408a", x"a526cba2525eeded", x"d1112db1718f7f52", x"16a1e4e72a4052e8", x"4bc47f30926969f8", x"05f170599cb33545");
            when 1376644 => data <= (x"cf2e9ea0b6abc95d", x"a446e01863438347", x"b06387888aa417c6", x"08056688e835910c", x"16d42826179cb5b3", x"60c5f560e2f418bd", x"7ef2c6c168254bc6", x"86d49a9ddba242bc");
            when 12779030 => data <= (x"4491f802dbf74581", x"b3ab2b82b53eedad", x"0aa6b29fcd0e4333", x"2406744f00731d35", x"36551397d854f3e1", x"6e8788e49563472e", x"4e8577d726f70403", x"8e7f10095a2f5fc6");
            when 29401351 => data <= (x"7c3f14aca58860e5", x"75cfdad1344bd316", x"55303970008dda0a", x"43673bda5df141b2", x"072c275e2d227810", x"0fca8938d173dd87", x"17e12bdae9949fb6", x"0347a334d3d4aa56");
            when 28080086 => data <= (x"59f9b423bc8415b6", x"02990f79b9999ad0", x"22dd5351b3787036", x"9b7de9cc7a78542b", x"0e1483090219238b", x"8fc06a0ad9ce80d5", x"93be29dc8784557f", x"672927d6dc8c6347");
            when 27394549 => data <= (x"fa3c80a5df94dfd3", x"72db44910582ae57", x"aea2998eecfab444", x"e955b46585101705", x"4f6b45c1a30d0beb", x"a778478aa425855a", x"0c73101261c4bb11", x"a07b39494041069a");
            when 31280601 => data <= (x"0750a0a0360a44e8", x"8a0928c26f9a9ed8", x"c0fc312429507f84", x"3353c1201bfd19b2", x"54d4a83fe982d8ec", x"b33a472b52f99b69", x"1ef26ff9399fd257", x"6797abe3e549399d");
            when 23218837 => data <= (x"59e7cd00fd0666a6", x"2f155074d86c586f", x"2066494d091810ac", x"88e5991eef78c07d", x"9fd923e80a60c622", x"96c00e9fe163d830", x"aaf4ef187645b437", x"8943e15c158b5944");
            when 15174181 => data <= (x"b3385a3ee64dd74f", x"4dc82cb89fb5b02c", x"c59b43d5947100dd", x"c2ede1da381d7251", x"2a12cdd61bbecd5f", x"4e9da874d18a065c", x"4f968ac00c809402", x"789089dd4af41fc1");
            when 27276643 => data <= (x"d07d69c14ea860de", x"d40685a08555403b", x"464f3b53f5032517", x"359a1de05b1138f1", x"9d12359e6a96a71b", x"7a25bb1f761f76dd", x"6983299f939e6647", x"c887cb3b9158f5cf");
            when 28045317 => data <= (x"df39d32c58929ab3", x"38bc67fa797303ad", x"47fbf9c909130ce8", x"732143b89f473364", x"c49fcc3c2535d521", x"f36d4883177f49a6", x"be566ce3d6ecf619", x"3c7cae75c2cda953");
            when 32526619 => data <= (x"cc0da05c08a78f2e", x"c4ebd7b53631a2f2", x"57afdacef77feae9", x"0e4c76b8f3c84bdc", x"169101d7254ef50e", x"63ac69cce66f9d30", x"b0476f3025c8d195", x"f59e964988f33ef4");
            when 26401876 => data <= (x"8fcd327dcec4b697", x"0d61e7cfdee7640d", x"198939875f55336e", x"166d697dd3034e7d", x"8a1597ccaddcf7b7", x"7bbda164b8368c2c", x"fd4304af1661ec18", x"30be5e0ea08609d9");
            when 26694564 => data <= (x"74c52a642b7ca99b", x"ca84b2364e8d2d1c", x"1affd07191b15adb", x"8b2880ed7c464942", x"98a79531edbeae45", x"2e49703452b16256", x"e926ecdacfea400a", x"9998951f94d08ecf");
            when 30938222 => data <= (x"d26f6e6f227c7225", x"c5103deada6d21b9", x"bc8a66ea2b4ca4db", x"fafc939db064ea75", x"94751c006895c29e", x"7e2f5314af35a92d", x"71d01a23f8b32036", x"6ba6ac9b44bd5bb9");
            when 2147791 => data <= (x"f8db7331bb8fe33e", x"30a03e1862f7352a", x"383084c0464a2ff7", x"de68ea8eac5dcd69", x"d84abca22b9b6769", x"abfde53f72dd87aa", x"4fb89d01cf9cc39c", x"ad00e95e42c17280");
            when 28390873 => data <= (x"09ac5ba3e40c29a2", x"e07b0629ab28b430", x"fc5702cf76f14707", x"d72379f6c0848739", x"2c6bf8c6da01b7bf", x"2ffb438de9907392", x"863eb35d972a6ea8", x"a0da5e819dbffadc");
            when 8147115 => data <= (x"ecaa0ca6591b1bdb", x"2f761fa5f310316b", x"3f3aa63a6abd854e", x"58c181f14d282bf2", x"076ec23ad96172a7", x"92d20a7840b628bb", x"c07b369ecd4062e1", x"e2a8bd61e7d0fab0");
            when 22940993 => data <= (x"8c09ffa92fd41d01", x"5427dba1727d726e", x"165a483d84d333a0", x"627c6e65030eedcd", x"a6d875f54e03a1ef", x"bbefd3422c7b716d", x"b6d3a5a81ea029bf", x"0d04642d56bd9ae4");
            when 1608309 => data <= (x"da714c97e2be8e79", x"027e926869de19c2", x"3decf70feff8c28c", x"b6819aa793aaef7b", x"66dbb7cb5abef676", x"32afac897ab8fcf9", x"7d82c14c0454e0ee", x"0be5b4155dd49342");
            when 18341825 => data <= (x"7efba4a8686c0c3a", x"0a392fbbd6b7fb1c", x"0098510059c0054d", x"e93bd2c98f341c3e", x"9eee0e648a6c7262", x"6532c189b6ae3563", x"96d4453da61f585a", x"b61d12173df6cec4");
            when 30732673 => data <= (x"b03cf6ba20d70d0e", x"9a3de5dad468c6bd", x"f54520d1f9a6a284", x"9faee42059d83b64", x"4d861b301b6c61fe", x"52b1f741622e0b28", x"81ab24be5463e132", x"3b8202a7662dcb6d");
            when 33755426 => data <= (x"f851631b3c376065", x"cfb711b1a81a2507", x"43434499d7dfd5c7", x"2f77fdd9a59ef80f", x"d7ee168dd75b7a48", x"74a44593749d7e49", x"2da530c2ee41e060", x"e6fcbd3041c94351");
            when 8031912 => data <= (x"90095bd5ec96d872", x"a8aa640d01001294", x"0e280bf613bd85c9", x"13f5486cb92b08a1", x"c87d4d42dc8c08a1", x"f8b1b6258aba2c37", x"a21a8c2b78928891", x"641d42df621f6311");
            when 23491041 => data <= (x"33e208e3f848d496", x"0e67793446750f08", x"ed8ea41c7c7a9bae", x"7aeec7f369216eaa", x"4242b2b33dc6cb09", x"051f9907c267ac08", x"6237e53a0eb84f9c", x"a1338735b6f22721");
            when 1549083 => data <= (x"dd034ee2921d756a", x"2139002d0f8a6a91", x"04cc0fa0bf0f81dc", x"4ff75e447fbe55d3", x"7e7e34ff37bf2afa", x"c8b9fc2df9b4644e", x"a102b2b14f6e6788", x"12931798ee309a51");
            when 9624505 => data <= (x"c6ea6ad3e229b188", x"a7c6667a12006e37", x"e7ee2013465a2c67", x"54aaa5390ccc0b68", x"0b5746eece2ac114", x"af4c503e87561608", x"33b4b915fc8dd564", x"fbb8630d824c5c60");
            when 13280181 => data <= (x"fabba55952408782", x"86be14594b7ff52f", x"e40b6235c862c06c", x"b14d4fa80ea4207c", x"18e8db910cf901a2", x"8039be9395ed596a", x"bb4918650d64f3ad", x"6ce370df74a4dda7");
            when 20962357 => data <= (x"5ae559888fc64ddb", x"b602d928e7168ff1", x"8a3ffbc41b0d7a00", x"39c717d9f0b196cf", x"c8170ee52a1a155f", x"df0ee718defe85b9", x"9bf0886624767b4a", x"618b12f80bb5cac2");
            when 29144206 => data <= (x"1cd6e1908585a190", x"3ea483ae753dca69", x"94b0b85780757488", x"8d451d0e10d8dbd5", x"95474f00b5650d4a", x"0c884b3ee3aab6b9", x"1ace5aff0390e480", x"b513331b64bd6778");
            when 551700 => data <= (x"bf3586a6b8bcca9e", x"04858dfc4bcdf2e8", x"a363c8d824eb9630", x"ab8cbd729ccdef60", x"1d803814900c3d31", x"b82099c50901128c", x"c33d8ee9382ade77", x"a3fb5b372d7a5b7d");
            when 31276659 => data <= (x"e51763a4dd5a656b", x"057eaaa216d710c0", x"4be0c11962fe4e0f", x"35f3af7348f6bbbd", x"a7e32b583c6098d2", x"6774dbe8fa8378af", x"7e4b7a225c151080", x"536c9b3443e9488d");
            when 17650296 => data <= (x"8319feabdd7f38a9", x"a07ee2338032ea44", x"b65094694ef692ab", x"c8f3f7d9ca0d974c", x"2fd6b8a974ee6fab", x"23aef5a06c70cc2f", x"32445832a15998a8", x"211819e66115f585");
            when 2640547 => data <= (x"c8bfdaed682c7bc8", x"44d66145a368e58f", x"3df0fd0d5b1ffa70", x"2ae22481a51e72b6", x"8f513b4c35b4b634", x"ba766ec4a83b1c20", x"fb8062bc8f7bab02", x"97968b8d7a18d1b0");
            when 33451874 => data <= (x"751b828ddaf6ea0c", x"6dca02b5a2f49812", x"c8cb9117f4da7944", x"b16d6a0a7fc85623", x"426fd54c01932d2c", x"4cb6e19af627e9a0", x"ed14625de5eb1e3c", x"3c6c8613ac3b3a88");
            when 10813563 => data <= (x"a731e09bb499be57", x"18a3548495946a08", x"e321ec6a3c0ab40d", x"98a77e1d9d69c39e", x"53f9c1c7437e8970", x"4abf462aeac90756", x"8dcd3e4a99005488", x"788789d596cd7898");
            when 10581618 => data <= (x"ca61cbda6069f642", x"599d99caba5fdb36", x"ddcf1fcd6a0e0463", x"968b1193fe442e3a", x"7375675f9a139a45", x"035d27c6f3463355", x"0a1f911c92fd901a", x"7e81bce08e9aac70");
            when 15978992 => data <= (x"1b04ed8e200ece6b", x"a619bef99224ff51", x"7f5df6cb333bba75", x"b4bc838f8f9991ea", x"b4256c255a4c35d2", x"4c9a14cd071cd3c8", x"e3ea235a9e58937e", x"5547400ed3141958");
            when 9347288 => data <= (x"2be9ac80c4e3ec9e", x"2c069d03ca1d8cfe", x"af3c957bd2c37249", x"de9652dec7505d89", x"8a622388aa84a4b9", x"0152301dfecbf601", x"29442184678fa0dc", x"f234f047c07ed76c");
            when 2030972 => data <= (x"b154c65b1e63924f", x"4a6b02abeb10b726", x"a82569a95a972bb3", x"f20e4aee2f4dcf8d", x"0ac4d5dd9850a316", x"5aaca3dcc81a779b", x"c2cd955809674b76", x"b31a43610da339aa");
            when 8797092 => data <= (x"866cd8a4b3c8ec97", x"e2657e082dcec8e5", x"9d00de3ca1b61c6f", x"036d29a765f1945e", x"aa6f068663ec9b46", x"5db51ffb9e6cd43b", x"26eef9d490d0fd14", x"375f523e2d0073b1");
            when 2137907 => data <= (x"8f03e8bde8c282dc", x"6118701c5644e1dc", x"efac13cd5972286b", x"8d18278d33e05915", x"a19ddc26200beeae", x"bf8e95f131f03ef8", x"a5cad1237fafa6c3", x"991d6dd16b48b0cd");
            when 29684118 => data <= (x"f9fb76b3beee9a30", x"17305c00ff5762b0", x"4edee08d84761e3e", x"620d8cbd047589df", x"1d6ba12b419ac7b4", x"5eef5b2ebd83d3b7", x"c5935b1614e9e244", x"d966110c821609dc");
            when 17217942 => data <= (x"89100af0a9b62cbd", x"1c123127756ba184", x"2531c1ab3a8149d6", x"766b891450648a8b", x"8c15c8c451d919d6", x"6cf964b8273dd102", x"ef2db31028019f1b", x"b5aaed928a6790a4");
            when 540409 => data <= (x"49102f48dbad23a2", x"981a9425378af674", x"0048fe127e0bb644", x"aa7192323eb59d8e", x"e3d93d71636a2c1a", x"fcb6a501ab754ad0", x"dc69356ac6013e31", x"19dc98db593b7dd2");
            when 10789176 => data <= (x"b77ef5463b35f819", x"140af2bfe8c8923c", x"0b970682da00dd66", x"b84ac78fadfd773d", x"131bfd8c2e01d0f4", x"caa9371b5eb28fda", x"1396e0cf6c00117b", x"65c8806a1bd748c0");
            when 22790425 => data <= (x"8b7b3128eb7cddcd", x"5f3eb0445263914c", x"43a523b4a521e9bc", x"3dccdc665a3f506a", x"d5553cb13af15a5b", x"c3eae6ceee556dfa", x"97d78fa2631719df", x"ff235961eece198e");
            when 18652627 => data <= (x"5470c243a2be254b", x"7cd7ded160c4f1d4", x"4611f792664f9572", x"faf4bec6f2e3e170", x"73acad25ee910360", x"c0294853cd1cc8d8", x"f67130e65359daee", x"cb75172a6d4354de");
            when 21899930 => data <= (x"3e1499b90e029854", x"358e6107a4edbb71", x"116de293697a2626", x"ed0dbf495fc8aa50", x"a181a55da549df68", x"e45ab50f891428d0", x"e24c47b91575822f", x"b1ac08140615bc5a");
            when 13959143 => data <= (x"9e3de5a5038a9fc4", x"9b28f50e4e5f3db8", x"5bca7b536325a791", x"86f934b8ae05bed1", x"db275502af571624", x"921c85d60a1b2d2f", x"69a739993a593754", x"752a7b8dffd460e9");
            when 32859039 => data <= (x"523da9613444b4b2", x"656defbf4266b488", x"63e2ddcce4785cb4", x"fcaa8cd072c0d059", x"7290228980669ebe", x"c378b1f6c105cd6e", x"31798986becb06bd", x"6e0be879e211d88a");
            when 5722677 => data <= (x"e59fd30ca36e9033", x"df4decbe7b98b7c3", x"b4e1190eeea991c2", x"403b3816069d280a", x"e0cc676047bfac4f", x"47f1602f108c4790", x"8128bd3cbafd1c1d", x"aabd99aca47bbe48");
            when 28713534 => data <= (x"3a9860f6c9d4bfd4", x"f2ec8d1a1a72f094", x"54a738cccbff33a6", x"a9ff7ebe6ac8cafa", x"b31a74da04c9b1c9", x"5234589d01a3e1e2", x"f99405312280e5c0", x"14d63d545f7b49ba");
            when 10276843 => data <= (x"4b24fa38207ffea9", x"f9572e38b56def79", x"f928c603afb229e8", x"dd07b0facf7841d0", x"c10a0e0937999de5", x"e88ac89fb8b19a03", x"e97d5707f1ca2d9d", x"6c45eb89c5073991");
            when 26935244 => data <= (x"355b6d9e0c0012a7", x"b9031de541d90004", x"f4aac05d7a062e3d", x"7826e1fb210acbd9", x"ae5dd2ffc72fab0a", x"7388dd818d958864", x"649260f9a25c6cb6", x"e203be955173fbe2");
            when 6744758 => data <= (x"1def3fcb9da58f78", x"216559e79fc74494", x"0ecf5fcaaff07a9e", x"5741800a616ad20d", x"94b7b37fea9c8bc2", x"7998193c8d12be4d", x"3baa01d6813a0e1a", x"6bb9a1359abc60c3");
            when 2139469 => data <= (x"ce2b1ff1b6848fc0", x"9e4651016b2e2a0d", x"db44c195d709d142", x"199142969bfc55cb", x"7b3d6a29f367dff7", x"985c852bac696bbe", x"da0c75e2c9af03e4", x"715deca73485940c");
            when 23036575 => data <= (x"8640a249a686d08b", x"ac171bd7d6d4839e", x"80386834c91d1f93", x"35a44c2ce03a0b0d", x"7b4a7409c5cdde51", x"f0af7e5603d17dd5", x"718906a264327c4a", x"f45cf8d821ca7fce");
            when 21846887 => data <= (x"4fea1474c083ebda", x"34c131dd86785190", x"33e7417f56f5fe80", x"ebee2a52cc6b2901", x"9ece3fc8eb91d420", x"23bb3dedcec25da9", x"bfdf9e40f58856df", x"bb812c751437b977");
            when 9850469 => data <= (x"eb776e0430bfd820", x"d20b63561de6cf32", x"3bdb74af8ea2369e", x"19554e15dbe1dac4", x"14671674afc9d2e3", x"6867044b89d79d70", x"22ef2600903dc528", x"a8504134781f6cb7");
            when 31169993 => data <= (x"631c7764755c1a67", x"0dd58f713c0e6979", x"2c4cf90da7d1898c", x"72a8e54644854406", x"1577f1317e609c01", x"9fbb2dcaffe94a38", x"dadf7d1f9be95496", x"b3e4f476c64520ea");
            when 8999444 => data <= (x"630936e82f555051", x"7056419b7f51c2f1", x"224364c731fbfa9b", x"e152856594368042", x"fb2a8f2c96b4eb1a", x"b0d13afb45cd98e6", x"b1a8082844daf568", x"107a60f14e58118a");
            when 12652389 => data <= (x"b77a14017ce27eb5", x"b6e3ea4625025d9c", x"e250dd519a6c2ce5", x"e6b3bd0c1d546ec7", x"896b7f6bdc6bc854", x"7f2af73b591c7919", x"56385f38116ac37e", x"6a4e4500d071d23b");
            when 5582287 => data <= (x"507f421fd2a3e8e4", x"695834a887a8106b", x"ad2e03190100354a", x"3731739c039a357d", x"b90aa5014ef9e93d", x"a4f80c83cd45e186", x"8882d4f4ccadfe47", x"6b19ab2a60d6ec24");
            when 13121633 => data <= (x"e0c6932f393010cf", x"1498de52c04c61a6", x"765e2a7cf0724802", x"883a484b68adc42a", x"d9630c07a456c028", x"d797dfb649b828a2", x"8de7938b2d3cb2a2", x"ad51ad397f3722d8");
            when 12007298 => data <= (x"cb0895842684cbc3", x"383be6f8c7e51c37", x"b21b39cbd685e12e", x"8af9fc13d0a5267a", x"9e19db3dd964f47f", x"2a1d712b3ef49c37", x"9aece66ddfce5d35", x"d7c1ab642c8d7a83");
            when 25785652 => data <= (x"71ec3d922f610d47", x"d7f52df6ed7cac90", x"5338968425a60aa8", x"79c66ffbbb16e40b", x"8f225f952c742501", x"c5934fd32869c3f2", x"349127d2f7d1f1cc", x"fd30bd0f7972320c");
            when 27112906 => data <= (x"bc4851e83000ba62", x"e1c84076eeeaed18", x"42972ee4996fbb5e", x"1a692bc3e7b03d22", x"9a4842a9ae8f116f", x"25a59b389640b202", x"1c096d5a4b7d43e5", x"75edc80315563b2d");
            when 10358450 => data <= (x"0c86a08ed9f3df17", x"df37c526965fae00", x"4b15201715ddb5be", x"2dfaf457277f4ad2", x"86017dc9d21824a5", x"a67557dc9cdbfe25", x"d8bd7d7513cdcaf1", x"f17a841aedf4c6a2");
            when 17419212 => data <= (x"f393be08ade2940f", x"471bfc2fc5d8062b", x"ebc0d0253e2c3b0d", x"db66ef3fb59b704c", x"e4ca00f1cd857910", x"c5e4cef4b6200f93", x"f945a90763d14e76", x"35326d2d88a20245");
            when 13693567 => data <= (x"707fd65d1d646db8", x"aca2932fa810dae7", x"c972b143b8a47bd9", x"17c1604aef9ed94a", x"4c617bd861d6b32f", x"0ad7c1625e77e801", x"4e40a7ccf9db0300", x"6b6154de38e457ec");
            when 14497770 => data <= (x"f7a16d17a3905ba0", x"9640209174fe000d", x"31579ddb0cb88920", x"b125b73c902aa701", x"0a52b6924655d617", x"c2977db13e1bea8e", x"864d011c48c04b13", x"88b803b148ed2aae");
            when 11752199 => data <= (x"89a1f37aba034ec9", x"493804cf500099ed", x"318b4f0f4f318f7d", x"2d12f920b2329527", x"98cd22383a85866c", x"43cc0028be46d61d", x"308172209bb84a18", x"29b112cd65b1a0d1");
            when 26486827 => data <= (x"3150be85ac6bcda5", x"496360363941c7d2", x"eb0ca4a346b68c9f", x"7648b7f4cf799b13", x"09a7da3e516df6d3", x"d521f6d2fa49b83d", x"b333d962813db072", x"898e60c76a4d4771");
            when 16118840 => data <= (x"fc6fece5ee4c7c13", x"f62934ff94c897fb", x"010d3db523497e40", x"fd13b3c67c1518f5", x"ee0a35be8782be05", x"ca38896489110860", x"9830a5fc0a9e5a3d", x"562592d64a8a1df5");
            when 27977288 => data <= (x"8f65a89a7c8d51f3", x"581fdadd25092dc9", x"3ee8800603d63ed6", x"34fb601cc0487df9", x"4d2bb21a21e6b47b", x"283d44bc52d1b89d", x"3b747e93853d9ce3", x"13fa57b92ecc7694");
            when 3777080 => data <= (x"9aa0214dd5d80fb6", x"61dc2aa79d589b8f", x"d9ab8ea6eb6d8cc8", x"6cfc72205258383f", x"39c255e2e3de835f", x"a1832147e11a7e36", x"90dcaefeb4382241", x"e2c782c837cbe73e");
            when 30624365 => data <= (x"0aac0dd62a1d9c3a", x"a4b13d4627928d8b", x"07e27acfdb7dff2e", x"a49a40b9890e6c46", x"15548f16dd3ae7c4", x"d71e697fa570110c", x"515196e6357c9747", x"6f8f02f3c41a4337");
            when 12427860 => data <= (x"8ca38a513de5c6fd", x"2c9a3ef87b3ef5e5", x"cb8867c9a49d2e4f", x"71a49f5663707230", x"4d17a4faa55e1f89", x"6f8b743083ce696b", x"dad9953b96fcf5f0", x"83da2e4517ebbc86");
            when 2350172 => data <= (x"31c1d1c8d3e3cb35", x"b378f6ab128b9d83", x"742dc1039f9c59ed", x"204deaa4133975cc", x"f8e96fa2206ea7a4", x"6e10b36777108b84", x"b4ef951634b77e6e", x"079721bcf6161703");
            when 26051680 => data <= (x"8cbd1fe61322e2b9", x"dc2d8903596f2297", x"e1c6d8d3c37af49a", x"514115e6086dee92", x"a3f706ea41d561c3", x"759085407fb9e31f", x"6da848ac608f274e", x"47e597295240c634");
            when 25527354 => data <= (x"911c387fc8c4e3f0", x"a98b5ed0773d938c", x"7e9c3c9933996989", x"9cab6849f84f6cc7", x"19f929df1789bbc1", x"497b34a22a9dba82", x"a81743e77ac1ff4c", x"de1e07dba54f8e42");
            when 6610422 => data <= (x"9bdc301d7c6bbfd3", x"efafd4f02c445729", x"9a5fc793b6001d31", x"411e2825ca458b8c", x"cf81c8c9140c8831", x"3430bd0d7148bb13", x"c124cd4899451014", x"28b1cf97f994c875");
            when 6408313 => data <= (x"7bf89df2c6e144f8", x"af232a2bc6248ac9", x"8d88415f118fae12", x"7137030a68f787fa", x"2bf13b49735abd73", x"ec478deb0c65d5bb", x"162694d22ba7cd50", x"ff6fd06967dc43c2");
            when 18053141 => data <= (x"cdbe361241cca6b9", x"8a7de9ca7e7f1640", x"4e63a553f11aa0ab", x"ee5f15576ef2dc0f", x"e49c7bb4c567605e", x"d2b06fa66df0fd20", x"ea0ecf4187a801f7", x"605eaff17922a1df");
            when 16979545 => data <= (x"40b4510ec662af32", x"7d1866909fc051c1", x"cd821f22d37d972b", x"084d29bea630b41c", x"911163b51dbbfecf", x"b8110b23393c75bc", x"4825110682d217c0", x"58406ffb1513d00d");
            when 30086369 => data <= (x"af8fe089ce4ebcd8", x"854e5ce86127a32a", x"c48af159cb55ce70", x"412c993d48b93f5e", x"bc0695142d0c14b3", x"2bf0647e1f3724b3", x"f0c9445aa68fc085", x"c73fe392ce8dfffa");
            when 7670088 => data <= (x"181325762b8c2163", x"0dc281b6e0ac6f32", x"7047186b10f0af5e", x"d62c9929f2707942", x"18498fccfba28d35", x"cfe9832a1989f0f4", x"471d4e56558b62ab", x"af7a6d880c83d23e");
            when 2548669 => data <= (x"46800a58a3a35c8e", x"ce5f40faa22d697b", x"49df0a69b9184999", x"70bda9124fd07b97", x"836a2bac05a09d98", x"4202922b5ef229da", x"881b17697196f930", x"fb9bdc50c7f5f6a4");
            when 33539731 => data <= (x"bfe24a8487fe3b2e", x"c6bc60bf34d687a1", x"f8cabcaf84293d57", x"a921abf3d757d224", x"9321cd8006c1f5ab", x"28c5d5678fd21025", x"50977ac87547d43f", x"dd86f546bff77ef4");
            when 32077625 => data <= (x"c628062029bc074f", x"1bb409a7ebede44c", x"14873f817d35580b", x"6fe33b960f0f8146", x"babea51e051c442a", x"214431f4e09b1686", x"dc5db178f5373e43", x"91fe45ff168528ba");
            when 33045620 => data <= (x"75be809ef967bc2d", x"f574d0bd5bbd3995", x"8f8a26ff896d6faa", x"a795d0de61aec826", x"3833cc5a33d4a687", x"04d34669ce2c2c6a", x"9916f998603dca92", x"30f616d07faec24c");
            when 18908661 => data <= (x"b46de1eebf91750d", x"443c9152dfb36b89", x"3e56d5e291bf01fa", x"7134670d3daac8ab", x"d9cef546df36a545", x"66e9b6d5fe586ad0", x"4b5016d6a1adf2fa", x"c06273ca63410a44");
            when 15219150 => data <= (x"a201433d4fb496a7", x"192dd880c8fd433a", x"bc59d3888b5957f1", x"2bfea6b4c6b68699", x"e33db579f057204e", x"964f9f5d5091eb4e", x"08d359b49dd7a950", x"0fec4758da7aa821");
            when 7888216 => data <= (x"53c19f66f26e4c02", x"d5f687304ef220d7", x"0dc7c59441d3fa7a", x"e96e41dfa71dc83e", x"b738b404afa4ecff", x"e5031978693b0466", x"13b18510eb9d53cb", x"c4c40a2a5cf350f9");
            when 7181645 => data <= (x"2567019ad421ed0a", x"fa54ef411fbfe488", x"093ad482e5a3863e", x"a629cbc0dcbf0e54", x"dbb5ecf345ee10b1", x"107b32f0d3ccc2c2", x"c39d11efa68c0824", x"fd7ceb88abc33405");
            when 27962521 => data <= (x"2169dc9ee5def8c6", x"8e88f47c1246e6bc", x"a434c40a61ff6034", x"8606147b1175b3a1", x"23a023e49fdd5387", x"aa115439b9748cec", x"38c4e77a1857d0b3", x"8c0541ca36d40916");
            when 1898701 => data <= (x"861fd283c1e43b16", x"e4b45f62ce1c6353", x"6b0ce8f6035660d7", x"8f09e4680f6cdf4f", x"7b8d418fba7a1200", x"85ad3c08f4773ab4", x"34ff63f63a3715e2", x"c3bcbee53f2e48f9");
            when 26069058 => data <= (x"dcedff458b898797", x"7ed97453e455cf6c", x"228c1194d6b28a60", x"bccd575ebedf0cce", x"971ddd5d50911f12", x"d83604ebaa3e5383", x"4fff2f208bbd08eb", x"671773be8d69cfac");
            when 29738230 => data <= (x"d417b64e7bb6b1e8", x"70561784699c0bf5", x"5551cace207cc8b6", x"7c7ad7f37c9086fd", x"f34dbdb0caeee24b", x"c6f8922cd57979f9", x"cdf978bbcc983ada", x"f812cb1a5e755747");
            when 18369805 => data <= (x"da4534bf97675da7", x"392f4229456976f7", x"806f650a8ab8a1fa", x"09ad63508c6aac3d", x"36ab634817c69005", x"138fe0bd4001c4a6", x"b2a581b76da2c906", x"a498743bcd888432");
            when 23485497 => data <= (x"677761cb3f9ef2eb", x"1a0efe4426c9a26a", x"dc4987788dba80c8", x"aa707c5427c4f45e", x"159db6241addd50d", x"d621110c6f5d577e", x"953b1f9c66de24ad", x"a6e369cdbd2fe9f4");
            when 16824361 => data <= (x"16b99a259ab64385", x"5ce08519f244c260", x"40e1825fbf12e460", x"9f0172a2f39f4a06", x"9ec5f634189ed3a8", x"8bb41c7cc1412f4f", x"8e05ea89bc324152", x"d84d4ec9973e34e2");
            when 20728915 => data <= (x"2c3b9abc4effd812", x"56f4f27d623b73de", x"b3cfc035ee7c7c5d", x"8b5cdd3378af8cae", x"2852c95cac56f477", x"b1119802879a1e46", x"6cf8f3516ee4d036", x"5c5032910811b4cb");
            when 5694603 => data <= (x"0dc18d97318e4ce6", x"2803d26bce30c7e2", x"6a664447c9aca059", x"0578d7b77515a143", x"225cbcd14eb96a3a", x"fc5c5f7f29f63d79", x"9334928f40d98924", x"0b080dd739e21d21");
            when 9169419 => data <= (x"ca6f2880c4a8c830", x"31c3578b54638a3b", x"a7931e49fef4e321", x"b8a3b1987420fdf6", x"db4fbc5d40980af8", x"6b9c760b0632a1b3", x"71f0b27b960c71fe", x"bf518111965436bd");
            when 15777953 => data <= (x"bb4c266de15d923d", x"a1cbcb0ed0fbfa80", x"8a909717a61ccb9b", x"fcee1bc309136999", x"248a7c7ba9236217", x"9a1a6611844628dc", x"9a6d61e7c407315e", x"635aace6fae25310");
            when 10565033 => data <= (x"1de603308c782fb1", x"a8921b86553e112f", x"ac80586ce0be1725", x"a1585fa1550382ca", x"59351d1e977f5064", x"e89b128557b09b7d", x"3cdf3ebe1f701e5a", x"d25886dd1ebcfa8e");
            when 17236897 => data <= (x"475a00bb9f3fadb2", x"d7121638f48736f8", x"2f883611a3a3a1b8", x"d7ea2c055e141e9f", x"a5a71b0ebeb34b6f", x"2569c00b13d441a3", x"a51bc5f0f50f591f", x"b67802b1ab57e31c");
            when 33192148 => data <= (x"4cd4c7423461480a", x"00edbbb21c4c8585", x"58bf53364a5e81a3", x"5aa79786dc950629", x"d0d83e629533a0b7", x"882c8cfeabf4a4a7", x"bd3d9f4d0d2186cd", x"aac72a5339236f3a");
            when 33321489 => data <= (x"af1121301edce668", x"786ed7a32a92f08d", x"0fef2860538c0630", x"d671e7e79cb1c4e5", x"f32a1a73d10db042", x"296c6715e9189abd", x"b1a0af70d92dabbc", x"0118a740855090dd");
            when 15551947 => data <= (x"b072f389a33f344a", x"a018fad2afdccbed", x"78224b218613ccb8", x"616074c3e0c18da0", x"a2e831e446ee456e", x"471fcc936bb94a57", x"1bf77aac8fe9c2d8", x"e06c8b611dbd1d27");
            when 20724410 => data <= (x"f2ed696481bc8d21", x"b0f47eab929bf3a9", x"9ceed17aa67bcf55", x"499f6d0c710463fd", x"9c604414dc67ca13", x"60f9ee4233e6c3a9", x"08986e81606f0825", x"9a296d5306dd398a");
            when 10840194 => data <= (x"4bac333d2b348392", x"e79d76cae41d3463", x"f296abf496ed6b61", x"9ac83a105878ca18", x"22705b4f88cac5a1", x"a364b854f49bc103", x"a8d1b371269d6c4e", x"aefd63b744b17521");
            when 1534452 => data <= (x"bd6c0fd3c8e4fa11", x"39befb374aaf561d", x"e14226426f8d9ad8", x"df2157b09df159af", x"13510600a9298659", x"273afdfde9b46032", x"17b1ca73cf8a9936", x"5d13fc7dda9038b7");
            when 28570463 => data <= (x"d834606b0b7da7d8", x"862bc566aef072ef", x"d5cb8cfdf87a6995", x"f19583c3598ae87e", x"6960a627805bf845", x"31c14d096a946331", x"6152f30ae7b20592", x"1de8596d434fbe28");
            when 16583474 => data <= (x"bb348da484575370", x"d61d2c6e8659d46e", x"3af38311b30aeec4", x"2a887808da6c0249", x"d5c02097e3939dfb", x"64f6468e5611993d", x"5cb232a52bec390e", x"ffab1a9717c9186b");
            when 32903080 => data <= (x"14ca7191769d5f93", x"39c49b1656d12ada", x"2aebc50fbcaaa352", x"0acc73343b5228de", x"a8083eb9af94f7da", x"993c754aa2b2f948", x"af0c6e0c3807953e", x"dfd474a03cec1763");
            when 9463035 => data <= (x"38d67787061f4d2d", x"531e08dd7da1464b", x"93a091a648255782", x"38993638dda041c7", x"30771fc65d9b4745", x"a10951778617287b", x"cd1a8f63a5ee1c4b", x"bf6afa8cdb8eec93");
            when 14577397 => data <= (x"2c9370ea70eda50a", x"b2787d2437a5099b", x"fec90c1983e9964f", x"e3e1fcbcc3743fd0", x"f5f4f4056e2098d7", x"4f9be0f5dc8a9fc4", x"5afe4cbd3f86da3f", x"7b3f53682eea6069");
            when 4396542 => data <= (x"f06ef36d67508e2a", x"6cd904312ce9d379", x"dd09c7da2513f962", x"9cab4a96df70c792", x"af1c1e6e757d039d", x"243d9cb0536cb933", x"e6ae320ddfcf92f2", x"d3022dcf4216f8dd");
            when 17572337 => data <= (x"eae746adfaa816b8", x"179d03dfef54976f", x"a5375e2700c57e0d", x"db1b8bbd69ae25f4", x"cc1353d97b205033", x"f88675eabe55d373", x"3431ddc50ed7114e", x"e33be8260f9b1910");
            when 7103074 => data <= (x"39980378f8720cf8", x"aae9e0e1253207da", x"1bee3294537225a4", x"b121f9bc87a19444", x"a8095cb4ecf235ad", x"a9b62bffebe90981", x"21c4019d2a198076", x"6c50a6856c607db4");
            when 13988960 => data <= (x"3d6b730324272ae0", x"bbf8c6a15cb78afc", x"e036e3c29b18fc70", x"796378fe28496edf", x"8966bd14c12fba2d", x"efbeb6f2b37c5414", x"f9514589c579e9f2", x"ffa4f7cc3d8a4b8c");
            when 7580225 => data <= (x"0b4b29cb8c13a3b5", x"a492ce36ff17ffde", x"1b0d6ed9e2fec490", x"0ce719d690738144", x"fa69f701dc10babc", x"ac54aa6cf398dfda", x"828ada4560e4e907", x"736a148d254f56db");
            when 20808630 => data <= (x"0a8c28888493cb0a", x"eaebbe80fab9e589", x"e4cc58b31410e2aa", x"331dfc5fb18ee03a", x"1ef131a8ce1b86ea", x"2d18474de061bb37", x"86432c7619cad962", x"14ba565c53693ec5");
            when 16411589 => data <= (x"263740627470c903", x"ff63c3bb949e82dd", x"2fceb194c73d11cf", x"0121ebdb058ef8c1", x"b1e73ce355ff8455", x"3ec922503540f5bc", x"5fa4e2d3b73a51ec", x"32fd424db3a7e4f5");
            when 11259118 => data <= (x"08e85b22366c9b5c", x"37af96e955579ab1", x"5d91c32174d6fab2", x"5d162d16b06ce2bc", x"dc1810b4672e9020", x"5de97c17e84e0d0e", x"cfa78d09fee20a13", x"3018e2cf3b3b9316");
            when 22299297 => data <= (x"766b4e13182f7f41", x"d10066fe0c6af381", x"aa80b7c0d84ef699", x"62bc78f32c8c77dc", x"f7907044e0cea0b3", x"99a58a4f48a168ff", x"b03d709d69842198", x"26dbb79f521fdbe5");
            when 29361526 => data <= (x"2593b6a67b0ee796", x"3aa9aeca1c9d6476", x"607c588917d0c6d8", x"c186c7df4849b95f", x"dc2ad30539177671", x"11968e384c139cb5", x"90712b6f92fdf58b", x"ebe5e817fd093b9f");
            when 28115419 => data <= (x"cd0bf8564b2f1e84", x"d91a2c8d7042a246", x"682343464b4338b3", x"fa997d908a737bcc", x"47b568ccae277a01", x"c3574efa2676dd0b", x"449abcda96dd8411", x"cc6bdb4ac825db45");
            when 4676359 => data <= (x"ded9318b2828c686", x"a3c3138ced52bac7", x"408be27ec46ef122", x"efe012b586b46efd", x"a9207ab81d199129", x"eb997e949c3c8334", x"dcfe8e94c0c93b97", x"256430ca8aa0aa70");
            when 17786930 => data <= (x"ecb90c6092265760", x"8440407161fabe16", x"436df97cc7f90ea0", x"08dba3505cd0de3c", x"8c6b5b3b60302156", x"c61b89badb07e37e", x"1e0a6ad99f63c219", x"cc3a5456fdeb8627");
            when 32764826 => data <= (x"ec791adaab2794b7", x"5611e7e9fd964fe5", x"5e93e596e42a4465", x"026b6e4b22a287f0", x"9e36447d8662ee69", x"730263616c610cf4", x"6234720d17d495c6", x"d7face55ee27e8be");
            when 32192645 => data <= (x"5119a6773a4c84ef", x"771004923b16c048", x"d46730cb4033d710", x"4c5fa13fdda8e5db", x"d12eeab72d84cef6", x"76f271d5c5652ba4", x"68cd571d31648c9c", x"c886f0887e9d6154");
            when 26401124 => data <= (x"26036001b265f208", x"7afb17c559cbc580", x"cd285f059efb4d1f", x"14485a5084f27306", x"8953b22777a9fe50", x"4eb20df0d815b55c", x"d6b18e4f17038c6c", x"21a042ab85e6560b");
            when 15809692 => data <= (x"218481ebd7e31e2a", x"34c8f6b9f3e01f1b", x"c2d6b0387c12e97c", x"5539c0504c26e24c", x"e3786b98a5c758e7", x"1b65ac9087a27cb0", x"2c9e55d9b155e1ac", x"3301177f61bc9c83");
            when 32425413 => data <= (x"9e2e03f1186daf3a", x"6f4ea9855f01423b", x"45d81fe226f12b43", x"bbb3518f58a953d7", x"7b6d740e0c02b9e4", x"72c98532e1942ab6", x"de1d244d75a8ae32", x"801e7776ccd390af");
            when 14439302 => data <= (x"a790e46aa4c80efe", x"e7bb6a097fe6f490", x"e7d95fe7f72f8b47", x"b5f8bd67d8e2feda", x"4a2ab4a4d3007e31", x"129127040dc53fd7", x"4fa494f9670b091d", x"28d373f9250c4e04");
            when 11676627 => data <= (x"281c082e4532c746", x"bbc7a9f52680d187", x"b3254f67358ac8b0", x"35df4295ea836d1b", x"657ab081cccfa58d", x"d6f1e575978b4cbf", x"95e5fae56d105a25", x"1a26589d5bb4cebd");
            when 24209007 => data <= (x"7cfb8b07b85b1988", x"7ae036e3c7732d0e", x"468e4bd1f47bd413", x"b78b1bc45342ade4", x"f9560ca38da2ef65", x"2f653643b03c5ba8", x"714cadf921c3ee18", x"f6b837b1de0a2be2");
            when 17826120 => data <= (x"c255fa2a53449320", x"fcfb8f547be30a3c", x"0204813cee130c4d", x"3d374ff24031411a", x"7bc2a56d63dd84f4", x"a00650d4f1d75ef0", x"4248ffc8776824a4", x"ef4fb167db7d1599");
            when 13612857 => data <= (x"d0ca718b60c60356", x"8f5e1263f4dd8de1", x"0af0499e8ac254be", x"0e797d4f9e92612e", x"c0894ae303bc79f1", x"40a2cfc477203f82", x"139acd3464c6be46", x"8f79b7fc15544136");
            when 20354027 => data <= (x"1b2b83a6848f707a", x"c867336a3df395d0", x"bf1953c7735c39ca", x"2a5ab05061bb14e9", x"319366929310d711", x"8a753631d10465f0", x"c719d3bbfab90c3b", x"4dc3a8b2a4af9abf");
            when 32556724 => data <= (x"430efaa6e378ee3f", x"9e0065545e708dd6", x"7d20977c3ae206e2", x"02f5d2833d785516", x"9414562dcdc841ce", x"e9c03308a969848f", x"3d7296be952e4313", x"79f4bb75fd9b9c81");
            when 2112925 => data <= (x"858fbb9f2370ea62", x"f6b81bb183321f77", x"9f371b0f1ebc12d2", x"9e5a391c4a7248ea", x"b1a3fafe9e050cef", x"5a91d15a8dd1ba00", x"c65bec4b78368c43", x"8f9eb25d00b65eb9");
            when 1397537 => data <= (x"ebe9d5ede2f58394", x"fef79b28d6994708", x"b9f8a389ebc4bd1a", x"b27c3f1e93762540", x"3395938c16ccf527", x"6b66574dcb18d147", x"334eb52ca1451f65", x"9ff0244b29a91e66");
            when 23223104 => data <= (x"311cc1795f0b7d13", x"a65b96bab109d768", x"c13aa5f27893316b", x"75f65dd8b1c17bff", x"1f85681b87cf0233", x"c4e47919e48ca7da", x"6de8e3fb6d31073b", x"a7d4e6732a0a7834");
            when 17266290 => data <= (x"caed7545ea2398fc", x"ea21f8d8814dfaee", x"93f4b59d8838d8b8", x"d8ccd37c497becde", x"c139b760f7ef0f1b", x"150e6e75285c01ab", x"89ac9f0c80f64ffe", x"d319ed198c436a06");
            when 18410367 => data <= (x"2fade02401057b18", x"5b333c7c1cf3d356", x"8cc0543caf4c2517", x"662121ba3f194bd5", x"90cfa964996f1cf7", x"27b14d1eca56267d", x"70331146dfcf8995", x"d126b44fcea89996");
            when 32997050 => data <= (x"325c5042f2062658", x"ce5394b0e448863e", x"e2e029a430cb3d07", x"0406ceb4225d53c2", x"ae2431c466092820", x"413416ce9a8cf3c2", x"0429142c1bf8de3c", x"0706b4919830600a");
            when 32104876 => data <= (x"08a8ba6efc021583", x"6e59851421c43d2c", x"ee5a3891611cbca4", x"363092c13926f9d9", x"0a48f8af01e90def", x"cfd56c564f562f3b", x"cec2b71ed3694160", x"a04768b5b7b35b7f");
            when 5437957 => data <= (x"86ab5a617a9a8443", x"d42f434b197c95fb", x"4415b54bdf0d96aa", x"2425294a30c609d5", x"2c3fd18eed836eae", x"cb3f65407301f1d3", x"2d2eb1bc4f6f94a5", x"4bd296d01e61c576");
            when 32480678 => data <= (x"8b7d712f67d5f2d4", x"6103a60fdf63ab05", x"d4c4f314feaea0cb", x"76c4465358f7a54f", x"0d918192c1d10a4d", x"3e86ea6e47793561", x"7f12478d00862f3a", x"6eaf269e23866532");
            when 16388091 => data <= (x"2678a747e73770af", x"326996f1c2394c9f", x"149a4fec7e559dc1", x"21e56c547762ea8d", x"03aa54b8d8102bbe", x"507bd4ae1668458a", x"c8933591cb07750d", x"e7744aca58cd11d0");
            when 11742095 => data <= (x"611dab0868709a8f", x"7df329adfcecdac0", x"04f0f80f7903c340", x"3a55aec817906833", x"19d1cf39578582cf", x"85327910b4fd15f3", x"418c6140c2fc6d3b", x"a7074e0f6b2cdf54");
            when 9124347 => data <= (x"cba513cc949c8997", x"ec30a75cc8b8bc38", x"8cb57e172a258a28", x"9c5114a4e2b2b5c9", x"91e45c55546637a1", x"cf8d3ffbea41b459", x"20c2c40c2ce94ea0", x"6ae7fb38330162f1");
            when 11176966 => data <= (x"59f0b3a87290cfb0", x"370dff972aec9af7", x"8ea63c32c350b641", x"53401e5fb046fe75", x"647dbcc04b482ef3", x"9d53eee2cf696260", x"e5c14f8a418fb469", x"22652379352be283");
            when 25435577 => data <= (x"a89e465e7f806533", x"4054e559774dfaef", x"17fc606907317284", x"e46562a52d24627b", x"649dc992fe3ea48d", x"3846691dbd59f616", x"a4a67cca61450ef3", x"32231d600c3a1a63");
            when 21653000 => data <= (x"f98f31b2f5cb8bc3", x"64198105d2e17055", x"a7f3b7009bf72c4f", x"1bbad38469ac12c8", x"8cac3d8f5130e4db", x"3960cd07de0388a3", x"1675b6e4026fb9b7", x"7e605e19dfe5f71d");
            when 2803502 => data <= (x"e938ba968cd273ab", x"d775c20c22c2f7b1", x"c8fa06d7d55a4e1b", x"3079e56d641c680a", x"1edab5e4c493fb6f", x"8c248a842a22824f", x"d4262a69d8aa08a0", x"525ce3632763e7cb");
            when 21973317 => data <= (x"67f0ba5b61d7986d", x"1ba43a3fe82ef648", x"9e6fa4076c9e7024", x"1528da77b2ece8ee", x"73ee753a561d081d", x"f7bcfbaf4e5531ff", x"6f64fa7029808b6b", x"e0169b003f560326");
            when 16543637 => data <= (x"7883fbf2483bdbed", x"1f8ae26645dc65f1", x"b1c47f9b2bbeafbd", x"5a596b397288f90f", x"e02680d378f0090f", x"fa5b8926c17de729", x"a72a120e660c5c10", x"232eb4f6a5fa9e6a");
            when 24574012 => data <= (x"890e8a6a60a6fed3", x"e45049d4da7c08fe", x"ca7a084204a7d9a9", x"ca665ccff03cb8a4", x"1af6e5f45906e080", x"81389eb7f4f51da2", x"73b37208118311c0", x"11b874c23a065803");
            when 11938406 => data <= (x"5e88aa2043a29804", x"77707325070cf5d8", x"5ac880ddd5f13218", x"b0a3d91276d23419", x"c041aa38beb4a0e2", x"c53dd90488c4f924", x"ba6e85cf4f3964db", x"892cc75e4bcd7ae1");
            when 31245133 => data <= (x"8f9bac17ac6cfa4b", x"f557d488c99d8e21", x"28cb6676da49b49c", x"f6c405c527d8dcbd", x"8c98de4ced5bacbe", x"50b32c610d218c58", x"db628fa15fc795ba", x"3ce5808977a611d9");
            when 10458376 => data <= (x"e8a9ee0fee043795", x"9e7d0b732ee09c87", x"7c2b1f8d031ad393", x"700558acba31a303", x"09c273bdfc935f96", x"4ca90d6450662b5d", x"9424a62e49378313", x"849c21f22d6a3e75");
            when 15281208 => data <= (x"94afcbdb9501dffa", x"54e2356a3d22d2e8", x"4aa5b1e8548c3d0a", x"352e8ac29e7db499", x"e3b1fb2275adde0b", x"91730fde7670a680", x"8990bbf053c7c879", x"3a2413e1ea8ac3d1");
            when 26957377 => data <= (x"df5bf9f129b5c99d", x"2ad6805271591304", x"c26e518758dbd6c5", x"b309f8fc425a0214", x"b5177bd80850ffa9", x"f5f0e944f05c0144", x"73024cbe72aa0a03", x"80a3f36328bf0874");
            when 12827997 => data <= (x"3c460da4b658cd7a", x"91c65f26fb04714c", x"2caceb506f40bfa2", x"630b25be3a54177c", x"ba6cd76f8ae5caad", x"9906b5137bab10b5", x"296d6cf9e0d76a1d", x"3fdec3b529a47040");
            when 16862873 => data <= (x"f9256fdac642463a", x"7444304104c0bf38", x"3328fb8ce931ccf2", x"ee1e825f16fa7f30", x"49f95c4ecac71d13", x"57ba86510fa60005", x"1cf018fa66694cbe", x"23b1530da9706f71");
            when 1493377 => data <= (x"26f10e73b10ca923", x"1e365c82ac86687c", x"72047a159f421e43", x"db8b67d1f3b83cc2", x"d5ee80329edefb8e", x"4f9693945d90a2fb", x"bdedffd244d8677c", x"b9c3259b8127b578");
            when 30868225 => data <= (x"e0bb64694cce06da", x"7dc8cb558338cac3", x"9484ea39c1dea04d", x"0a2ff8d611d384a2", x"c28223ae2667fa91", x"1bc0a4d800e91b85", x"dd34835032fc7ca3", x"935adee1abad3ac9");
            when 32387449 => data <= (x"22d4460d9d560597", x"6ccdb6777937087f", x"33637318cb95a77a", x"e30e1c7df548b328", x"145a002ae0b2b623", x"ea4a6f1b1f994f3f", x"da1afbd97d9860ab", x"a11564056df0f29e");
            when 15405853 => data <= (x"81acc101036ceedb", x"20cddafd2ba5d34b", x"dbe239d9dfb7f507", x"9461a1702f230ebf", x"b8d411ae8f2d7c24", x"a80e9507f7fa343e", x"c25aa0e02aaafa55", x"a491817ef76b0db6");
            when 14382288 => data <= (x"78288796c4f47f4b", x"94852617115e5c56", x"512b5114746a5fed", x"638db5643e438c5d", x"c4e195e95986f76a", x"41118fd1562a3866", x"1ac4133986c461b4", x"6529659b2ec0c2e4");
            when 22279087 => data <= (x"9aaff073ebc1561a", x"8026e963ab62ab05", x"98f4f63d7a90d89f", x"6750a749239a006c", x"192796a6cbb8a167", x"54eddebab5f57a57", x"55314d54c6ef528e", x"c5f3d47b3914abf0");
            when 4376285 => data <= (x"f4faff03b4622ce8", x"dcfe697f9d2867da", x"0e0c2fdaa2f5d396", x"9c411bcef7719d6f", x"939fd7721b9dc896", x"b894758c05639650", x"46ebb58cea272f43", x"0a8637ac95524e26");
            when 3337125 => data <= (x"b2fcff39c1dff5d2", x"8b86c3e81a999620", x"fad21aadf2ba22e3", x"69f5d6b0723cdd50", x"3242538bfdf95c6d", x"79ccaacd914d4e49", x"04098fe1bc704880", x"493c285ae0b9ce30");
            when 8809639 => data <= (x"9f31f5e4542c160c", x"6cfd7d49096921d6", x"6420c64b1a119ad1", x"c0bee82f32176f30", x"5bff152ad223682c", x"af8dd6eb9d3dcb35", x"f913702a897c9a11", x"94f31ec7a524099a");
            when 20603166 => data <= (x"d4b75babd08480b0", x"5ae3d68c2b2e7b85", x"e1b564fa269cc8a7", x"06c10879fc925216", x"9b75c75c8e352524", x"e53f22b930eba503", x"ccc01be3e0123a26", x"fbf1e825482ee5a6");
            when 1010273 => data <= (x"2e0fb83a0ee992f4", x"142d72f8dd4167fe", x"d46a8b43aecaa08e", x"ad10d0e13311bc6b", x"a8d3c079d6abdc55", x"dbd97b89524d19bd", x"69701200326e7f87", x"3f57571fa00b1b06");
            when 19267395 => data <= (x"8d42a2bd89620440", x"102549040debde37", x"87598b7ca1803080", x"f6d2961a2a7cf305", x"91641acebf1f4faa", x"58644b18c035a62b", x"0f9f9e42595021f7", x"04dc5cd366944e29");
            when 5787644 => data <= (x"d3eda7ac3e449db6", x"b238dbd7b5aee198", x"d44c594fab297a41", x"9ac07c52251cc51e", x"4cf4863578bfc7fb", x"4bcd875fd554f4d8", x"cfcd78c309efb0fe", x"5dba2d64a815b8de");
            when 7341343 => data <= (x"f795d380be4e2f9d", x"9e3a60a1065579dd", x"0e41c4a1487dfe46", x"8d196ef5b3e66db6", x"7a8ace0ef2fb075d", x"9b77f51fa66ae37e", x"6c46656964573254", x"09191bda06949474");
            when 11677660 => data <= (x"517451637f3279a2", x"6e8b24c21d04c982", x"d844cfdcb4fb458d", x"2872565c4e46f7b1", x"770436d6ba4c6f2c", x"4a58437645ee89e1", x"08895843bc7a72b4", x"4e0064c51787f43f");
            when 25316534 => data <= (x"b65a4e85227bd8ea", x"cb01e6d81ad42cc6", x"c7d172b559ad907b", x"26cbf2a5c10cac36", x"398276319f114be2", x"b6c10f22b43dc184", x"5d0609255f090dcf", x"02b72474aa8980e5");
            when 5296912 => data <= (x"b103101372894da7", x"4672b2c4dcd25d36", x"146df3b0997c4dbe", x"75d2026faabea92b", x"143238c62c366cb5", x"4ae6f0df512923fc", x"5ee4d5e80337fab5", x"7b6b0e210ecb8e0a");
            when 28846495 => data <= (x"ed39f90e69c24ff3", x"7612365436228363", x"b451833cd15370ca", x"9449781e99eb548e", x"46164fdd84bb4d7e", x"ca0d017ba06bb010", x"6712a55faebcdda4", x"e54a8d0cf9991116");
            when 21731810 => data <= (x"daf1fad5a3d593af", x"f0d101cbf8eb3142", x"870539fb6bf5092e", x"45973ef191acf2e7", x"61a3e88371d775df", x"b61679964d73824a", x"ce15e994197245cc", x"385a8e2a059e778f");
            when 12885601 => data <= (x"4358d6736d907cb3", x"be9d8e55f3217c4c", x"bed70a128265ef3d", x"4bd0dc7310426d07", x"c695ca51d6e14ac9", x"a37045af49e0ff0d", x"a045c3ea7018ec54", x"2932fe7fa2789983");
            when 31165181 => data <= (x"7df32e035b57af4b", x"7538717c53e803eb", x"29f52d27664fbc11", x"691f935463e92b6f", x"e366c551b8488e41", x"4844d6eb135b53c6", x"9d719f4d251f249e", x"3b260e6d2db40e46");
            when 1794630 => data <= (x"19cdbe8cbad35c35", x"d88431e1aade1810", x"b0db9e2071ceec76", x"59c4db9147660a21", x"fa7ad995983f460f", x"78949fa419178e9b", x"b9abb100ad5ab729", x"5de46c99a764af27");
            when 13261749 => data <= (x"010da1462150ffe3", x"e0da9e843c9bb687", x"34689ba263f6f280", x"2bd06a3c6627a479", x"ff25e73b8cbe9d93", x"82c795749f46d6bc", x"bc21e654e51c537e", x"8a603678da84cb5d");
            when 13226931 => data <= (x"a7d5fed118ae3fb1", x"2c55f14757c9b07c", x"3b8c66c08a47e3a9", x"5b0d6ae1d410399c", x"0b37f9108ad87ee5", x"36721d361e8929da", x"beb1a7dd6624fc95", x"3374b8e6368b283e");
            when 18953838 => data <= (x"51b2c880fc23e43b", x"a9a4db9eb82928a0", x"a8b9250329daa113", x"da4fd44e542d00d3", x"8075ed86890663e1", x"381ff13495fd9286", x"cfad2d8bd3f898d5", x"4a19c028e442a27b");
            when 18651503 => data <= (x"19fe8520cf3f8c96", x"ec085b4b3be64f73", x"836294099753d01d", x"d61bafc083d86e27", x"b8c5b663bd1564f0", x"214a0bb0186ee858", x"768846ad177b7ea0", x"f2fdd5963de65e08");
            when 1508053 => data <= (x"cc645145a17fddde", x"a836990fa0ee7152", x"f0e43234d4c71174", x"a46dad68cfaec167", x"f44cb3196497c70e", x"b73c942fc638cfab", x"841190e9c721e0ee", x"5e00fe61519d3ab3");
            when 23064030 => data <= (x"2aa05cc25da59bcc", x"968a0cb023b91893", x"1fbfc80f04d81fd3", x"d437bf9c76fa9e11", x"609d3a92c86571aa", x"30c175edbb937ae2", x"320633c14d1743dc", x"8db19fc19f81047a");
            when 15723994 => data <= (x"7d22f4139d8a781e", x"03121aa220d38482", x"7bca2bed8c598cb8", x"a3be9e354c2d933e", x"5aaf5e04b4d56be2", x"629044e56f7b58e0", x"e3b5a8139195a6ce", x"6517d0c33fb78c96");
            when 14599417 => data <= (x"e828cc999f3c794c", x"d3d5ec6ad84e645f", x"aaf20aa90a0e2f1c", x"2feacc822cbc6252", x"114466d0c64024c8", x"b596725275924cb1", x"32eb4c0c5abd522b", x"92be72c7653e7f6c");
            when 31047279 => data <= (x"80ccca079eb878c8", x"e1574dd59435ea22", x"358b5cadca261c5b", x"fe3ac91870d1fe67", x"1a31fa1788f90ace", x"aa7456b7b52ee23d", x"799d58a4e321f72e", x"3f961556121d6e34");
            when 610856 => data <= (x"65f96de93ffe6929", x"da54bddcf39a23fe", x"a63952077d984358", x"6717d293d3951914", x"f6441fc7ae43fa4e", x"c494df04a5588a13", x"19453f86233ca7fd", x"72ba6145d6fee378");
            when 32656445 => data <= (x"fec90c2d21ff6a14", x"6a48659c663cdfd2", x"88c7dd014c9ef85f", x"2d9fcaa08bfa8387", x"69e28417b3ac00bb", x"a15e0befe43e0a8b", x"540a5073dc7f87ce", x"52303c904ced7973");
            when 1268312 => data <= (x"42c0b5214f9c995e", x"74bec2e4d90d67ad", x"18b387f4906b7098", x"66393e11256f43be", x"94436635c93a5a71", x"7adda2da791d8fc1", x"f20fa5025d302255", x"a1802d2c20fdeaa0");
            when 27519422 => data <= (x"7f9fae46117bbb2f", x"b5c7f4e6be94939d", x"942af464071dbdf7", x"c3e8891e424c4937", x"5abce488365ba9b4", x"63ab46f001a2ad18", x"acb4eba0869b0b88", x"2c2d58bc1397af53");
            when 32762356 => data <= (x"51f1516de8e1a7d9", x"0ba4a2adfe6ace45", x"6a8616d3484adf71", x"835af4dd10dd571f", x"2b595507fca2d097", x"b573110cfec0a2e9", x"23aad57e1a98c1d1", x"997d3bf84b4a1708");
            when 29621992 => data <= (x"4bef321e4f2d3dc9", x"3e905f97a2e4b070", x"75d05fe8839f6c0e", x"374c770a3482c14b", x"c9a6ead780952d58", x"609a7230f987c5e2", x"519c3df208e02c4e", x"7c8faf87813a2509");
            when 15038909 => data <= (x"0e8cc775f743d9bb", x"4072644070f3c3eb", x"7297cb8e42e41651", x"685c74651c36dd1d", x"9a65d1b28c1e92d5", x"7acfba2a2bd8a1ca", x"1954a39ac2348998", x"cd09c93229bec48c");
            when 13365315 => data <= (x"a8f413dcbd056698", x"d0ad91a48ef34d00", x"3d560fa9d15c0bdb", x"59eecd4611bbba19", x"2ca682df59c57476", x"13322b56b0b1dcce", x"8b505425590143eb", x"8f6d8e9ef213a321");
            when 16842521 => data <= (x"30c95ddbcd67acd6", x"7463b2a8e2c16eeb", x"f8ee1325a6902724", x"88372ff6d390d3b3", x"bd53c4d6248602e8", x"ea71856ad27a39dd", x"7739355011fec86b", x"295f8557dcd75e19");
            when 11351587 => data <= (x"42564d4bcfc8f3b4", x"e8549330e8b95b94", x"12a6ead7dae5086b", x"22bf242f66c75368", x"6d6a801fff263018", x"e8f81e2da068dddd", x"91ded8c5d340f206", x"bfe05595628f32f9");
            when 5718034 => data <= (x"8c2a8dc5d8f32ca2", x"9ce8cc70682c3fec", x"e1a86a89f1fcb6b5", x"2c56ef3a16aea782", x"3656779d89a5b593", x"f056adbc745bd728", x"f6c3f40ca93de43b", x"2d9fa6cff4b0e442");
            when 30268457 => data <= (x"da7b2b0c3dbb0809", x"d97c5f87ca7d0a18", x"4ae9d088fcd61189", x"267a3ac6b985704b", x"ce53873d5c0a7109", x"c14c5541e670eed2", x"8605c04bec3934d8", x"81bc47c258744cb1");
            when 23185522 => data <= (x"88da0746b1f86c34", x"fb5c8a94f921fbe6", x"1557714be69a1ecf", x"2dda7ee4f857d823", x"50cc30bc664926ef", x"a71ae470076140f4", x"4047264990f9b842", x"37f56a7b69c70e5a");
            when 15457337 => data <= (x"7d4275233576fd12", x"3381516a70feab3c", x"f10ed7fc999ec766", x"3ab2d083db1e106e", x"898d6afcaf8d24e6", x"e4caf113e38815c0", x"642c17b050d03083", x"2216ef62be65e380");
            when 1051563 => data <= (x"bd0498b27f039455", x"b3a147558129e1c0", x"a6ca66aaaa4d6bda", x"c916831c990ef12f", x"a12845c23158c727", x"584aaa5b06cb3ee6", x"0e16014150062266", x"96a3b9439065087e");
            when 16418944 => data <= (x"4019d00fa3bdd1a0", x"1548b1e0bcac0ead", x"bf8c7733c5efffc2", x"2fe6fc63fe50b43c", x"990e8585d431141e", x"9027ac60a71cb233", x"ddf65a9051407385", x"86e2017383814f17");
            when 33147108 => data <= (x"7c16d34c44a615fa", x"c3e8b4330347f306", x"0e9ce5661d98a289", x"871462fe4bfbdd01", x"03293b5e5c96d78d", x"8f2fee43e0486d43", x"afe0d854344e6a4b", x"04ef70a5ada9a6fa");
            when 26867537 => data <= (x"c9b82a6ed66ac071", x"54d27a6f514b4013", x"94432f2d57809769", x"01737a5ec1c817a7", x"07d3ae639d9db953", x"a8a30934491ac951", x"80cfa47c37828731", x"95fa00533e389ecf");
            when 29274912 => data <= (x"3c245215fdd38ef3", x"a0c91f4853818687", x"4d89a18722b3a24b", x"81e63f81528626b2", x"019191ebdd92f8ff", x"2724a4fe05c1bfb6", x"9d05e897a76265c1", x"1108ff5a33484c25");
            when 17899582 => data <= (x"e6a07cfa24f88ede", x"20e1710fb90b00ca", x"c5943f2a11a134b4", x"6deae3c26daf8b5e", x"475607bad70d1753", x"731fdc2b3348e62d", x"87230d68043a445e", x"5fa8b6031fdaf5c1");
            when 15674257 => data <= (x"4258c3b2bfd7f69f", x"83a38086d1cf255e", x"4f197a109830312a", x"ad403e0dc715ce2b", x"386ddf4f2d230f0f", x"92f5dddd7921c437", x"065a831d70d60dfb", x"6d26cdbe2913239e");
            when 25764049 => data <= (x"2277405071c27e9d", x"e90281348c722632", x"c5ac72c34535d35e", x"a9e92edfddc115aa", x"07d854c78bb57ba9", x"d3adcb1aa8b4e8ef", x"7f11c6b3eee439e1", x"8ffc2f662e014a07");
            when 29511106 => data <= (x"1633442b24a11cdb", x"f23f1f70cee3bdc1", x"938a272f62614d41", x"eafc308e407afd60", x"4665ae4ac0661c40", x"6b85896c753ba62e", x"ae18ee531810886b", x"d4568f8055bb1a7d");
            when 5444778 => data <= (x"71c4042e857b9260", x"6951775232fcf892", x"a20ab8233fdc5eea", x"e3354ba55afb4c6f", x"23da969db6f816d2", x"324ce8bdf06bbf85", x"daef4c455c4a58e8", x"eae2b2b70e0eb080");
            when 16017227 => data <= (x"a3bc5fec7c9fa8fe", x"d4703ed451a1162b", x"a7b8232ac6cbb57b", x"3e2aa4b3ec5bb5f7", x"d73c5c41f171475c", x"8ec264a46ce7148e", x"3ef6a90f102b6e5b", x"9abb0ba2ca2530a0");
            when 16162214 => data <= (x"f5472e21e8817037", x"b97d502ea88ae980", x"a0ff8e7b7902260a", x"771229430f2a5bb0", x"56e31694be23b36c", x"d62c28a8aa96c4cb", x"87e6678d69cf6145", x"963cf9a736be840b");
            when 32769463 => data <= (x"80638a61debdeb33", x"9afc40dae80b8754", x"722742e58e30191a", x"bbbaada889fdc0d0", x"eec0bc59e06bba5b", x"87147d987a5733b2", x"d857562f73455c40", x"72eeaf7582ee81d7");
            when 23615335 => data <= (x"56a84f8ba94b8f4d", x"6b50f1881a4411a3", x"3c6cc5779c1f3317", x"3f3063f5764fb1ea", x"02880b4f8677c844", x"e733d37c0c36a917", x"76779b18a4990df2", x"36ea07a2e7510801");
            when 27165684 => data <= (x"ab56cf58c182c2eb", x"7ddb99ca9caafb33", x"c437167a3b65ee17", x"4ce4a97c3a15a26f", x"f3c9ff5c22c9a123", x"9df63e3b1da6aee0", x"fa83bd8e140a9548", x"5ad086e64977162e");
            when 11148039 => data <= (x"89e59edb9dad184d", x"45f4923a23378e0a", x"23c5f9ee8c4becb4", x"a699df87d7d04b35", x"eae5e54ab888e9db", x"5f098601b7e5d84d", x"ab155e4d922a70c0", x"3433d69668563824");
            when 1582708 => data <= (x"4b3889d0bd60ddd7", x"3b9f47b17e7a4a51", x"e6a4eb74235a7c04", x"6dfd3f2e4d3a8c3b", x"2e4308a54906b2e3", x"0c2c433daed251f7", x"ae645b41f407961e", x"bdd5715d21974b77");
            when 33231175 => data <= (x"e70f99bd02137e35", x"3a75b593cf844650", x"439896e3f7eaee92", x"f328f39328b8834d", x"6995c5a00bbd62ba", x"aaaad2a334243523", x"2fd373beeae84ae4", x"ee34b93acbeb6c80");
            when 13864414 => data <= (x"715e733b12e3783f", x"676d250e79ecfe71", x"6b9f6619841ae5e1", x"94433f3f2481b3ba", x"450f9b6b71bf787b", x"b4d296448f95bba7", x"6b2a1b3aaf83fe9e", x"52448c760bc89f00");
            when 33367987 => data <= (x"d75904c105afff75", x"0f5cd65c6340223e", x"e658a32c4cedd390", x"e0c5e6d73ab4eb95", x"38ccd501c7ddb228", x"b36988d2f734a597", x"12ce4167b4461d72", x"020e1393ea480e3d");
            when 25986820 => data <= (x"1ae6afa16a7e5385", x"44fae49c4ace1d67", x"db55d7f0bf40e229", x"556b5ed73cf4e599", x"15de41bc95aa4571", x"6855ff10e806388d", x"6ffc0ef1776129f6", x"55c6fca10eb31f8f");
            when 12351685 => data <= (x"b073c8da972ce6da", x"2becb7e2f4ff668a", x"96198197f513d5fb", x"8d0f526a0b502edc", x"dfc56ae0d3c031fd", x"7f7aa0a53718c0ce", x"1f202c3364ea811a", x"a17a0318ecd09b3f");
            when 27869211 => data <= (x"cf19ea45386de908", x"bef32a4e9bec1864", x"db5bc647329c8782", x"4a707bccf5f15a2c", x"f96cee5b4ab7e42c", x"7aaba598a5ba2379", x"01360056aee876e8", x"656369c9c4bb1de6");
            when 13647194 => data <= (x"36205ceaf41145cb", x"1e5346275bee84c7", x"8067d40ed2e25c63", x"2b9f2223f3a24a1f", x"684b5fda3756eba6", x"5d2089ee922c0ee6", x"fb5646ea3126dace", x"89ae75d5207f7042");
            when 29203264 => data <= (x"7ee12f28e930791f", x"a237ca7e2370f6f2", x"28630a9b5fc97782", x"f9379909396340f4", x"b6725fd5b38b9663", x"87b36f208d8644de", x"f7133ac8b2fc1b45", x"e9009e1c0def310c");
            when 17940432 => data <= (x"05fba66cbed5a86c", x"58d98898be382164", x"aca843af62abf577", x"fe784df970c6c21a", x"fb1c39f562ed2d26", x"08769e16c3da537b", x"ab61cbf979cbd9cb", x"01b99b6549a2ab00");
            when 20499904 => data <= (x"6f5270eca4c5a201", x"22e913a4c3550b8f", x"f83dda2e56a7cd20", x"957022fdfb18f844", x"8903405e571ad4a2", x"e32a3a386dccd1cf", x"8e5bf3e04393a395", x"c651e182bb8325b6");
            when 20219171 => data <= (x"05417ffc2d35253c", x"69586b73e17ed1ea", x"35ad2a3dad439851", x"8cebd9e8c50a8fae", x"4e38e7e44b739a0e", x"797030aee9fe6d1f", x"198e575010436ff2", x"22c7853033690183");
            when 29362773 => data <= (x"245a28f7fb6a1be8", x"211358c50df2ef64", x"c90faca26a5e7e53", x"34b08e5d626cb252", x"70b22fc19eccc168", x"c36bc5f344306924", x"7da5ce68aef2f17c", x"5dfa998112956cf1");
            when 19217683 => data <= (x"a5fb941c677f9172", x"a1a7745bde959eb9", x"e7231c86a0a5b687", x"4eda1aa15af19a4c", x"544db827807a268a", x"b6651faaf1cbd3f7", x"8bcfaf68c06e3065", x"366e95d1bad7ae4e");
            when 7806614 => data <= (x"16ff400107956ff3", x"1c5326b71e2f83cc", x"2321e79024dbe10d", x"67a2dfe1987cd35d", x"1f8eb6f18a8e9eaf", x"d26bf91a57f69561", x"35fd2975f66a30c0", x"897322591e8b9918");
            when 31180728 => data <= (x"9b259b5cfbcbda13", x"13abd779aa51e550", x"4200135817fc0000", x"8777a3b54240656d", x"f9d9b618c65d6d11", x"6b1bfe61888b3fcf", x"90cc2519602b1d89", x"fa9dc1a05ae7f59a");
            when 17904871 => data <= (x"74e96ce18309e3df", x"66c9eac38f27aed6", x"a2124642377e845b", x"d824fdfbd82b0965", x"d98d45cfb0d40f74", x"225e8aafe2d0ad0c", x"a3ef281f9b9a579f", x"68f3261e4c83c8db");
            when 16633029 => data <= (x"b9ab9ab20a141ce6", x"fa46b19b5d9afe1a", x"e8ab31045f1f6ba0", x"af094b4d70048c7c", x"0574668d62cb97c6", x"6545ce78535caf3e", x"081f4c62e5dffc22", x"ac08fc4a0ff1a924");
            when 13572509 => data <= (x"032b5a1b763751f4", x"843f0f9770863669", x"38f037f0434862e3", x"38c6f38bd6ad1bb7", x"fc381d51fb10aeb3", x"e48cfec536efc759", x"dcda3f4f8dbf1f3c", x"1d45fefe75ac00bf");
            when 30644743 => data <= (x"68df2adde6466dbe", x"e970bd4d9467d6d8", x"dee898bd994e40ce", x"006fbfb3c959279b", x"4250a13bb668063d", x"152295e5f8c5a91f", x"c15c906f997e3403", x"7526e8dd56f3d6fb");
            when 5784929 => data <= (x"1475c3c2a0f3cd54", x"a88f0ced40d871cc", x"95fc56b366c5f4e2", x"2eb5a497cf45b56e", x"987c9c716f71e66a", x"b3393fd934eb03ca", x"792d74da89e004c7", x"82201d85bded051a");
            when 22893815 => data <= (x"9a3ea0abe6b264b3", x"5444ff7749f75c21", x"40f71a8e076346ef", x"3013ffc4fea3270c", x"c4527b64c8ca87bf", x"0a1f44603424abb1", x"53d21db2eaef3096", x"af8ee726e69123a3");
            when 20637672 => data <= (x"a15f91d24ec93a38", x"f2155d175b1b5b0e", x"63b5c1103de29245", x"1f1b199c93c53856", x"fa27cfa55cd9c800", x"bb4a21d760790f4f", x"31bac17f3c39b702", x"4efafc20537a1ddd");
            when 8438536 => data <= (x"1d22ed6b4061d431", x"2297b263825e15d4", x"4f9e98dfdcf275fb", x"b6b647f6a51003a3", x"4e949f9fb21cf768", x"36c4c6a9bf0fd897", x"4346f3ee590a670c", x"f471595209599122");
            when 7732889 => data <= (x"42d2088b596a21a6", x"41818f847e4b29b7", x"e3631a952f583e6d", x"08ba6474b3848a17", x"351a7827b85bab07", x"c89c6152f4feca73", x"c19e8b53b01d7769", x"7147952a6d1ffa67");
            when 10312685 => data <= (x"b7d8a9623acab4fa", x"4e934533f54387e1", x"198fd000ee17f0b7", x"1cc274f04cbe60e9", x"e39762f1a912b834", x"5eb3d19addef9ebc", x"137e40dee1351c79", x"22b370fa22259a99");
            when 1532055 => data <= (x"c4ff1350c2a79555", x"8861f53f8f445c9f", x"5e1c1f89cbcbc3dc", x"6862820e91a04dcb", x"0989a2e452257206", x"88317f85c8f6c1fa", x"082ef8277cc5b84d", x"0bc40fb46c1685a4");
            when 3291669 => data <= (x"37417fe70a182d53", x"5dd4ec003dc0a224", x"862e5ba1fb0d145b", x"d4c2ab7675191dcf", x"6e5564e555fc5a0d", x"8a3f443d14bcbee3", x"afc66022a2c94604", x"f30a6c716c6c02d0");
            when 12555767 => data <= (x"651bc95820a35c7d", x"c3edb16ce27e4602", x"501da866141eb7d2", x"eb816cfa3fc589f8", x"6d88b8b829d80933", x"0e862bfd5ed50082", x"b3ba1967f741b0cf", x"07be171f156d3cb6");
            when 4156978 => data <= (x"0565efe5dada8a7a", x"bc24af0690b0c900", x"7e5d61f2b519c1b0", x"977c7ce28134be54", x"c13485f3ad924261", x"14b86de656bcf22f", x"662792bd1c9bb918", x"3f73fee740ee5243");
            when 26148050 => data <= (x"5e76eab6ca654e4a", x"0131d2815c3a2f22", x"b2e7f54f0f54892b", x"95280079c4f8ef06", x"a2563f037287f7f0", x"b6806058107c74f3", x"d67788d959eab6bf", x"25e3124c345fc895");
            when 18224131 => data <= (x"934a21f9810a6cc8", x"2299616b44ee53e8", x"78f724dd5cc701a9", x"b65aa697622203b4", x"f976a858e4399f1f", x"e2f5615d22b4064f", x"a229feeb6fa767c2", x"b9a5b43c1112968f");
            when 12700296 => data <= (x"f6309bd6ef0a4352", x"6ea3af18787fcc3e", x"58630266c0d791d3", x"0a9f0741fd56a645", x"8f262534f6ebdc9c", x"0cfb47dd29b626d0", x"e5027aaaa1c7cd38", x"5b57e5cb63455a2e");
            when 26782568 => data <= (x"6fdc131b30c43173", x"6890baa97642464c", x"0a0f50c8425b93b6", x"15f17be313fe23cb", x"de795e2705fe3af9", x"2d201a6b90f3a298", x"cbe69647a27fda71", x"f142db5a61d55902");
            when 4431252 => data <= (x"a05cc786f8e188c6", x"1a1f53ec00d7f41d", x"cb17606dffd3c8f1", x"e706747536317ed1", x"133ffa8d2e361476", x"429c50890a800483", x"dbb1d9b319687fb9", x"0a3da3b414880e93");
            when 10092832 => data <= (x"62698308f69d60c6", x"7a0706c7d63bffc5", x"1995ba558302d164", x"d3f6c1a7e786808a", x"12c642923779785a", x"95a760a32c2ce596", x"f9e25108929883e0", x"97023448d6085dbf");
            when 1424417 => data <= (x"80a6b5148351e469", x"4c403ef29bfa4543", x"a6fbf819d005e6ee", x"d4ff2b4d0b3996e1", x"3b6e6482e10ba450", x"cbcc76ddb299673c", x"5b32fc0fd7217ac9", x"77761fb77e510b7f");
            when 4711002 => data <= (x"272ff5eab5ebdb6d", x"6004df9671b9fa93", x"30941b71185abfeb", x"e1a36ec120f05240", x"29ab421ce913930d", x"94907e7e6e1ab492", x"95e76a7d16b53834", x"1fafcab650d64f52");
            when 1111397 => data <= (x"f342a5c2342a99b5", x"ab6524004828560b", x"9a3dcb2b7fcadd25", x"5a85e06b8fa5b318", x"20ec451dfbcff426", x"3d78d2f27d8e9e91", x"3abc3891e5020f6b", x"e4c95a36f5db3bb3");
            when 18334999 => data <= (x"ab7c3470cfeacd5d", x"59dbecf70cd7d01c", x"377adf9febcf6a39", x"11725fa4e2454270", x"431adb3b6b2b2532", x"f55f915a154de09d", x"00d5dd8da751739a", x"e8bf19c293894b20");
            when 10432746 => data <= (x"cfe40153ab1545ea", x"dc58840e096c4947", x"2d2f8fb1bb909951", x"6b48e14a3aac60cc", x"54fc6da414b19879", x"d19f033f4533602b", x"87e8f58c2abc90d2", x"0e22179d2eee29d5");
            when 24599375 => data <= (x"6a5147cfc7d968ce", x"25ea656452bc83fc", x"c1e8f52a3b6b6650", x"ff024116bc72651e", x"ef39d562e43f48f3", x"8f306b63c648bbe6", x"c025d3939120dbc0", x"f1f4ceb029b4e6d8");
            when 11125601 => data <= (x"965a6d07955ac082", x"2082d04009ea8397", x"736109391910f59f", x"83114a7d457539f4", x"9725311abeff6006", x"c9d56c364c56e3e4", x"03ed215ccbc30868", x"ed5d53291f4859a9");
            when 18093706 => data <= (x"cb7c62c6bb767935", x"018216a33cbe9042", x"915caaa9570d37e8", x"196eaf0e8dbf86dc", x"5570e096bc7d4470", x"bee0849acd1a387b", x"df56182974589709", x"4189b0a6b12699a4");
            when 1215142 => data <= (x"43426e32ba3b9476", x"900b9771504079c4", x"487bf8068d56c494", x"cd774b343218dd03", x"2e408b3667ce92d9", x"c9f8f1b72ba728c3", x"93ab03e13a972fc2", x"8a9f58fda9b3ec1a");
            when 30978068 => data <= (x"9dfc5ab5a11e2b90", x"4c9814adf161883f", x"8e925fcf135bc4c1", x"03a141b48bbb43f7", x"e03f958b5f838507", x"63635a0bdac3fc97", x"cfdd083ebbc867b6", x"84ceebefe70c824e");
            when 22736503 => data <= (x"bec89412f9e745da", x"9b500820755bf4ab", x"69fe29b29b7bc611", x"5d92c631a7dbac77", x"7e56e64d9a6b509d", x"b349d16ffd7ae252", x"452ac05ad5ae8860", x"8214bf5da357cf57");
            when 16885133 => data <= (x"7a0ebb78526ce8df", x"cca51f6f7987d535", x"388785ad0f7a9c12", x"0a1d49591b1fea4b", x"55ef71a7e92f45d4", x"c0c21448cdf6903e", x"c3206112833ce63f", x"a67ac19678c0edf6");
            when 30972316 => data <= (x"04cdd024f5e23502", x"41bceab7ff5c17c3", x"4532ec0ed00f7386", x"fdd549e2497fae80", x"4a86c8df1ae86b9d", x"b89829d75af4f07e", x"183357bb0a6deb16", x"6f04f2e5156caa2e");
            when 21496755 => data <= (x"f7c81f701cb09b82", x"a0c9827042ce2cd3", x"120001df69028c5c", x"5299c2c5450021a6", x"c889e8a004062697", x"04f31202126417ec", x"599dffa78325336b", x"8ab5c3495a166734");
            when 25022868 => data <= (x"974bced9f20bf44f", x"8fb171d4a643b068", x"d438c6ebd07b1ee6", x"2d7c802e455cb495", x"48cd4624f2428232", x"46d223b713fb0b45", x"dea65626b3d7602a", x"a198eddec6049b29");
            when 10364643 => data <= (x"0076d96a2e36f18e", x"bf2ffe1eb7960a3f", x"4da401fe417b9f92", x"44372db64db082c6", x"aab87de404cac9b1", x"3ee1cb266918b389", x"92f9e9f3d6e8e370", x"a4cb8f26f7d26605");
            when 826008 => data <= (x"abf36410fb4d4abc", x"365446277583ff8c", x"92d3170e67806b71", x"3d218cfc46cc71d8", x"d6378c0d65ba366c", x"2bff1d7be740f1e5", x"60aa8b852d4fbd12", x"9c861bb75e49afa5");
            when 32588363 => data <= (x"347fcb5f2e3f7118", x"5f337e53b2fee14c", x"a5ee2b28144fb5d0", x"6fc9179abd3b3d4f", x"f5bb58b90404aaf8", x"3c569bafddd8df22", x"fc06fee48eb4c8a1", x"cb269d1fee9f50c8");
            when 29331787 => data <= (x"10b20655a34e0d64", x"3ea7e3b9b38c0bec", x"0ac36ae23cf356e5", x"ef77601709e5193c", x"0355d4a9d48575b3", x"d27de7953b5410f2", x"82cfc2bf8fa2c699", x"829ba473c0e4a8a6");
            when 12424657 => data <= (x"2f7b79d3de772691", x"0ed77975275a4331", x"6e783bc9c9a2d54f", x"aed0bc8029cd0924", x"95f5301a923e1be2", x"e86bb74353cda6c7", x"7791f43e516b6141", x"e72f7ac6f5fa0eea");
            when 27933776 => data <= (x"726b1801c349bb1f", x"7e57e06a8372fd82", x"1a8a63e75b6c2608", x"952772ee0125fdd8", x"a8d35587c49386f9", x"317815d1543e7f43", x"f0e1ceca97d2b3c5", x"ad6c933fd7df5d84");
            when 11463054 => data <= (x"4dfd34863f5d4d44", x"2738e466d1bc7010", x"a319ee4ece6f5d1d", x"666a9e4ecdfeedc0", x"4381e5a53d42a4ec", x"eeba4a7aaf5318d0", x"3e12c0c477377edc", x"3d268895576faddb");
            when 23210902 => data <= (x"c0e959947c2dc748", x"140b0eaa748c731d", x"01cab02277ab1253", x"532b7b4716cd4e00", x"557d82fd220ce99f", x"92b1a3d6f2eef5b6", x"1a673b619c1493be", x"a0dca99f1756e34a");
            when 29714886 => data <= (x"c70846be978c2341", x"eb33755dc27cb278", x"8ea85ffaa8d656cd", x"5f3f529bb1bbdac2", x"e469db06c98d7af3", x"cdf941bd4b8f20ca", x"affc68f56ce930c8", x"bb61647fae542db2");
            when 1051686 => data <= (x"542cbbfc9f0a36da", x"5686c93313b96fdc", x"aaf1d732860a3d79", x"980447d69f7a7ff8", x"ae64651347c80ef8", x"3575e243a52d2d19", x"c17e486a7a5627c3", x"102547c9f678c1a5");
            when 30503168 => data <= (x"b77491daa0bbf19d", x"1fa8b3ce7873d479", x"37210e7909f7e7af", x"40e2635331a1043d", x"ccaabe790e307bb4", x"728f2aa2dfd03d43", x"a78ea898446e7189", x"6aa98ff6ee677a83");
            when 15082846 => data <= (x"e52fd4d4a1eacf41", x"4cd91caf8da08b0f", x"49130a64482f3e99", x"d88ef4a87d816172", x"3e85832fb57b4771", x"9d9bbd7a39a0577c", x"5b5c3632496cfbd0", x"dcc42d1a333dc3b3");
            when 27347554 => data <= (x"5200f3c40c762e30", x"808102c05b7a2e15", x"0b441c3cb93d2453", x"ebab3526039a8c03", x"7af29f13ba68d123", x"d323c77321b6584f", x"e4189d1ab2a404f4", x"098ccab53f6b9525");
            when 27457735 => data <= (x"d06b82aa34446482", x"bf828e176d08b29f", x"c76544342fbf81d9", x"861f48b305d42782", x"6717cf56893aee7c", x"86b3a08372c9e4f9", x"bb6a404d96c22c30", x"73966b88a8154b8f");
            when 10993444 => data <= (x"91356885a4b13bcb", x"94cc8dbe113cffb6", x"97f6aa912660fbb7", x"22798ff72721ac55", x"95e3b14bcb950954", x"9e7292bd2e0560b4", x"f26bfb442045da83", x"e38d59638521d458");
            when 28603107 => data <= (x"69debb24a25ee6b8", x"6c356044ee84c668", x"d386f67427ad875c", x"fb4b7248b6913d94", x"6238e82c4f19f8d3", x"15af787b230e7883", x"b2812ca8f6ea51ed", x"3c7013f6aae32de0");
            when 20767527 => data <= (x"06e9a0a82b283463", x"b7aa0adb5dafae9d", x"423b443a19e07a25", x"3bab2f7a4c40e609", x"3d5215d98580b195", x"561ac765371b547b", x"d6d32f9933fc2121", x"3b82709c433efc59");
            when 12035340 => data <= (x"b8c050310d19b2d6", x"5950743f9f3ad42a", x"bc569dd7e56c0098", x"7da378a33a077dff", x"5e1931f88518ae0b", x"ccc3b3ed01ba1ddf", x"2f3d2bb202802e26", x"76320d32ecc13150");
            when 24514065 => data <= (x"343f6afd8d1bfe0a", x"58a18f5247776dd1", x"b416f3a565b6a4c4", x"d81acbd0f66a2807", x"3f04b9905ed32b3d", x"dbee7af1e7760ae5", x"91d0b600ef147f83", x"6bcddbcb68a398e7");
            when 11047102 => data <= (x"8a2bc106aed2d96d", x"328f604f38ba38a0", x"9b01f478c2b38073", x"e8cd3b80b87fb3ed", x"8a5004cb4947d182", x"797e4c969a180544", x"4b0170ea41a83ad9", x"bb7fb908b2d207f6");
            when 33534753 => data <= (x"c224d5efb88d98b4", x"e84fefaf8d689d0a", x"66bb2de0bc63a6a5", x"64ff5e53a0d69381", x"9c0344ec81ca8e03", x"3e068494f131a672", x"891216c2ff12bd55", x"b3e2891cb1b17609");
            when 25996363 => data <= (x"03c7c543038e9775", x"a73c7e90602efc64", x"90b1fad11d3f4b75", x"62db957d04a07e24", x"abbbe220a3c73c92", x"6949f793df40ce46", x"bba6f006bd4b0b36", x"3b8b7b929bd94fa3");
            when 27953815 => data <= (x"cf31d33c23954e06", x"cad9ee0d1f787df7", x"ebf9123328a72027", x"9f66e948f0cc9e5f", x"e23d543d930ecc61", x"7f0902fb0bc0ed92", x"4fbc8befd38a5ed0", x"71ee12fc7bb04ee4");
            when 31429108 => data <= (x"75b71864fe37168e", x"ac202d894eb6cbaa", x"45d854d8ab6228c3", x"1b77a006fc268ba8", x"5ce0946a3394d236", x"c69e6bf95c990503", x"99fe4bd5f8eed715", x"82716ce072bc00ca");
            when 14636684 => data <= (x"215b92a7b4927e5a", x"291d6ef1690768b7", x"15248336b6311ec9", x"7f488da6231b24ae", x"d0fc9cb01681485a", x"68f1674601bafd38", x"2dbda33fb9e2efab", x"c2f5e75d9a65bfcc");
            when 28883784 => data <= (x"5fe2bf4e81c10e31", x"e4876da9efd44a12", x"2f94235617a0e450", x"47bba2422d4149cf", x"8b1b3bb95d051c3d", x"0f57ed7b3792ee45", x"7bb38358294ff5df", x"e7cb4186660f663a");
            when 15553960 => data <= (x"defb286e558859da", x"8f1b9e62c965ab39", x"a50cb58312e57689", x"f41983cd705595d7", x"9d45df041425e51a", x"2b5c92b311c52007", x"116e1338a2e3d525", x"366b5e89edf70c51");
            when 11149039 => data <= (x"a8dfc8e38f7727b4", x"134df8e8f145dd93", x"5321d95c31e677f1", x"001f3a6be4c463cb", x"317ea77c7f83e1e2", x"04c0a576e7dea8d1", x"0496cca1a43e6673", x"ae056734d3989b09");
            when 26312278 => data <= (x"07242c9d80add8d5", x"129f34c73447891c", x"399cc11aa989e1c1", x"e3f0735923502205", x"3eea0a829ec91d95", x"0862301dd8ef3ca5", x"d094691a534eaec6", x"b250ccf67666f35f");
            when 7272954 => data <= (x"621086e25be178e8", x"b6506ca2867ff233", x"71c3ded983fa5dd8", x"d0f25ca3bd3dd0a0", x"b15743d36d2a5061", x"b5acd27e12222585", x"82475767456792aa", x"ab9ff0432e0adea5");
            when 17799498 => data <= (x"b6a2022f544e0bdc", x"3f9c41c34a33e029", x"2bf1bbbbcfc9a5e6", x"29a464d2b048b358", x"e5cdf9571b32c2df", x"d87e9dfdf520f37b", x"884e9e2b2792226b", x"b7de519779f16dd4");
            when 10380168 => data <= (x"bc9960f219bdbb5d", x"888fef37695931ac", x"36ebdf0fbcf90b5b", x"ba28fc69da7a3013", x"bd5a64011b7e116f", x"2c9d27622366c71a", x"6f1c3f58dd990c34", x"1bf4208006e83a1d");
            when 13806678 => data <= (x"d401053914e456d1", x"5238412ffa198909", x"591c4c1c9f07c5b6", x"053ddd51dc104dea", x"a2ba161c92b7a317", x"ca6aac0c34fe7a1c", x"aef0f59a5556daa7", x"26ea3a2f21898151");
            when 31853821 => data <= (x"fbfd745ffd078124", x"ede727886a6a657b", x"3f02edf13931cfb7", x"0a33e91e1bfae6c6", x"4e5a1ea5edfef275", x"a218caa0576a2ea2", x"1d5a3d5102ef2309", x"ada3ef92bddde42b");
            when 6703794 => data <= (x"f82f44922321484b", x"154e803f40421627", x"4b8bd24e7bf63dd0", x"8dacf68ea00cdf66", x"a695bb447c86d514", x"94877a88ab59401a", x"b94e8f35c348ab41", x"7fdce188833d3c50");
            when 10396044 => data <= (x"40ccff6025960687", x"1399f26bf8708601", x"6b4a0a5920ed993b", x"89d11ce5d4b1e801", x"25562263ee27e25b", x"45fd1e1335c7893b", x"109cb9e58d16a050", x"eeed5c2f7e2ec384");
            when 23753920 => data <= (x"6c25497f34776185", x"94fe384c674141d0", x"176a96bdbf2ed2bf", x"f6476ac4bbffb2c3", x"853ddcdca8f0b75c", x"7a09c1613ff18d1f", x"fa34a7e1f9c5e4ea", x"aaa6c2d1be7982e3");
            when 14296648 => data <= (x"a21b50eac596688d", x"db6f6fd79a31dc15", x"6029d58b1b8d3e10", x"342184dff4334e9d", x"0b8f590b3f84df3a", x"8347ac1de7fe0648", x"f5aa7e17a7960903", x"c9d44e898aa4b669");
            when 26667309 => data <= (x"d0baf232119c5c77", x"54e7e70fe2171043", x"3c5a0b10f9c103cc", x"8a1951c4079ee242", x"de414b606c9f362b", x"ec49efe10acde13e", x"32f1e86880016de5", x"a3d2c0e87183c1e4");
            when 15703042 => data <= (x"60a31033ed7df578", x"e1921ae96a1bedc9", x"c951509303a558bd", x"c47cbb3a6307667c", x"c57f46e025738c85", x"1a122f5131b5b621", x"490795e920aa0580", x"21ca0767cd23efeb");
            when 11120574 => data <= (x"af307ffb0ea1176c", x"806cba2035b7ef9f", x"6172627e4e54b65e", x"955d2300ac525051", x"c9ed4d5a6ac95405", x"7ea0f7e308b6c5bd", x"986e55b3a9830e3c", x"9a8206ba7d9851b1");
            when 14603596 => data <= (x"50444fa675344cd6", x"ed04022f850ec919", x"0e25bca12b174bbe", x"5b802ffcd1246ad5", x"30daa67b9bdc1528", x"898112b293e6ebf5", x"4d756cdc63dce24b", x"41bc6621031181a3");
            when 729532 => data <= (x"0323bbd589fa5d4b", x"036da8e24ecb5991", x"9747b091b55166d5", x"e8115ad7f9bc19f4", x"f154cc0a30b8d6b9", x"362ac10039669da9", x"678a41a20b26f808", x"525b7d2d1e9bb8ec");
            when 7497229 => data <= (x"8c014fb7b468f713", x"98334be567f336c4", x"15c83bc9fd4aaa07", x"740f3b0588f43268", x"2e3e0b4fc67812b3", x"85c5f6c65777680f", x"8f2aa0c245cf7ce2", x"b4a834dc08d34478");
            when 24257144 => data <= (x"4c1520ad14f9f84d", x"125f63ed6ca640c5", x"752a6c8b686b0fb2", x"6cf637c11f1ef9a4", x"9a31e5dc20b279e1", x"a70de60efb79b4ab", x"1e6550895f745e12", x"2b0f8c97c668049b");
            when 4477027 => data <= (x"488f125536008765", x"d96bbbcea4a0d398", x"6f954a74dac4758b", x"7730d59999082f69", x"74b79f2072bb058d", x"9d81c8f0705d694b", x"21dc54215ee74ab6", x"4827cccd8cf128c3");
            when 29401191 => data <= (x"d0fab2df44c00b86", x"6ce0c2b68df2c895", x"a72e7baee8b41561", x"8adce575ccfbda98", x"04ab74789186fa81", x"8093acc8e578ecf0", x"a79e3111de148e5b", x"3e06c248851307c7");
            when 18357557 => data <= (x"5b4435474df6b573", x"d01a1fdf837da3f2", x"b6d51f741a40f366", x"006f8678c7a277f7", x"6293651b1a8c2cfb", x"252ed9faecd4a0b8", x"d0f948e1a9e5983e", x"158c23c96ef0dc1b");
            when 22403303 => data <= (x"5c6214c48432bd19", x"cf34e54bc2eea1d3", x"4fe0cde1011b63a3", x"0d6bf510d7e70bd2", x"1b79d66fe20e6245", x"0777ffa953ac5e03", x"fcb91e29f7c002e8", x"e99b3863985251f9");
            when 5591065 => data <= (x"7778f2be25370f2b", x"614997e40e320744", x"a2d5a5ab41923e97", x"e9e880c4ff51d6e1", x"4efe19dbce534ed6", x"14b564b5ab08834f", x"630ee8e4eec4ab34", x"c53b25e70eed659d");
            when 4201925 => data <= (x"b32821d738bf327c", x"1986aea61cf2e0f9", x"24cc8e8eb8d2e5fa", x"ae5802f60e126c51", x"b12fd4b605022d96", x"20d84f824c6cac89", x"1f86ec39b96c3ab6", x"310eba349ada0dd2");
            when 13796950 => data <= (x"bb495301e9cfdae1", x"e28e946bb6b008e7", x"a6022cf51e8460cd", x"559fc869ac40a978", x"fcdb760d94e4c912", x"33020faf93f5784f", x"5d56714d221c4655", x"7ba9af0eac406a97");
            when 8869128 => data <= (x"8d4ddf4124a302a5", x"d7b404216f9ceaf5", x"e865800f426bcb44", x"d672e1e5be1d189b", x"32a22b3f6fdd07f9", x"c156509962f5b86a", x"b2274db8d2877f83", x"483342311b0df2e6");
            when 30552480 => data <= (x"6880246298d5a875", x"5a56aec1238398b9", x"1083a065bfc39a1d", x"4bb3bf1853b58208", x"34b561ec9d89e3f2", x"f30b08ea1e74fcfe", x"04140d9facc8369c", x"1c7b52a951caffcd");
            when 12151005 => data <= (x"b8c0db9c5561181c", x"b5d3f187f4b99271", x"d70fbd93de37d9eb", x"6c753748ad835fcd", x"2aa6aa98a63649bf", x"737e6c172000c06c", x"24f1fc5e2050aef2", x"04258e906a6fb551");
            when 23574971 => data <= (x"e294c21ac337eb88", x"d02a110e53a873e9", x"f745e596ca0844a5", x"1fceda6edb7b7ef5", x"b582e8d7785e4a03", x"af454a714af187fa", x"d63fade682b50dbd", x"a7cf0ba6c57f97e6");
            when 6079144 => data <= (x"3e8a4f2ed2486577", x"f5392c30c7357a9e", x"5c7d603c3beb390d", x"4a2b1f7971951e1b", x"1f20baaef9ee398e", x"9c7437f42b148252", x"bd940a26ca463e51", x"5fe48e81bf8770fa");
            when 29679738 => data <= (x"ef5f8782665d834d", x"7aea6a5be584bdcb", x"b937f569a186d1f5", x"3a18052149e9c20d", x"54a5cdb362a9baf2", x"092ec637a556d94c", x"69e3456c853aedd2", x"212c73dd306fb95d");
            when 21985580 => data <= (x"6023eeb28b1d96d2", x"e538894123ad30df", x"bd2e6fc6144bb76d", x"1a38b47d9bf1dd42", x"c1b23ced1ced0b37", x"972dca388af8bd51", x"1b8abc2ee0463761", x"abff1e8a6e554d71");
            when 1725887 => data <= (x"1fea86a10268382c", x"bb54b8db496496e6", x"a152fef96eb00cd7", x"2909e6094e68d677", x"804f75598554f407", x"9b3b489a6d7b2357", x"123ade3f53ae8b52", x"da77d8b337e2c750");
            when 18094316 => data <= (x"f022da2388ecd7e3", x"75bfb7519d04f058", x"7b6b3013b49c8140", x"8e0295608706cc68", x"85dbbfe34da993aa", x"708bf579205fa31b", x"74ce72a6751712c5", x"357e4c59c85c3841");
            when 14092078 => data <= (x"cd0e943f6179a49e", x"cc22c55537e11939", x"eeea11a6d254920b", x"b61cdb60cf693467", x"14bb587389bd93b3", x"808f7eafee69f54e", x"fecc1edd47b8f440", x"cd89917008effae8");
            when 16697515 => data <= (x"a44b7eb68679af28", x"c13d20ebc4527b06", x"fd0b3830f6098276", x"aef9b60041aa3a03", x"e3d54f97189d5db6", x"80b508b127ff7b4a", x"a38c5d1c0c1cdcde", x"16c3dd63500173c7");
            when 1324215 => data <= (x"5b5c34814909cffb", x"90e5c9309e8706ee", x"1f817aaf8f137bbd", x"ced1db6ab3c4cee7", x"aef81f1e59ce1455", x"4cc5da2bce0db26e", x"a1c3c6027f184fd6", x"298dea9220db4b61");
            when 22565610 => data <= (x"0a1b9a9b51245c90", x"89b15740b2280b2f", x"75246fd931f673fb", x"0c7ec85826c652e5", x"05c0af282134b74d", x"1e81947f6d867abe", x"0a5f5f39cc2d7590", x"34cefde71d4ad15f");
            when 13447473 => data <= (x"19e1ffe146a31c4d", x"791c98ad0c262c01", x"9fe2755850e274df", x"2f9e9de5a2315239", x"c400554f4edd73bc", x"f87f6b6066c7ae49", x"abc877c1c4591fec", x"c59a4b3f853afe75");
            when 17314585 => data <= (x"b6f12b53ae0a5b7b", x"1fba6556a84b5264", x"0cd27d3a10a19747", x"5b6e48186a34d91c", x"35b00e2c02ce4102", x"4e06582e080177c2", x"f76dd13293d28ab6", x"031d6ee3c26823d9");
            when 9098068 => data <= (x"a248753a94cdcc20", x"81d53d8c06f8fd54", x"032bc4d68a50e452", x"ff66ce8c6f3283d2", x"401762062d62e3d1", x"ee722d291cbafe39", x"bce96b0ddab628f9", x"fc50013b9adaef58");
            when 1029040 => data <= (x"0b78dbd9e87a1342", x"d81fdac7481f9426", x"2fc33c3fdc4df188", x"2a0b5aef455c89f4", x"706965db78f85e1e", x"1a7603d32dbe02c8", x"c642424dd5260607", x"ac1b2f365bd1f0a3");
            when 33098026 => data <= (x"9dcb156dc5f7ae0f", x"d1a5da83dd8abdcd", x"a6680c98d359a9af", x"86201cb82236a256", x"b6a906dab49b76ea", x"01115cd1a734ed65", x"c2df6cf8ad48d90f", x"777ca590bbdc7477");
            when 1096935 => data <= (x"930e194b5b6beb95", x"0ba576371c6f5b07", x"9dd83308853cbb41", x"7bca502931c93b25", x"3739b128881b3ac3", x"1b6f01d4647c4c2c", x"0bb19f97c8e50f83", x"f809fdef8bd71450");
            when 30518332 => data <= (x"a4710ae083ba8315", x"bbc883cafe806123", x"b357550c8d87095b", x"c1d04405f127e112", x"b8fa847524df69a1", x"e5827c54e3b97cba", x"bb3144f4dff8e6e3", x"dc662ff3523e0162");
            when 25739684 => data <= (x"e33352758e0e7f47", x"5b40eb6dc54d5c4e", x"893fae73807231c3", x"af4da6ab5deda843", x"d0baf4599e732c8c", x"2e3954392197b7ae", x"6137dafba2fa24b2", x"eabdf26eb3906321");
            when 8014170 => data <= (x"0225c36221ff5ead", x"2ebe9c63c803fa96", x"8d5c11d5e722456a", x"c31cf82338ad6087", x"da7e842ba41cceb3", x"fd5f2b549b93279b", x"5ad54af46132e584", x"38a5742c5ddf4f56");
            when 16652400 => data <= (x"a1861aa36a795a9e", x"a2042ada87c5c631", x"ac821f0967d5edee", x"43eb23e45fff32c3", x"3e3877fcff1a1d52", x"08e112545015764f", x"30bca22ee0aa1c66", x"b16a088199f99765");
            when 7463412 => data <= (x"d192b54582065c9c", x"8cc7d5c874e49c8b", x"6a99e4818b4e9fb4", x"60bcdee154d85d45", x"c3ace06a95b9fcd1", x"f456ed15fe22f150", x"e452eec2100158ed", x"d11c25434b4bb9ba");
            when 24203723 => data <= (x"934b1bec3a411ceb", x"ed028ad55fcc805b", x"02c867327c75d64b", x"16e5a85c5d061d34", x"6bd051f937c206c1", x"40ac1790c41b2671", x"4ca51032994ce2a0", x"f5ba114ca1640e8e");
            when 25822384 => data <= (x"4d21bed4f3f095fe", x"da87c47c5c3b2d8d", x"7a41ef8765cd4209", x"be2faf047229e50c", x"16496bc82184f4a9", x"a66942ccaffe5e32", x"6dcb74ae5a9c3c83", x"7a29648106fa0029");
            when 17850501 => data <= (x"61a28b15473c4800", x"ce6bc57e66e28cb9", x"d11f7d796b43d204", x"d224ec084117268a", x"a0882d35cb7630b9", x"9765c04109e43e14", x"27998f6423db9ff4", x"33b873eb35f1edcd");
            when 11369004 => data <= (x"5d07935194c240f4", x"d50ac4781a58a1ad", x"28d18dce77874df1", x"a1a953feaefc91fe", x"5aba22db57a958a0", x"790475e707347a54", x"7565cc6c4673bddc", x"5bea10718603296e");
            when 25572177 => data <= (x"f62f122da0b0eb34", x"b357b50153d48864", x"3d563fa77f488393", x"f19f25c9b480faee", x"fe4aa79094a7c126", x"e860488cdf66f831", x"bb0d249b63b9e960", x"440876e19f2e883e");
            when 1957178 => data <= (x"173e799d91720910", x"3238c10d1c79e9d4", x"b0043fdc4ccc65ea", x"e2313fc03bb7eb9d", x"a6b359c8fa6aa6fb", x"43bf41d488a077ec", x"b1d046aacc3e4ec4", x"54bc3c241ae88f20");
            when 4500452 => data <= (x"cd3649c1e1f2017e", x"75007371008f7fb8", x"1359d3828d847621", x"be574eb62ef4655d", x"333101b41b0fa1fd", x"97644fdf4bf02ee7", x"87fcd49e1657e87e", x"68f0e5a53ed9c976");
            when 33510843 => data <= (x"dd97b56091e07a5d", x"f6e029a09639aa87", x"610710eb77543ccc", x"24ebc7c39aef315e", x"e2a90a9839cc32a0", x"3784b4900687f74f", x"c2b4dab3e5bb38d5", x"7ab708c860dc7214");
            when 4858097 => data <= (x"6ac707261f3747f7", x"bbfdc486defb874b", x"da45a62d7fed130e", x"67e8bef598901d48", x"7643d077c60c0c5a", x"9b6b57ef70973221", x"58353716bd662826", x"756308ea9a3e7a71");
            when 25204446 => data <= (x"76ee2d8658d87933", x"b16be20244fe05e6", x"f39a7e204162c4b3", x"03413fb2e5b3f76a", x"c0fc9e30acdd1504", x"aef24e16adc8f9ab", x"1cd5797a6c3dfcc3", x"fa858e1fc546fcb3");
            when 542645 => data <= (x"276aff407572f6bd", x"fbd660b14ec0d491", x"8f4bbf74d6d1bdbd", x"7b0ecb6da2f99750", x"5631cf19edc7cb70", x"4c218da6a97ec600", x"12154bbd00d0e243", x"26a822027f0774d7");
            when 21057863 => data <= (x"8b13b89ef63c8c85", x"78d2a0d2e07acfa9", x"b37d4e14991f613e", x"6435448792ba29da", x"4956f34a3dca63fa", x"8c0bf566aa10a046", x"668fcabafaacda36", x"862c1bf7aa200cca");
            when 25265445 => data <= (x"bdcf91155429ed1d", x"1f8acb6159b80f61", x"3706b989788b2e81", x"60dfa14eb0b2f698", x"2545f09dc4aee048", x"78a724cf8c9d7b04", x"ea73ee29050cbd48", x"27b9a21f6eeb1a23");
            when 16339276 => data <= (x"b72152ad88975399", x"d467f2f7f2fb5875", x"d9d3dba372e56597", x"847454f108f07330", x"cc6b0b55295b7f9b", x"98d5958b8b389b16", x"6de302d0c8f1b5eb", x"188e848a923a7ec4");
            when 15578462 => data <= (x"cb9e0bb525ca5671", x"794f34ebcd75296b", x"ab3ee8de620944ee", x"bb5b8bcea86782c6", x"24afae56dc05f912", x"80bbb24eafeea7d5", x"ba09c96c08cea947", x"b8d3a77563c020ea");
            when 26905406 => data <= (x"3aa48619e7fe7ac8", x"118a6b22920b9e89", x"9bc89cd1233c6075", x"5e8048e8d1cd182f", x"03904d3b2ccfe08a", x"2f0348f1cef0262b", x"d6aa20f2d96b5287", x"89c14ec4a95c36fc");
            when 5102544 => data <= (x"7f9f61edc8472653", x"dfaf26e81c27e31b", x"56ea4d3cfba64797", x"d7f75f29408f78be", x"4fde1c304be257a6", x"1a82814e58d01c24", x"674e4a00b1bfe52c", x"90f607c779d25ecc");
            when 29358205 => data <= (x"a3bc797d7a039d0a", x"d620cdda3d6892e5", x"b8345f6dd329db4f", x"f190d44f52217494", x"1fb4024bdc684b87", x"af9238e55cd53683", x"37c3cfb1c8c6f75c", x"0d0cfc948f9882ba");
            when 26433835 => data <= (x"464c169c8df158ba", x"5a2446b2fa8fb118", x"aff288df84dd03f2", x"4f99b0d192f73dce", x"99025c99c75c8094", x"e165bdc84a6ebb06", x"3ead51cfbfdcc554", x"846ad6c5bf742af0");
            when 25675192 => data <= (x"fb8113c8f185b216", x"6346096980a67cc9", x"75a9e8e9f7d78e66", x"1b254f7d288b4856", x"15a9c790fe3fea95", x"8bba05874552fee3", x"71c78db0d894408e", x"00f04a61f5e1b7eb");
            when 9728482 => data <= (x"632906fc444832a6", x"2f0d7f3826cfa71f", x"0f68aebedbad4385", x"5ea73cf3120baa57", x"7d22b2f0c7c50240", x"0eaa6aef61e832b1", x"9cc091c16375e435", x"9412d44166d42a34");
            when 2639094 => data <= (x"569ab17f118ec987", x"7c40359b67ac5265", x"aaddce6a1bd67896", x"b97dc781fc43d3c0", x"cf4f0850dbb971f8", x"d7d998287a9afd20", x"f9448ac0b3146c81", x"2da8dc5927424268");
            when 4607178 => data <= (x"6741db0f4410da40", x"de4ddcfb778c5dc4", x"6e00eb77169ca8e6", x"57983e5875e268ba", x"0f96c293306351bd", x"4d1a92ffb347f1d1", x"adb7c3450c4a4513", x"516d0b3fa66eda23");
            when 18048881 => data <= (x"66d8a2242c216a0f", x"83c5a6ed60eb8a4b", x"99ea823592426a30", x"6d735d90a286c784", x"22529ca62b21ca2b", x"4370bd3c37b0f4fa", x"391a54c8f6a53039", x"9a7a457420989171");
            when 19040727 => data <= (x"4f77d066cd3e5fe8", x"b59967cbcf8c7f4d", x"f68f5620e45db9fa", x"4a5d953c4c25f811", x"ed865aca7792870a", x"1dc449472ba3159d", x"ce726d9542fcd032", x"2662dcd2a2c3be72");
            when 33824145 => data <= (x"51532d28f899f47c", x"650dee9f09321a86", x"0b4cb7497245d364", x"6b613fa163ea9073", x"653651dbe5bb49d4", x"b3a40791b9512084", x"176049ba3de81c61", x"275f4d24ed66bd90");
            when 12453007 => data <= (x"7f29b505184e3524", x"b7897ea515f78a8c", x"87a36938c048e39b", x"378e3aad2f171ff7", x"e600546b5c8cfb3b", x"67e8eb51d4d8c5b8", x"ac325172591c099f", x"7d8dd7a67277dbf8");
            when 20851198 => data <= (x"8acaed904b9c41c0", x"e1deb237aaff4f15", x"e748668a1129a236", x"896ed44f3c54f146", x"7ba06fe94e883b78", x"92b33d586f3c15a9", x"441829794bf4f663", x"b6a62837702ceb64");
            when 26073290 => data <= (x"fb05d64129a361db", x"a29a63381119a0c6", x"971223259cf1732d", x"0f9471908a8c39b6", x"a61224b72da100a3", x"d0b0ac8314119904", x"98252bf89ed27138", x"3ef25ed3a373c950");
            when 3248605 => data <= (x"3dfedc443d75096f", x"30f2f1ad6640e412", x"082192118f6e2be3", x"b9cec49e6a62f077", x"0f44e94180bbe0d1", x"76419554b1902662", x"479ceff3b06e1285", x"6f6ea1ad28f7f97e");
            when 28295586 => data <= (x"e856e245c1aa56c0", x"a50d6c6f1534a047", x"bd0497d3619774ba", x"e0af9c4c3b7d9e27", x"3e0728a7c34c501e", x"4f59a319d0975f1c", x"20bc8a15cf8576e7", x"5db6489a6a54a32f");
            when 20630233 => data <= (x"aff639095bdbcb08", x"6078981c51a6f1f6", x"73d8fb3d90dd8ead", x"a34eb61e8e72a131", x"9cc79f84a1dca03e", x"bc8bcf1b2151b36f", x"81e710db12b0ff37", x"b2e885f0b59f4abd");
            when 26138287 => data <= (x"e2547dc28e493d50", x"a4bfc9a9b9c639ec", x"d8180e80460f8a78", x"01fb30e4d777d9f9", x"a1a1b7c0d6316b38", x"7ac9f4bc5dbcbdc9", x"be8b55272eaa7845", x"f6f6d5885a228c9d");
            when 20474807 => data <= (x"7ee3e481fd609f7d", x"b03c4a51b1c948fc", x"798c8dbc4dbd9af4", x"34a239d7b6021924", x"97bac95d1ed29f1a", x"55ebb4285f63504e", x"48531ba26abd3860", x"4864eb661f0445a4");
            when 24037077 => data <= (x"5c2b5520e37e1c9b", x"1eabe4fa699ea7cd", x"c3e42d26ec44f4c6", x"a252d495a93102f8", x"8c5e5e338060289b", x"943071db6a26534f", x"5808dd8df7fef0dd", x"eb148a294f386853");
            when 32738291 => data <= (x"8db000882534f13a", x"01f03555032d98f5", x"4f0ad84b935e0c27", x"880536ca7cd095b8", x"37e207525f686a4d", x"c3a8894dca646a37", x"80a5e5f8e3bbfa92", x"9b5c5918840de247");
            when 33143113 => data <= (x"1ea6f591b3c93936", x"e59245dcdcf7a187", x"368e7da7aec202a1", x"efe23dd12c8ed34f", x"cf823acfca562c5d", x"2be70be9eaf2b4e4", x"c6823e9fb247db28", x"28e27f05c602bc1c");
            when 23579858 => data <= (x"d9f6037d66b50c91", x"a854ede311b8f00b", x"f74a3c0814dc35d2", x"b800be1c6e2a6381", x"4fa4f6609f8929af", x"9e0f25e1b8436bf1", x"92d91e61542de949", x"58282b3e956bb076");
            when 25548494 => data <= (x"7efed975783beaed", x"f3cbbe804d91be44", x"352763800826ad8d", x"d8fc4d194ab86eda", x"25980f304b765208", x"9a0a3e575bc0eff3", x"03f0c075cd4a3675", x"232185839387a27f");
            when 17318242 => data <= (x"ad4f1d08b9947494", x"79256655b1ba2d4e", x"f4431df0edfb65fc", x"6e848f97a2baa151", x"784c121a94517b4b", x"125ce79c6e166bb1", x"ee19413c2a3a2204", x"b75b89b89967b532");
            when 23516383 => data <= (x"5833a15bdc10ccce", x"577387ea87a033ac", x"13330e05b70875ca", x"a3388a9997c7e8e6", x"12d0dffae0ada307", x"7a67a3d71a983387", x"019930b252213732", x"0db969aa46a49906");
            when 1385819 => data <= (x"f651b2cab9d12819", x"f402785375730b32", x"b545cf7202ccc83e", x"9371553339df2060", x"56437eda216974e5", x"26f0975924214e50", x"f2dba1a7117b8d66", x"d8368708f3dd8515");
            when 10854411 => data <= (x"3851890bc5d2209d", x"8b0c999b2a8f9d24", x"18ce3ff51a963f4f", x"cdf859cd7d860fbd", x"bb9b825661a26183", x"18cba0fc7f7f0ba1", x"6b5ac422ad893957", x"447e4398a988bc98");
            when 2809853 => data <= (x"8e7f969816038490", x"378cf9a44c8cd105", x"e0ff9a083710f8b9", x"13cad7868267751a", x"b9001bff77409d91", x"f96a44bba4314390", x"c556f39f65edaf2e", x"c7b0a7c6c9af77b1");
            when 33303732 => data <= (x"09a36414006db7b5", x"9f88b7f1a04020e8", x"8b69182a01f30942", x"78e80dd206a5157f", x"1fce39a9eeef72da", x"cb614f5e0f1c89c4", x"6803a9e3c32c6c40", x"deacee2c11be0d68");
            when 6414302 => data <= (x"b76b3be270e2b2da", x"629e17bb587ffc95", x"6fe8caaf052e924b", x"08b96bec4a7bf26c", x"9a3744e8a9c920d0", x"6e3e9356d4530cd8", x"298b2674da89ac6e", x"69605fad184df616");
            when 10231471 => data <= (x"73390932b645d916", x"ec50df24330cbb78", x"c821e2809b7e1c07", x"909c53a7e89a57cd", x"6f90bb5e789a989f", x"d5213c34674de799", x"614333bc5c26a799", x"cb49837f05708073");
            when 20973404 => data <= (x"e96b71630d9afd02", x"5893c1b7a0ac740e", x"24e8eee0881e6464", x"c5a7aef6d54af1e0", x"532d3b324566030e", x"6fc107ce0359a133", x"bbe5e659a2396b14", x"23db503a44193a39");
            when 19852753 => data <= (x"10c66c65849362c9", x"5ee4418826257de7", x"de11c9895f3701fd", x"d79832b22e3bb664", x"ca973d9e95d98f1f", x"76e6a7009b9db172", x"6ec85c9fafe1a4a5", x"2f3d9e8bb03a989f");
            when 10884647 => data <= (x"2c58602b49e61a24", x"793e8bb09c1fc35f", x"7a25d63e915d9a0e", x"23d22e6413ccbd43", x"9084c1352135cf41", x"31aae6c29c0b505d", x"e3b5c6f5080a21de", x"f8c168c75b2050f5");
            when 10895200 => data <= (x"b6ea9e5bf31f39ba", x"a3b483e01edad9f8", x"f218203c3ec4cc0b", x"33c8e009ee70df28", x"63e89922c45011a9", x"3558ad19e79032e8", x"b1641dce2de39324", x"d57b863ff6cfc53f");
            when 9428748 => data <= (x"c32d873dbe4eafd2", x"67b7af91ae9f2500", x"a569a9e87b3c0d02", x"8be46e56d642751b", x"53af24be2e093d5e", x"d1897832e5af3dcc", x"d9a00a34421e7251", x"ef8693bc37795244");
            when 9226185 => data <= (x"b4ece46f5af63999", x"a5c902aed83b96c7", x"694798d1ac9166c9", x"fb2401459476e3d8", x"362645b1fb951430", x"0de19d45c633a4ed", x"e00bb302f95a059b", x"70f3ebb1712f63cd");
            when 23804036 => data <= (x"3bef95c8ac21b489", x"0abc66f96519f538", x"2d8419bb2a95bf19", x"7b926f5674d6e557", x"02754d7b2b74e89d", x"7c550569d0671a15", x"7d04ec5063f6638b", x"8a781635ae22a309");
            when 30282662 => data <= (x"78fe5f28dcca9674", x"3523f0ae6c17187c", x"3ad98bd54377748b", x"b71d03bfc9dadbb1", x"a35b2786af8d1d1a", x"9c98d2d1da54755a", x"17bb9aea29a36541", x"2f1b7d79b68e9b62");
            when 16191681 => data <= (x"7f3bebfef39109eb", x"f484050b84a7b195", x"fc8a184ea8cdc576", x"cfc76a11dee6be01", x"30ea251ba9217354", x"245e0a6b433e75b1", x"49050aa922e40377", x"9c199af45b0730ac");
            when 32475751 => data <= (x"16485d12d4b6c002", x"feee3485aff16e9b", x"d206b54279f7ca24", x"e09545c156180a13", x"ea8bac3f42bdb696", x"70117c80fd12f30d", x"78c4c8df45a65f9c", x"2e9ef903c3108512");
            when 32844093 => data <= (x"7f2c378dd97d3003", x"2dd43978d272da2b", x"4bdec5e91c42a02c", x"6279d4e8f1295efd", x"0513d1741c2de297", x"f06810de23de99ad", x"5c20e184f843e071", x"abc3d864afc29adf");
            when 3749167 => data <= (x"3e6462ab645d7590", x"b43be3bbc1f385de", x"3d74db9532781046", x"54430e9071216d8e", x"5da4cd8df3e3304a", x"b55622041f0d6b79", x"171978b5d2c6f3fb", x"cec44ef9192d5e85");
            when 8039857 => data <= (x"c2637e06227111dc", x"45dea006ab0f1faa", x"c58e489b2cad3780", x"a2e3622998914625", x"f182a855e6de34f2", x"9776b1c0f10ce2b3", x"d0bbc47fdb0d9225", x"d8f244bd45115a76");
            when 17847846 => data <= (x"9a551d768cc4464b", x"a9cc44db2591acb3", x"3f3a3f5ed0687b07", x"828631a5e690161f", x"ff60f93fecf0ba3e", x"cec00615881b82b0", x"c5dbc1f790b07bd0", x"74018bc7979c2c81");
            when 25736258 => data <= (x"24111b81009dd030", x"5547610d974116c4", x"9ba87c5af49c4819", x"db7686472519b22f", x"7d04deefe73e8d1e", x"39e8202222c29d4d", x"d5ac2d55c469eebb", x"49446ee8e4e87caa");
            when 26924424 => data <= (x"dcda16b8e60c35a8", x"ab1b86d525fe18fb", x"deca9aec7c9deb99", x"ecd0ad76deb7f091", x"6ded0b281d81c5a9", x"bff601b53f7c6dad", x"6f65cd44dc593f79", x"42e5be93e3fa1da9");
            when 33284986 => data <= (x"3acc9ac12eca8f33", x"670dbf6a94aa442a", x"042b708e7a47eb2e", x"d17e8f27ec7737bb", x"86e5155f9f52dfbd", x"f214bb26ba128053", x"4a3fdfda8da2938d", x"41e0ead82af4b226");
            when 22295850 => data <= (x"32403cfeefe9d6df", x"a0d6dea3ef241ea9", x"1280ba960dda319a", x"99028ed885cb1e62", x"d6364515a6b29028", x"07832ce2e196db96", x"6a08beac41b19ae0", x"89adc8021e1b7ced");
            when 30368969 => data <= (x"5109d8d2685ec56a", x"fd09b8bc5f21d396", x"70402fb91b85bce0", x"45873e3c074f1a87", x"a3cc96cdf737476b", x"c13614024f1c391f", x"462d52b6f7def105", x"e80e04bcf4edfedb");
            when 28431808 => data <= (x"eff424a8f5149bb9", x"93f774313bbe2a6f", x"7d2a9c2fb67f067d", x"896dfea283257847", x"9e6965c83dc26206", x"1848c34fa29248bc", x"f3de70c457395efd", x"2634925d5b994892");
            when 17466239 => data <= (x"6e9ec9d7244f4fab", x"9d85d505ea7658dc", x"e576ac7269dd955c", x"ba3adb027a852ac4", x"f9fdeb388cea6b85", x"691304a3bfe4ff22", x"a3cd6b0aaeab8d4e", x"5d8b48ad2f78cf8b");
            when 30244961 => data <= (x"969029df6c631b6a", x"664bac03a4656fd1", x"efa9ceba9dee7733", x"e11ca53aebb99640", x"f6552231081fb1ca", x"bd9cc88dfcc020a4", x"cdcab9225d0a747a", x"6174002a2ad37f9f");
            when 28435683 => data <= (x"431aa759a37b7724", x"45df5056596a9bd5", x"49b672a75bc7c9c3", x"d0847e044547c35a", x"81055fbfd1c7357e", x"e0f3ab4d406f9e9c", x"1b049cd1d97ff82a", x"e49963fadcc63655");
            when 14978119 => data <= (x"878c9e60df080359", x"6779b1b8e6bec131", x"3198b94274b9676a", x"bad284feea2c3328", x"a16b2851ad04ec1a", x"9e8e488e3d4e5e1f", x"ffa02519e76dbd93", x"6b9892d44a5fb598");
            when 4421429 => data <= (x"8525024de95d52c3", x"badda8965dee1d24", x"208a4df6618b7d83", x"0aa1a62d801a9e63", x"e98c66280d1c2945", x"3ed8b648bfa2a1bd", x"1653b5508b01ce3a", x"0b0cb2092368b312");
            when 4068959 => data <= (x"814caff76295b682", x"02175021232414ef", x"e4a0714d2fa75fe3", x"65c01938f259bda5", x"e7d36c1600a2704d", x"8fc16842b72d0927", x"d48a85d2b5a8a8c0", x"4ae492a06a4213fc");
            when 18291515 => data <= (x"fbaf0e27e6b4ff2d", x"cab3da40f228f839", x"22a222f472aa28a1", x"3c2521b823c8cc1f", x"02ae42c4505bd363", x"e4e7d986b6a4db9e", x"52122a955f4cbbf9", x"b31204234f749683");
            when 24876914 => data <= (x"7f9721030dfa0c85", x"faf6f7bd77c6a494", x"a4f4fc0c656ef572", x"67526b5cac1e6376", x"6c2b03a81c355aa1", x"b7831fcb0ad73079", x"1b6b2974e5bdb0ac", x"8c803f7f20941af0");
            when 5994608 => data <= (x"e257021e95433d49", x"0c551fb066e3b13d", x"b63eef67c20f7b84", x"9829fcf469e1c17f", x"910f59b629dc4d8c", x"dd97c94fc7222141", x"4c6cc5980321609d", x"861323f1545dfa30");
            when 15055169 => data <= (x"34a267e21149fa61", x"76e470b8cd83a88b", x"0c67e8468ef556a0", x"3f441c83fbb92081", x"309f46065ce152b2", x"ebc77a2d4f4a96e8", x"0fa13cddbf5caddd", x"4314608581518665");
            when 32701078 => data <= (x"c72e5b4fd2a70bd5", x"f5613010599044cc", x"5a384a3a0a42c493", x"34c7d5408dcb4b14", x"f0c394afd6468c7c", x"c6378d51735d7e2a", x"3ee6b0298eecf98a", x"58eff33d01989117");
            when 26363263 => data <= (x"dc3c863e44df3aa2", x"5106db3a71cf7770", x"aa7a3abe8efd4293", x"c7dc6fc737c4c766", x"0a13b2203ffb71ab", x"cc74fc4cb11f78ff", x"f217fc1f03f17c94", x"bb625e05353eed8a");
            when 2349165 => data <= (x"4f6a3ff2d99761a8", x"c36a19af3cdc7ea5", x"46133d7873fb9f17", x"c6a3bf4880280ae4", x"bb377ccab53e8674", x"73fec7a227d9e501", x"6f3b22b843fa0348", x"c79463bc2f19b329");
            when 23145585 => data <= (x"2114679f0da7f71f", x"f3fe8b7b72c07673", x"b2ca2030ace5a9c3", x"6a665b1eb6171ed2", x"b2c1c374691dc96d", x"9869a8bef86b5b26", x"fd0c1ceecaba7080", x"0ee93c2d43187c08");
            when 17500447 => data <= (x"bc49b85648f58bc3", x"848374395797f06c", x"cf341b14d3730141", x"18a714f3f9edc1e2", x"b8ba08ef6631aa8f", x"c2d0c9f8dbb6c0fa", x"9f4ccc41b05cb833", x"bba30d1746d983bc");
            when 13038267 => data <= (x"dc2ff733ec46cd10", x"d2e058c468502fbc", x"68138520e5ac43c8", x"ee2e9bcdb6b88f6a", x"3172fa63382e8a7d", x"7c5e3549ffb9e0a8", x"c0d25a46c64dcd4e", x"469eab5b970bb978");
            when 16265792 => data <= (x"113ddc601e16a3ad", x"84b930ca324151c4", x"36c86a6cfbb04e6d", x"bb8d852f5adbd4af", x"4fee8eeb56710520", x"689a2ce4c4c27077", x"3776204f7abef741", x"9adf489ae35cb2ee");
            when 33344822 => data <= (x"0dcf3f6ca83cea9c", x"46a1667d538fc31e", x"5d7e298beeccc5b4", x"b2490779d8f800a7", x"bfe785848c2e583c", x"78563274b6f25535", x"59bc8fb63318e917", x"c5a2eeee3b8fe439");
            when 14494102 => data <= (x"78ac99c0d0e77e49", x"df55d22c2dc3e2ba", x"b33bbe0c0d922e7b", x"bf1ffee3473d3fe6", x"98393c0cf0c1f6ff", x"5cb4567a542f8764", x"38bd63425175eebf", x"ad52e4ba0661def1");
            when 3522365 => data <= (x"26c71912ec6ffedc", x"2d15947b08d70a51", x"1a4120626585f550", x"7b5382098bb0b832", x"bc7a19347da03f5f", x"54da3fac8e2ed2c6", x"2b8a3dc56f8243c6", x"db12f282653dda96");
            when 20155770 => data <= (x"aa4c130ded48203b", x"61958a3771bc39ce", x"2e63fc88cbe679da", x"159c48bec2a7f0b5", x"48edd5cf5236728e", x"439eb336c1d59cdd", x"5769829849229656", x"4fce9ac0989ce869");
            when 18917373 => data <= (x"99c008135a6795d3", x"fd9afc07690d17d3", x"ebc9bc192c54e418", x"f780cc4beab557a4", x"a58697b8212f2099", x"41a68a3605b72614", x"a8ae5962f8bff26d", x"a042162ed778d2cc");
            when 18569487 => data <= (x"466b3b22a8e791fe", x"66307ccdc453fa00", x"30a42934671c5f9c", x"572d65802ec99250", x"e8e2f71938adc8bd", x"4ff4c860461a4d57", x"f7d336158aa65627", x"9251dbb231f92a19");
            when 33417387 => data <= (x"25ab596e91f10627", x"a2edec457744e42e", x"f457e42a3bb7340b", x"91f0c72544f29fa9", x"3117e50c7436d214", x"7fb2a10811be33d8", x"084699c34d318b5e", x"a776e1e28b734da1");
            when 19066215 => data <= (x"3c5951c190f511af", x"502d0f8337fd68c2", x"484dbb302084a724", x"78faa223145e4488", x"546c21733fe366c9", x"85c24e705d1a6faf", x"cac5a65099f69cb1", x"f28e762dc50bcbee");
            when 20575123 => data <= (x"9adfb14671256233", x"a42085e095dfa3bf", x"2042552227f228a8", x"9da733105707ca7e", x"dad32bc98d3de89d", x"db0431a5b14b289d", x"05e5a7cb33eb8363", x"7ce88eb2598c0569");
            when 27483422 => data <= (x"c9f8c094af55eca3", x"7591176e4d5d883a", x"78eb4d2852b2677e", x"60958fd4aeef8b40", x"bdb844591f454972", x"6c2be361b27b1e75", x"7d7408c0b6b1263f", x"535a5a7c06a7f53c");
            when 24641107 => data <= (x"b70c530f81766f95", x"3aadd5effbf3f32f", x"41d4473a29b31e09", x"184b2090571189dd", x"9e84e7d9a10f6985", x"90923d315ca55672", x"2a3ccefdf7114e48", x"49d5c97a3105aa1b");
            when 7196598 => data <= (x"3716ce0973e760cc", x"9d35a546616c2715", x"725c3af685afa7b9", x"f628c75ac7ad66ff", x"72c8bb48bac1272a", x"8408a15a65471b72", x"132c1e039ff4cbe0", x"bd35bd235b183a48");
            when 14433175 => data <= (x"81942d78b8e10499", x"d97997be83c828db", x"903db752eb6feeae", x"c7e79406bfaf891d", x"41f76b2870e35e86", x"da127ca4e7f5e311", x"b806cdf366bb533a", x"e9a4062c90d9dae4");
            when 11968895 => data <= (x"ede02128d7798c37", x"08a2dfe1b2fa0c95", x"1b2e1e9e4e2e6806", x"b85d42e6803563cb", x"6492992b2569226d", x"33da13e056d79757", x"a6035623b91386d8", x"8bea572abd77010b");
            when 14583273 => data <= (x"2dfaa3a28636a53a", x"4074b7158ddf991f", x"eef30ed7e4685214", x"0aa7c418a9eb9166", x"1ccc41e124c17d1d", x"f3117e1fe48a224d", x"570e0708e0b4380a", x"63cf2c1acdcd27d2");
            when 22655332 => data <= (x"8e8ef2227d556cf9", x"13f67d2818a4d5c7", x"7e2df085afd6259c", x"3b123e8ca50cd013", x"5c679acac9491f95", x"b99089b409e5f8f8", x"ede5a87c5ec172ca", x"6e4feac0491dbc5c");
            when 33056309 => data <= (x"044317f5f8ffa8e3", x"553d5c17aa38bf4d", x"4d7ae999df1f84de", x"2baae89fc932dab4", x"7a25948091bde2d4", x"efd4befdd1b48464", x"dc3fb35ca63b4e03", x"9a99623bf4c2057a");
            when 20888291 => data <= (x"9924de4fa5f3f739", x"941cfe99d5de9752", x"23965e77416b3b7e", x"71695ffa47f3bc5b", x"678fd75658c2d958", x"5383e8f461d3652f", x"3a6584bd274d1834", x"7b17284c6423866a");
            when 15803584 => data <= (x"5793f39c1f0894a6", x"809810c983d494f8", x"100d4bca11f1a39c", x"ab1fe29c638e55ed", x"d0ad6fdbdbe5af5f", x"7cfa26358797a12d", x"b21eb0c7b547adf6", x"f8c6e504d0c8d3ed");
            when 25556489 => data <= (x"208d797c0e22deab", x"8fd5c739208493b2", x"6ab9246e42333f3a", x"cd40db3dee09b100", x"c4370da0d9e8fc99", x"4dd3e930bd1b9e4c", x"b9b9871a36b8f703", x"ee0afcc4779a9a9c");
            when 32467530 => data <= (x"332cd78b64589fa3", x"96a7d50bdf850a3a", x"8863c7e2fed06429", x"f3a6f13a67be5351", x"fd20a1b545e908b9", x"4dd02631493a71eb", x"3dab00cff6a0fc57", x"4a3dd20e4f05cce0");
            when 4685537 => data <= (x"d8b49a9150095e7f", x"15534f2f210ddfd6", x"b146bbef8f825b81", x"5b7bcaba78c72fd9", x"13cfbba8c39d5557", x"d7b1e40573fb2852", x"8dd4222df49f165c", x"8f5bc0aeaff2ac1d");
            when 30172034 => data <= (x"52d69bb201123c8c", x"2504105b168729c2", x"69b5e3cea3fe211d", x"50dbe82d7682e7f5", x"df2a638d0e2995e6", x"f944ea11ac48a35f", x"1e37ea20e98a0774", x"53f7c6a09dbe2b75");
            when 10400949 => data <= (x"774f464ee86c32e9", x"1f59bfca6797ad87", x"4fdfd93f478af243", x"fcb563eda36665d3", x"695b1480b7725c59", x"4959b1e60ccb2966", x"5213e9d54858917c", x"d8a4930ba6ac332f");
            when 2965925 => data <= (x"391f874ca69b8b0e", x"4a518e80ddc476f2", x"d01639aa565447c5", x"54a9d6d6fef4539d", x"85babdcc691149c0", x"9614dd3e5f133ad8", x"33f245becb230055", x"b97846cc252ad0b1");
            when 3678427 => data <= (x"65b0b68b7289f88a", x"5cbe1f33032a4332", x"5df5d30983c73995", x"bb6eb124b46cbe1f", x"94badb2667f67d97", x"afee00954f47158f", x"e2a9d743a17f6976", x"7242e08c306b95d9");
            when 13290344 => data <= (x"dd68d84aa187e4bc", x"00451e9612037635", x"25fb0424a3a6c44a", x"b1b775eae59b8805", x"6e946b7b27e68f9f", x"800341a9e573ec64", x"99118e5a1d18ab86", x"91667d241351abf1");
            when 23346216 => data <= (x"8c9369b7c5204dd4", x"a9a0bfd522fdb375", x"374bef62473b43d1", x"07f8d97ffb6f92b8", x"158191a59f1bd26f", x"44ea70877749ca7a", x"40bff9e9be8b29fd", x"b74c18d2a7cf3940");
            when 27071028 => data <= (x"26622b09a6f81494", x"3e26bc43054df5fb", x"4079ad993014e9f5", x"e23ef96820b53f6d", x"ce0db03673e8a0d4", x"24174f8db4bc7740", x"06070d9ae9f79be3", x"b1a2f53f1bb20094");
            when 29167039 => data <= (x"7ce929330801e9cc", x"351bbe889a153e2c", x"663aa589b8d8326d", x"b17502c4e07be220", x"906d7f755cbec2ed", x"ee5ad43becf22451", x"9e0d5f3dd555db5d", x"b5b7ee6ba375e5a1");
            when 4453711 => data <= (x"ac32769f425f34bf", x"9318e6c7c83949f8", x"d84844d507c0e151", x"e99d317a345a09fa", x"2c01814e0a9ad171", x"843cd9f2698debdd", x"e1aecbf2457a2774", x"6bbbdbc50d9f87ef");
            when 25497906 => data <= (x"e45585691bf8255f", x"4910f289947f99a2", x"77693def612ac44a", x"07fc17658895660f", x"d6697796a754c6a8", x"7380c1e647857b45", x"52d64c51acf924ec", x"5689aa3513694b39");
            when 8402311 => data <= (x"4f24bdf1dd142a1f", x"9d24b901292ef71c", x"f4253988e7ec50d6", x"5d970eea2a8f60e7", x"9a99ad904f3e2463", x"1d4ae33e5d379eb7", x"c823ef43908f1734", x"6e8792cd6b85c3a8");
            when 4644555 => data <= (x"f75123247ed73dbc", x"26aa58619f558feb", x"7531bf3f7cef5745", x"f2a46d3ba623e649", x"5fcc2f00fcd4f248", x"9d2cc481a98483f3", x"42d2a07e4701ba24", x"37622c307632ddee");
            when 25883161 => data <= (x"6ad20387e0722ebd", x"4fe9ac4982617621", x"4cb4b9ad0b136c54", x"4c20a665b322b996", x"2b6a28a73a393fab", x"0537e4b43164500b", x"58141f16fe76b3dc", x"b505cd1c5c5ca242");
            when 16335523 => data <= (x"abd736d752a3fdca", x"25fd80c374659c69", x"ca4fd4458c39827b", x"585436f6bc3d503a", x"de1604785fd2862f", x"22c5db338a195f28", x"335478e06a83de19", x"6a03304f578e5671");
            when 16909749 => data <= (x"b4511cb4f4564129", x"cf6405b04f9663b0", x"65102dd0880ac3a6", x"fbfd8d3ca77618e1", x"b9e770b27cbab155", x"39cdbf3ee18d0d8b", x"545b5e6d46cf363b", x"718dded2f4add9be");
            when 25522743 => data <= (x"39571a7169dba2a1", x"b279518e4c041358", x"7b3359c7ceb74c12", x"509ce866720d70a0", x"405f64474f844b19", x"9ca979e2b261d00c", x"a3d7667eea05420a", x"64f1a0e5d4970a33");
            when 23258358 => data <= (x"11efb56c533d0335", x"89fcea7b9fc56553", x"0b2fe6280c2ab948", x"ea17c11a34facf96", x"bd0b9f99d4380fc3", x"f6ad7980547ec577", x"49008e2dcf7abccf", x"7adbfa9ca86c0c59");
            when 19381272 => data <= (x"114f6d765b65d676", x"f677409839cc178f", x"dab27b749be83fd1", x"80c7ca0526b038c4", x"68e59e519478efcc", x"34979f2b8ce3460a", x"b41e439f297fa5ea", x"2658398422536cf7");
            when 27671707 => data <= (x"726d12d31d5d6248", x"80e829b846fb8227", x"e55b69408e013f8c", x"7c0c16d3e2b6b288", x"79d7cc3888dfcd7b", x"33a1e7e164ae0d99", x"d9f1bddecf291036", x"95aa4e921d5bc824");
            when 15722110 => data <= (x"1d1290f5ce20b8cf", x"98a7aa37577217d4", x"02118fa3db110fea", x"279bc07d00aaa8fa", x"0e9b2292a757c4ab", x"916946bb1c80dab8", x"bdcab44eb0093700", x"9a1fef75e7866088");
            when 8597567 => data <= (x"a1c67a53b4fbc236", x"124bb7f3be7d1cc6", x"e686fd4aa0df453c", x"62cfeef42b38593c", x"387829da7b1eeb53", x"63989d3b1a5e0abf", x"048354db6e81d738", x"9c8862c5a3f3394a");
            when 12631087 => data <= (x"582263ff26690113", x"fcabfc8c828b4a40", x"41c78449383c1d9f", x"7b3299c54f77ff50", x"45cd4fe95ea32ebc", x"bbb8d81c87d6c94a", x"0592dfc3dad62e8b", x"07ce4e68b774cbc0");
            when 16321032 => data <= (x"e75a2d5bee64b0d1", x"89c58e45d6571c35", x"4e0f3b5108fbce31", x"3ec42f7159f908c4", x"bf43d64bdd28ecec", x"7609296bd0a70564", x"3b625c3fa52a96bc", x"1be44644ed27d837");
            when 28328115 => data <= (x"9a922d34180420a5", x"ddb023c12be6b945", x"896131d89f25349a", x"36aaae8e49196dec", x"f844391ee92b8371", x"be3ea6216f8f60cf", x"e61db066dc6b51fc", x"704080a3e39c1862");
            when 33806918 => data <= (x"a6fe543e47f3c1da", x"907bdc9a5847d5a4", x"62bbbed46d2d6bb3", x"ffc4b1d061cbbc3c", x"a84ee95de4a1257a", x"ed358213c617a1b0", x"749ca73b71f75a5c", x"e741a65c6478c8ef");
            when 8498480 => data <= (x"546541f176d23dfc", x"057ced5b4f6f9570", x"17038888cec12714", x"8a89b0b103c3ab43", x"1375a1f60dd8423d", x"4394958947b24cc6", x"361d612b823be3c2", x"5fb5ff244be179fe");
            when 5028190 => data <= (x"f7b3e7c10d29bd5e", x"c6c324146c216b70", x"c33b5d6862edf8d7", x"8f9d80a0dfd97eac", x"e6f8a835d43bbc52", x"733c058282cede0b", x"490ff65018cdc8c7", x"44e7c58507398ceb");
            when 17099905 => data <= (x"b917be876cbed2e4", x"bd5f0444f2d19937", x"d44176973827c320", x"da3333d79ee39c1e", x"a4b6c52dcb6b25b8", x"321c99c4447ee160", x"19e3b2e0e4a89ba8", x"41a75d37f5b2bdf1");
            when 24718858 => data <= (x"edfd0ca39ab7a053", x"9ca04179b7cdadae", x"77b621fd787dae15", x"d0e63976ad9e5ba2", x"b9fdcaab78b80dba", x"8f1aea21dda0299c", x"a080b67373dea80a", x"f2440f61eb4cd6e1");
            when 7965680 => data <= (x"ba5517179f673801", x"b21bd6a42b2aaede", x"404615b57185f4a1", x"118e954d8b40fe53", x"8e39d752e3263903", x"909b9444a8366549", x"61cdd31856ff69ee", x"fc4fc00cf93b1a2a");
            when 912512 => data <= (x"f9724084113dbc4d", x"183189831be7819a", x"b6ce49243f6f357d", x"68f1d13389e8c020", x"bc9f1341508778d1", x"523dd6fb1e0bfeb6", x"d83fbbdfe849bceb", x"03b3d069d8bd6581");
            when 31627078 => data <= (x"8a67cab8ee72fae0", x"640ee7a7cadfd36a", x"893547246430a38c", x"f7c00c4def26cb43", x"b8df281f7826d90a", x"ec887b632ee07b45", x"c51493594ea3abf6", x"e080455e341c7b98");
            when 2268745 => data <= (x"94333facc7b6b349", x"b8674e00ec4d9e32", x"b4c107be3b269c8d", x"20ce9967ebfb9adf", x"ff64a4c943e341ac", x"40109e107bd43565", x"b035f240777fc361", x"a9c76594c5fae705");
            when 28806788 => data <= (x"fe0f05b2e8bb235c", x"1d66b0536c896a4f", x"65f32c56dbe86226", x"2777459180fc9026", x"51d4cb55985801bf", x"d35fcdd03c4dfa7f", x"85e6ba8afb25f7b4", x"963ef9fe90e12960");
            when 29876085 => data <= (x"441105f545b77f87", x"bfa266289069859e", x"485480a5c38cfa40", x"d9884ca5811703d6", x"d48e61e9ba45d150", x"fd33cabb219b720f", x"daaa08a068983441", x"26267605a3c3d453");
            when 25787726 => data <= (x"9ebf58b01fd39feb", x"3d6e069681f420c7", x"b7286f7c76b94dd4", x"be2594b6456f7e5f", x"f2f1a5cde6ceee3b", x"537e6a883f76476d", x"465adc9d449cde7d", x"c3bcbb3db17aa62f");
            when 31050737 => data <= (x"640a7e13e04d7374", x"398401fa8e249068", x"eaa38566bb35084a", x"fbc12cf556b8ac7b", x"a6b4eb3e038ae5d8", x"6109d3aedd8ab48d", x"31be1933914023ce", x"02bba828cc048286");
            when 18199818 => data <= (x"1682ed223b8b5bef", x"73bcfa01f4a0c7d6", x"c9d75363d14131d4", x"ab00b71164b1577f", x"89bbaf5bc9d96a22", x"337385b4b4c055ff", x"a18b2db36c46f7f8", x"aa12d8893030e48b");
            when 4614306 => data <= (x"a8d9b61ba9f5173e", x"23a4a74e749271b8", x"a66d24341149c90e", x"45f4f2c37d314b40", x"8dc2f8356d0456ad", x"86b22b5332bd3fc0", x"f732e61d4ae73a7a", x"382dfae91eae5eda");
            when 1327823 => data <= (x"d39352d0f7c661c7", x"103cb59db8e32f5d", x"682da7834b4bc502", x"3d50b0a8311feab2", x"aa663a6842a68ee7", x"58fa44169dae905a", x"8b1c1400694af525", x"ae4f499e8cda1241");
            when 27928633 => data <= (x"c4ff399f4c317f38", x"8c0daf0caf371097", x"64cbd83b6f517e61", x"b52dadb8ec53e0f0", x"29c93f666acf38ed", x"58ba453e7aea8d1d", x"a313624a294374f8", x"644e4a7b48bbebdb");
            when 20608662 => data <= (x"d7ec8153fa5604cb", x"5b41013dc3c21e9e", x"0e898112689d1598", x"9069939ba56b7837", x"00d8c40c6b498eca", x"08d0f7f88cbc8917", x"89531dbb68f2dcc0", x"a849a5b9b4968cc7");
            when 33220338 => data <= (x"fb6196212dd2fcd1", x"0a4b40baf82585ec", x"930619f1390d51ef", x"4a2a1b6b51eb17bc", x"99e9cf92a6a23383", x"0cc8b3fd6db8d1e0", x"c988b89f45f2b8ac", x"a3e647a40a44c0f4");
            when 27052707 => data <= (x"15582840bf002e2c", x"1e588fba152ada7b", x"0704baea6be8a9c5", x"24c7121d271ba4f3", x"4f2650a1c4b746c6", x"aa33ec2187e060d6", x"893364cbd14a022b", x"b808c30967da74a6");
            when 31957779 => data <= (x"b68ce5baa306ad86", x"02b6cb121627ce1b", x"36153e2913880b72", x"1e63678baaaf98d4", x"084e1868a1a5bbdc", x"ef31c7a047127ca3", x"028d97381a56674b", x"2f1df5ab7cc853b3");
            when 10288815 => data <= (x"7303543e51862a16", x"bca21b9a1d9e5939", x"e613548d430a27d2", x"30cd647013627948", x"c16d9ff3186d5d96", x"b0d23a35356d9858", x"47f3bed6272e04b8", x"2c691f20f05711fe");
            when 1197584 => data <= (x"88497aaf93fe0e01", x"df40ea29fbb2864d", x"f0de0ca652e621b8", x"bc69c451a83483b3", x"f321048a90189cc3", x"1344c2433c5f3c75", x"2277871c77438b07", x"f677e407cda9480f");
            when 15453510 => data <= (x"2d013b71bebd79a2", x"4685fd8eb5d76c3a", x"5925f69b7424ec4a", x"fa9b7fda4179e66d", x"6d2d08a99527f97c", x"ba64f7d863f3730d", x"9cc1a1c16617f5df", x"e314468be448c194");
            when 25482319 => data <= (x"ba06158b6ea7b4ae", x"7ed0fb61c284b5d2", x"44a374ff31e819b1", x"f1d89b66dac87472", x"d14be4ea407126b7", x"336e3b7281c914fe", x"00ef7103c3db9695", x"2aaa1651c4cc1bdf");
            when 12781726 => data <= (x"5db2df52eb9acbed", x"3173a6cdbe541f57", x"f975ee0a1739a9de", x"5492dd536d789364", x"33011a99035bb977", x"a87b7e13a1c41835", x"ff6105ceeb50e859", x"bde756259ab0c594");
            when 5081134 => data <= (x"084d1f1e24709490", x"86ed9ec36483d7be", x"8d4c5f2c2cffe2ac", x"f622d7a4aeb9e1a2", x"0918c4326f6618a0", x"59cadcba2a87b29b", x"cda2de7c524a859e", x"4b56fa761af61a88");
            when 15209640 => data <= (x"9a39f6363edb564d", x"756e0f7b95ed7874", x"94cde8e852baac1d", x"1eccb56fe022751c", x"6a7d452763a737d4", x"0363ee8b7ccb3437", x"d384fa353b685c3a", x"9058aa539dccccc6");
            when 15101978 => data <= (x"be55d9692c52121d", x"b2bbd140f5417e30", x"b5b72db6af39f1b7", x"b4f4d7b8c4820876", x"5c9541529312be86", x"b67783354fa586c5", x"b9a554a8e211692b", x"e6ec0283adbd8b4d");
            when 14686810 => data <= (x"bbe934ad984ceae9", x"057e5619cbc8ae81", x"92025d8cf644a8c2", x"070612968322711d", x"3b08f6b7b931982f", x"46b6d03854cb69df", x"c6fb5dd9cf3b07d7", x"c769baa5b97abba5");
            when 4930786 => data <= (x"b9be819ad4b9592d", x"87ca7a8ee99548f5", x"249d5188a80661e6", x"90ae42293ea30fdd", x"699b02b9846b840e", x"5ce3c3533c6d1e3b", x"7c5c6fbfc25c00e9", x"1e842cfdb4021bc3");
            when 30096989 => data <= (x"e3970669b522051e", x"b25a3c91af681448", x"022cc0dbe46f2e9f", x"99678600c827ef00", x"fb80214f161e66b4", x"96650606ff8cdc63", x"f9f3c24c53a5b30f", x"fec1946d40610e69");
            when 2190894 => data <= (x"2107508825eb8b1d", x"49fdaae663711c13", x"6de56d86247d8bd7", x"9d1c0095739e90e0", x"02d875bc261e72a7", x"02bf95e7b4ab5dac", x"819cc3cf1641338b", x"721267b25f7d02bc");
            when 22642406 => data <= (x"c6f64d7f1c5f6677", x"f492b57abac70179", x"a736c54ebb9b322e", x"100b1b7fc6d3fd19", x"8625744e59ca9705", x"3c2c04fa0d670bc9", x"d9e073b4a74ff017", x"dbb7cb1bbfc7fbcc");
            when 13542373 => data <= (x"05b184eceb89eba9", x"67c8cb2e0e21ebc4", x"3e232cb0cd93d245", x"e495d01971e9e03a", x"09e5049061655abf", x"567acb0a834c01d9", x"0735e5f9b698757b", x"2d3f95a60d432110");
            when 12256249 => data <= (x"417a0c745109c622", x"c75ff28590e6cc31", x"74988055603e7fab", x"4290928a262df907", x"bf8d7f0e154867b8", x"4e21f56a859f0978", x"fa0b274e60426455", x"7b6293e3eb2f494a");
            when 33357279 => data <= (x"44c41fc14a434787", x"cd6121f2450234b0", x"bde494aa7b110eaf", x"56832a8470bef49e", x"aebf28b93cda60aa", x"6a96f28683cd0eb1", x"c0be94ee5a0a5198", x"c5a29353e954621c");
            when 33383879 => data <= (x"c91922e5683e8f0e", x"6e6b2f077c9d4f01", x"89d14424c0cd003f", x"fb9c8077416a0ee2", x"33914f0c8596f868", x"e5a04bc7ae6c024c", x"e8f9f4e94bb98759", x"355281214fa4623c");
            when 24831017 => data <= (x"49d3f139177b9e23", x"7e83c9cbfe91c2c6", x"9958fc3398c804db", x"71bb20dbf45bd538", x"627aa38d01b7b07c", x"03efea86e87070b0", x"7cd837e709496e7a", x"78d9e35cd2f0aa41");
            when 30396718 => data <= (x"900531e86c15ebd2", x"d2df8fa91de37950", x"51d7e265d8b50f92", x"09fe029199fb953f", x"fd4f88b7e9e799dc", x"b682fb9a4be1b763", x"54293fdce7493a98", x"a60b4ca09cad9d21");
            when 11859240 => data <= (x"0085606f01f1afbc", x"99c453d58bbde43a", x"bad0e5f3c8e62441", x"1e9a9ecec5e320c8", x"33360d6bde7a6e8a", x"1b3932f5419d0651", x"2416de74f9a0d290", x"3f2993bfc82c937f");
            when 1190270 => data <= (x"640b648f3959539f", x"a22e7c32c092dfac", x"053c7a3ecd18622d", x"f3444b948a6ed456", x"b14f1db74b8d955b", x"de90228cc2d89bf1", x"40539814258717e3", x"cfc0a0959734a07a");
            when 2451832 => data <= (x"f5c8ceec7355a24b", x"578b69b74927fceb", x"9be4c76d5432fe1e", x"93e63a4b50edd77a", x"0bd7acdac5768e08", x"0379850052214165", x"340e5cdf4bd86a08", x"5ac2ee9718bbdf95");
            when 28053023 => data <= (x"ebd680ec3de4e884", x"4e4199590f89a9a4", x"686bc830d6d48d0e", x"35ac69e22240e303", x"d8a458393b1d9f4c", x"004007b4bd2216d5", x"0debf576a80e8cb7", x"fcfec1df193b3ff3");
            when 28986080 => data <= (x"38bf3ffa1a337633", x"745f4d3f763df009", x"b8964058fc6dc69c", x"655b7d8eb4a5b8eb", x"ce878f21a2d191de", x"7671ef0de85c5141", x"8d0bc26728c4fd67", x"93635691ceffd187");
            when 9825657 => data <= (x"8475600cf2373054", x"c581409eaea37b99", x"104fe56ca9d9a2cf", x"a15560a67c2e8205", x"21f4ea0a4aa46021", x"4ec93d344bae1ac3", x"69bdbfb3d6598f1c", x"3b68c9160043ac2e");
            when 7033890 => data <= (x"50cf58a893dcd8d7", x"4f71e3eaa5ffec51", x"6fb2b56c7918d475", x"df3dd9cdd519a52a", x"cad4258d35813728", x"77c380221c1fcb51", x"b12efcd23c4b3f34", x"60759119a139cc3f");
            when 15510111 => data <= (x"21c0bc484c1a4d26", x"88b3dad67ed97a14", x"133ed4c615f6112e", x"4171445531332503", x"4d6e4d1a7ed04dcd", x"f033a90d928fe4bb", x"ab6235817e79d27b", x"7899f14fd16716b9");
            when 17208398 => data <= (x"2208b5c0b3505839", x"7c36d463e58b06bd", x"be2ffa292b087dec", x"73eb574bbc90efc6", x"08b946cb101aa09b", x"94a457d8e7be23c1", x"316c891b89c4d846", x"982125ea0da08344");
            when 23206377 => data <= (x"c638092c1a9bec90", x"cdfd9b4be9c5dc1d", x"29c3753bfe1cc5ec", x"1522bf01694311c3", x"3c9e83c693fe06ea", x"2c984bdb6e7d936b", x"474c6d8eed16fbed", x"d759c6e81eca4a8e");
            when 9736343 => data <= (x"0f1230c8538c5a15", x"1fc166397df2ece1", x"0df204db5a09ba79", x"c901f329173ddd29", x"b7cc7943c48ce1bf", x"cf4e0bd8a4190ea4", x"6aa174cdcf22a2ad", x"84e17f7db63a3b74");
            when 7070163 => data <= (x"7316c77a35d8983f", x"efb3a62e6071954c", x"8e458e989727325b", x"3a0959f41a57a2bd", x"740e33e67d224f59", x"29deba935d4ca5b1", x"fda0c4c45294dfb5", x"05756625ded7c01d");
            when 5925841 => data <= (x"7d83b2bec177c8c4", x"2f1a1a7b8e69c0e9", x"ccde4c3b180a0c49", x"5f578dfbf360faeb", x"fe5a13cc7ca99a91", x"c6028c2341fac52d", x"d88f8bbb04d186ae", x"f46d5c2f441f4d56");
            when 30849086 => data <= (x"bf40a58199fed673", x"bc0aff6ad3cf7f37", x"61938bc2586e34c1", x"c2e48490b7c6eb0a", x"0e97246531d55efa", x"d996b3d680b3265c", x"32554e7ba1b9a6b5", x"eadbfd48594c767a");
            when 31793006 => data <= (x"d35bad93f01ba3fe", x"f66fd95f484d0412", x"600958150d096f73", x"875a9d369441db7d", x"e10dce99d812847e", x"370db2536e1b7191", x"0899f6b31dde3b62", x"bb7c47ad7d657ff7");
            when 31843533 => data <= (x"91875abe32d56043", x"cfe8d141e25d6553", x"da56a5b02ba9ef62", x"98d25f992df1f97f", x"e32f18b8f75401d6", x"107a0e5bb572f225", x"378c371150d594df", x"fc61ee5ebe8cccbe");
            when 33189762 => data <= (x"a4161c416bdd98a6", x"cf8e3781389c76f5", x"ef5526bc9b256131", x"0175037f2e8c1a91", x"141f87c7e754780d", x"17315fd67d889015", x"8e26f2d8600af86d", x"fa895c46bc5a1f5d");
            when 20253788 => data <= (x"c23bf07e6b96cf73", x"cc18b654d4f4030d", x"7b098a90a354d6cd", x"8bbce3b8ee49f995", x"34aac0a9f254592d", x"e5616bef6f634197", x"a38b5caf902d418c", x"292c10af04453543");
            when 3448674 => data <= (x"c8deecb0b6e6790a", x"b79a883ae6e2b471", x"e03d828886ff9cfc", x"5ff71ef4425bc2f3", x"b67c63161d29305d", x"70062e77b42b61ee", x"6a899e9e42facf04", x"b211d5efeee65c78");
            when 12454132 => data <= (x"5b9a0a20507b4ea9", x"f38abff5722f10be", x"8d7bfdc2e14911f2", x"dc5536abee067f60", x"d5b0fa8ce815d2ac", x"01a7c1dc856cdb9b", x"a671cce321f5b864", x"eadcaa48e78226e6");
            when 32406169 => data <= (x"3c1127a2f23f56ff", x"5f56708dd3f523d7", x"1410be2df302862b", x"260f4d68ea1bff59", x"a28f51e4f25b5a3c", x"4364bb84be810721", x"273c20550a65e7ce", x"a31982068726d68c");
            when 20234270 => data <= (x"3b24901bf8eeb8c8", x"1e99e2d3585e7275", x"0d755e28ffbdfd15", x"29c7b1d28dabe561", x"2c7ddecb3c064274", x"e806397902c31948", x"eedc154526062cc0", x"2044476d7753963f");
            when 30731749 => data <= (x"6b2106963365b45b", x"c59d748a0f0a278d", x"98ad67e362c4a504", x"61538df43278767b", x"9d6951dd4c70157a", x"8aaff6e5a24befab", x"daddea008371f7f0", x"f04e8c0310b60ae6");
            when 923891 => data <= (x"6f5a835132d10929", x"9e88a26e767bb3e1", x"fe83f0ef3efae6f3", x"e4b34547d1f202ec", x"7d806802847b23d4", x"3be8814e2812ce33", x"8c177a2ec829b9d1", x"6146ac1939821011");
            when 32195184 => data <= (x"2d7d5fb5c11093a6", x"d9f948da2aa7f794", x"7b5a66cc1394b412", x"8fdeada04c90428a", x"7535c8d9d9c5da65", x"799b5315e170d713", x"c637f6aa7fad7158", x"86a868e1a5754846");
            when 6165072 => data <= (x"f2a5d063408225a7", x"4116135f35a54d13", x"5d389945a6e546c0", x"20159a2dfebb9be7", x"a9ef20981ed11726", x"8c306a06d228699c", x"5becda0e543c7b18", x"0c4a3e543f3855bd");
            when 2197713 => data <= (x"3759831645d36285", x"184dc87303e76477", x"865b15ee0f6a37c2", x"5b1641bde9a73ced", x"2a15cd2691ec50ad", x"c3bdff24f6f7c4bf", x"de4598472e9bfb5f", x"88115395fc5b77ed");
            when 12390194 => data <= (x"a48bccde376db0e9", x"b630ad49fd028821", x"a2724b36e5130004", x"ed62341f95ac1ff8", x"a4e844e307a52274", x"1a294703194036f7", x"2d8ffcd94ea17ada", x"2c1293cec4385f41");
            when 19815718 => data <= (x"dead120314ab66b7", x"dead381b2b999ef8", x"6888c664579c7ff6", x"22a773792604dfb2", x"84681c5930b3c957", x"1d3703a993326b1a", x"bee729fd03c0b048", x"eaee6c34a2a73373");
            when 30617857 => data <= (x"5d8444e55fd17d3d", x"bdd57e53801762ed", x"41239b71e51d9381", x"68bc87d21a7b9829", x"8a89d8ec39efa1fc", x"dbe1e274b210bfde", x"4610e50db686484c", x"4c0a9c2f3282c6f8");
            when 9525876 => data <= (x"7fc09c689c3b7e47", x"7294eeeeb9981870", x"91e9586d87e3552e", x"01478b5e7d4af118", x"2a2a4fadc49496ce", x"cc8c8e738e4c790d", x"86f9461b67c8520e", x"e056ae8821f063e4");
            when 23855376 => data <= (x"c19e700b5b995a46", x"8c03f49719ad5e9b", x"cd223ea50fbf0b75", x"addfa3a44a79163b", x"451691f2b90b1d88", x"215fc09168dd9446", x"5a5e94a7d91c19f0", x"3e2ccae177aedbbe");
            when 2983639 => data <= (x"03fd45048cc1fa89", x"9fcf01b99e36a4c2", x"a8e15407ecf4ceb2", x"45836365a8bb58df", x"0ee0a0dc8fa1af67", x"0e8171292b7bf534", x"df072e75b92ee386", x"32aa3713e0b94b94");
            when 18454680 => data <= (x"c64538ebd5c4157c", x"0820d22e141ab74b", x"152dff8b1d2594a1", x"8af4ce40d843f86b", x"c33b60586443d0fe", x"8ce7756126c769fc", x"828895ed16937912", x"ee08ab9572a0d79f");
            when 15254004 => data <= (x"a572d0e09e6ba804", x"d023d1f789d7fae1", x"64785f7efd82fbfc", x"f427fd7d721b87a4", x"8dc02aaff7375b9c", x"2bf69e705a33c351", x"48a72aca772ae2f3", x"a372c16098f78934");
            when 19457455 => data <= (x"155565f255f90c46", x"a1164dd7dbcac0aa", x"32162523fefea3a4", x"583d57f351e5c17f", x"495d30a9ac6ded0b", x"eac2b53cc7084d10", x"4244e55e2501d2f0", x"d2d6dc8c69317ed7");
            when 28945210 => data <= (x"fcbcc3a881830511", x"84537883cf1fccfc", x"44ad2f097b8104ee", x"500df846c6d525e9", x"92b568f9c2631286", x"f100076308a0173c", x"2f0d4337484cea39", x"6d3d908c20105a6a");
            when 15589711 => data <= (x"c043f98b172b0ff0", x"bc6c05cca3e2e507", x"3dbaf927c7851518", x"bd727464c56b6c4c", x"dd8d21e268e1799c", x"b60dba598b7427ae", x"043827de01bb54ef", x"3ef592b94d2dc249");
            when 1116453 => data <= (x"d0446e0282fc9d52", x"dce47d5b512decfd", x"6aee8f35af3b1cba", x"ded5f0c9b88e3208", x"25d0a14a212d474d", x"eea85716e750e0b2", x"51e955a90b515385", x"4f77c644ff4d010b");
            when 23344760 => data <= (x"5f099133aff4b965", x"b710bd17161b27dd", x"18ea843e43b6b628", x"1af01aeaf1bcca0e", x"d39c9b31d767184f", x"cdc7c75c85ef00f5", x"1b883c830cc713ee", x"560ad8d12ce9b3c6");
            when 13181814 => data <= (x"77fc5a1505fa7159", x"b88696f89dc26c99", x"a26881150c2fa24c", x"8ec5e66e9813085e", x"a6a1fd2f2f9f9df6", x"f2aa19ceb5ba2cf8", x"99ac3a4475b54885", x"8479d09a7e023db7");
            when 1835314 => data <= (x"9a3e60b7b6f353e3", x"7a890325d4f96359", x"6e23ec6ea65d4640", x"3834b5eb9238202e", x"019e59c680c98c4b", x"b3f27248203278f5", x"8e6db85d6e69bce8", x"62b25c7c34324f05");
            when 813134 => data <= (x"96b0c5b15bf31ba5", x"dc7f2f8de311139f", x"836d1d57b8628e4d", x"c81d472b301932df", x"ba994851b199c0f7", x"b29e94b1729d09a7", x"bb84025421770809", x"ca6c95766a600f6d");
            when 33292327 => data <= (x"4fc258964595f76f", x"673cd6e377cbbe19", x"cf4261a90def549e", x"fab1269f5cefbd5e", x"f0e89aba6ef69e1d", x"c63ecb8d0e4d97cd", x"be9f601b09070c17", x"098187c3fea6b4f8");
            when 28098356 => data <= (x"96880e24afdad3d9", x"e1b99a6d55395549", x"e10d7628a1227bee", x"346c263a7ff67ed0", x"79c16c3c0362b79d", x"8a98e700fd1f037a", x"ed6ed19fd66ab4ab", x"75bc4e77bac30b9b");
            when 4639765 => data <= (x"179914a4bc4856f6", x"84515d388c5fd53d", x"f5b74cb8fcf27e2f", x"9df44b09911758c1", x"84df9f25fbf1e08f", x"d4496681b79f7a3f", x"a304bd0d115e730e", x"6965a3b2ed68002f");
            when 7394548 => data <= (x"e186cb4c6fddb982", x"f35872015adc1cbd", x"ef63dbf14a27ef42", x"960bc2e5e094a024", x"e04e97fd234fe565", x"cd970093c561f844", x"8efc25e2186863cf", x"05ef251b32dd541a");
            when 19849674 => data <= (x"9f9a2e3292d49efe", x"431fd3da7e3d3b26", x"371c9cbdf0e24585", x"c89e4434ef77cb68", x"e1f080f658d41e95", x"84e6747c7db77918", x"6162b2862f540f02", x"aab2518e0c4cd41d");
            when 27422056 => data <= (x"8dbb620f5d5d35e1", x"f36f13e8c5c1fc19", x"2baffd3a0eacac5a", x"d5da1085b53babf3", x"bb2b1620e39d4949", x"3eff749113dbbf11", x"df2aad1cc6277871", x"d965635f94fa6dfd");
            when 8127058 => data <= (x"05bfdeced8af1f04", x"27993a902b08820d", x"c5b1a6c843ef78ae", x"8cb91831364e5107", x"2753bab9d723032e", x"0f7e7d78157ce1fd", x"3b34bc71e91cd268", x"3a3ce57391378941");
            when 24353636 => data <= (x"f4fdf8a322474f72", x"236d3eba2579f446", x"3bcc6c883b32bef1", x"fbd1b470207eda66", x"3df4bd3f28ad749b", x"738cb3e5eb4c1b86", x"5ce3cf5939c57a3e", x"04ad8f400d1b59e8");
            when 32060392 => data <= (x"0f73a9451f7edc21", x"2a25ea2351a1360c", x"4b90fc9ccc689fef", x"0a04499fc45c356d", x"1f0445d5871ced01", x"6ac2ad72b65c8f2d", x"fb38cf819fd653ab", x"8de003950ec13568");
            when 1017376 => data <= (x"06872cd2da635e9e", x"4d62141b035baa7b", x"77540050183ed7d3", x"c4dd44d532d3bf69", x"ca69b34c7270c0a8", x"1cda2442658706ef", x"846b256c1d54722d", x"435cebef4d47b8cf");
            when 9259761 => data <= (x"40390e3bcf8648ee", x"b8e15a0540d3bf1f", x"d96e2ef0907b07bb", x"38d7ad71f79c941b", x"36faae3aaa7666e5", x"80f131849002431c", x"aebeb3b1eddfd550", x"1f96ca0d06f8647f");
            when 27948794 => data <= (x"2fda600ce815cd95", x"74d3c22c0f7bd967", x"6b1fb46d312c9587", x"1f22c933114ad64e", x"636d3fdf6cd52241", x"5de20a0b609934a0", x"4b00e4065dc3fd54", x"daec0200c5f52c3a");
            when 17291935 => data <= (x"66043501d1808ded", x"12b166ac4e1f0f1a", x"d17c1e7a21d4a174", x"60ea550ec8e8bf55", x"885dfccea1251f7f", x"05a7e479eed70644", x"2f83df70c5fa94d0", x"413017b8e9379851");
            when 26684579 => data <= (x"36145ce9da8233a0", x"ec7b5183cbbb06ab", x"17d38c22b17e8ef3", x"b97306a7f99fad99", x"e936ed25e83b6c6f", x"db2f5296ea9445d5", x"0e1137e7258bbf9e", x"f8ee0f63eaa25814");
            when 2208598 => data <= (x"4fca32db66617117", x"7a445255e6b56284", x"4f02e06efa4a856a", x"d61657fa18668174", x"fca4354e91696065", x"3f7c4b90cda74619", x"c6971fd42098279e", x"329e2a0fbb250714");
            when 17593178 => data <= (x"a98cee1fe479ba07", x"ecc6847d047abc20", x"7faef717c6b21361", x"689f39975460e44f", x"2d2c22809d359a60", x"52142df2a32e8c65", x"3891bdf4abaa813a", x"c96d02deea9697ee");
            when 16227534 => data <= (x"48a80f3a5218b80e", x"4ac19bcdba23bcb4", x"f0950967a750ff3e", x"f35176bc56c4cd66", x"8c2ee495222fa97b", x"8255237a6f4bd2ca", x"1db7efc25e0fce35", x"d3124c853f5f9fed");
            when 33503733 => data <= (x"5ec4e585bb95400d", x"494e39099e1f38e3", x"833cbd75f2bed34a", x"a9195fa173a7eba1", x"a5e5880fe2b47368", x"42c9aee292cf919c", x"329efba1d6e15e74", x"64bc37e87271e4f3");
            when 7512865 => data <= (x"4f949c013a481881", x"9454794736d61d6d", x"58d2683cabfd9c88", x"53fb86a83c7f79b3", x"4a2c2c20194c7070", x"1af7ee14012e805e", x"8296e8d3bfda9599", x"c09693b3b0778c05");
            when 19763594 => data <= (x"d73df53e522f5ab1", x"2cc3fe061f51ac64", x"efab63a59f044a77", x"4591278c0c19a122", x"ae65c16304bbffd5", x"27089e8baec73b0b", x"343d0fc35c3da844", x"93c1e755916ccd47");
            when 1620265 => data <= (x"1adbc7eee0ba3e6c", x"6df52c1b17e26eb5", x"fd900c0fc8bd23dd", x"e242d35737857c8e", x"e0ec75baf26e303d", x"e800c9d96dde72f3", x"0eb6b665554c42be", x"1eb454f525545272");
            when 3207669 => data <= (x"6baf708525e4d230", x"f0e35a2ca22e3acf", x"36adab2582115a67", x"529f8890f4734151", x"cbb3c1deebbded21", x"02a44cd3f0be7818", x"046b7935d1f07052", x"c74189169ba712d6");
            when 20815751 => data <= (x"0f00846f83b63c4a", x"2f0410cf0864608c", x"a95e20bc5f38b8da", x"06160423163468c2", x"30b977da31c49069", x"f4141a02529bad29", x"10416c248297c0a9", x"5040ed627c89b406");
            when 7404675 => data <= (x"e691a71504304cfd", x"1d5037db17098343", x"4febff8b73ed0004", x"1e0cfc221f595a32", x"be4c0b6f66c4e181", x"5efdc262416fbb7d", x"f462447765abb6cb", x"d94456659aa733f8");
            when 8016876 => data <= (x"0fd6831dbda9ffd4", x"1f408dcfb3171928", x"bb128d553215cb7c", x"72d457eb23000e6e", x"8ee549c6081e683a", x"9244ab933820d127", x"c0e59561b4a62ba5", x"2b2949ababc500f5");
            when 32446036 => data <= (x"187cd4dd19849324", x"eb69918bc77ea1a3", x"38dd53242789da1c", x"61ac8d271605578e", x"52356892fbbeb181", x"a69937dd169ab43d", x"d041b2fb7c04c7fd", x"18191f4b8c197d5c");
            when 11676393 => data <= (x"ee44cf217ffde788", x"6f81295c2ab416a6", x"73f69be5d36f6454", x"707deb9bd2788078", x"455bf4da3ab0f577", x"8ee0cd5399d2540c", x"c07c902b919fe26b", x"6870ebdf9c16308c");
            when 10218681 => data <= (x"fb575bbc87819fe3", x"9615e4101cde1d69", x"c4f7867c5a904d2e", x"0acdd8d852749975", x"151f3d4418f74151", x"82ed49aba57fb3c7", x"04b5abb31c6e02d2", x"3001ce0ca83451a4");
            when 21810780 => data <= (x"817b10ffefb0c991", x"4322babcd6313af0", x"f7c4e08998e7b7b7", x"30a055bcab1b1261", x"a098796d1826174d", x"3a0141dc82f5c4c0", x"c920aa3b65602473", x"3537f5f9836074b5");
            when 7471571 => data <= (x"093d0f760773694d", x"fed6a20981b8f692", x"24a0d523323249cc", x"853c2044ffdb71e0", x"06544ee5c18ef34b", x"50b8c882c06b5738", x"2b5d14ec3c9b926b", x"6a1d29fd8d2eedd2");
            when 25034548 => data <= (x"7aaae4c105f46101", x"01825f366b9ef15b", x"37ba53defa1f3247", x"b9e9a7cdab41fd44", x"48a818f9049d738e", x"e666d908a48d40c7", x"0f5ff67c499c544b", x"29a41be71a4b3bc3");
            when 6461033 => data <= (x"713f883f2de9a21d", x"01f3c5592e01d592", x"360a8a27919b6754", x"bef0060e6c5fdb21", x"965d0e212f7e9ea7", x"466c28d8be23e762", x"2a653dbc012ad217", x"0ae300942e7dd949");
            when 29979698 => data <= (x"0e303652342ecd27", x"d60d6258199d0113", x"22c099f42108cf6b", x"f8ca55c88e8e4b93", x"113a246b27748cd8", x"35b9af61d79915b4", x"868a973906ca0932", x"ea49ad7c89644148");
            when 27466881 => data <= (x"c299022b51fc4e19", x"09da71b7b0d03f56", x"dd8f01d394eec23c", x"b20b340fda7cef96", x"c0bc81f67c178441", x"09d6b3471c853046", x"af4f4471f97a8b0d", x"2751cb7240bb144b");
            when 8088315 => data <= (x"2c3dd24ab651670b", x"2c79fd1a1703fc0c", x"7a81ab06c6366ed0", x"c9936a85c0db2d5e", x"7ba36b0dd9172cc4", x"c89dd398737f5a27", x"fa14c9d253b50be8", x"ad056184be771495");
            when 31814231 => data <= (x"97a347e2b0e8f4be", x"2a1a7a6b36b53d2c", x"92e459e07ce55272", x"baf7681b21e88df7", x"d5ba4f3dad8387a7", x"7799d4c63ff5cf14", x"e0e3aeae01bf2a0f", x"5dc214e359cdd318");
            when 26409581 => data <= (x"8376268e09112190", x"18d5be5826ea8f59", x"3e1f3240086d900e", x"0dda41ef9c965047", x"94ca74743ee905d3", x"51079ec35fa861d1", x"e699c511c85b9d37", x"aea98319361e22eb");
            when 8829531 => data <= (x"723e5040aca43533", x"4952b61efac3e43e", x"e56971e40b6bcce5", x"e96242bb3ddb2595", x"fbec2aca64193e84", x"d4fe0e39275abf47", x"16084a9b7ad52e54", x"deb48973c87ab19b");
            when 26804407 => data <= (x"f5ced70200a66ba5", x"2af45734242114b2", x"d2d0d25bfe9a515a", x"6da2b740238e90e1", x"d1494f527fa48413", x"07b961aa708d1649", x"f7fec512ed16a5fb", x"037efbd7d898c672");
            when 25570838 => data <= (x"03547aecf32bf69e", x"cbb18e13cf1e6475", x"01367df9ed6684cb", x"1031140545f01a49", x"35ace9144387fb12", x"f69b864aee1826a5", x"acda35c146869117", x"598395141d614a9c");
            when 9666564 => data <= (x"5830439faed34ead", x"1facb7ad695cbeda", x"dc7cb6e3588ea362", x"f36c9e0e47857fed", x"763d57008e68fc0e", x"2e9f640e314d438a", x"d4313055d378839e", x"b9952233746fc447");
            when 18804546 => data <= (x"8f2293cbf4c95b85", x"251601a2afd1ff33", x"298c57602a03db68", x"1a04268043b3aa32", x"ec6cb5c8da66a336", x"d2326cd4326be8c2", x"618e5c0446f92cb5", x"a1c8b24ad14c0000");
            when 6506813 => data <= (x"82cce66383fee783", x"37c7c368ceeb437f", x"a1b6e531e3dca519", x"11f307e2365a229d", x"5c40d91fd5a7ed89", x"207f1eda422805e9", x"f4563186e34fe1e8", x"176ab8a1ee9cdd15");
            when 17487264 => data <= (x"2221720408cd21b0", x"c2f0f1c8a605743c", x"e41114e4ac565c7f", x"33e2108ef6534cb5", x"61217a0d1c7c7713", x"50637826a7049a21", x"4bd857577a8f06c8", x"1bc95f2d6e29d2bd");
            when 7023066 => data <= (x"9438f8773538c72e", x"0c647762fcf4f4e1", x"0d97a58fa05780a0", x"3661c4f491490800", x"6ea9a109746b2eb6", x"fb152aa7c276213f", x"9395786f0afb23a4", x"3acfc3a5e5ee1809");
            when 19606650 => data <= (x"00b211d879ff30c0", x"dbb10feed7fbfe67", x"eb0f82739b3ed847", x"a8321c1f0e757ebb", x"ed9cf2587b6d5ccd", x"6edc91e12c55962c", x"137f0c023df39241", x"36ed89bdde0f7071");
            when 30574974 => data <= (x"4e41b61c8b7929a8", x"65e0b8823b71d0e6", x"e8b69bdd88cd40d5", x"54507be6c8aecccc", x"288a3a4b727ca782", x"a1d0538689bb7dec", x"50038722b88034fb", x"7340e4273b7a34bd");
            when 16144582 => data <= (x"a88c15293edeec6f", x"f5a9f09c3e4185de", x"57dcc9451905ea98", x"293a2c32653fb564", x"5915e5168136d4a6", x"6767e7b4f796d727", x"cac6742ab64c6aef", x"c222e6f8aef87e69");
            when 2459721 => data <= (x"0e2b599c02073132", x"68db7fbe57d86243", x"abf12a7168137324", x"1f23fb2f5b355ab1", x"bc6297e593e2b218", x"4a8a343cfb2a87f4", x"6fdfbfc7a8f12c90", x"1b79d36516f64adf");
            when 19897965 => data <= (x"61fb39319b3f831d", x"bf4c14f20eb556ef", x"a5873f188032f467", x"924543a47ed2a1d2", x"c1b20eefb610168d", x"5f061744c795a7f8", x"e7ed0c369b903408", x"ce01faac567d9262");
            when 25195147 => data <= (x"9a0a6230848d4123", x"790d89600a6a2e64", x"8937c3c441fbace2", x"5c1db489db90f318", x"40b19fca4419594b", x"db06a61c6f91e5e4", x"391951d6a674a512", x"d4f49cbbf36aab93");
            when 4643343 => data <= (x"7cbdee162c35c83c", x"a4835a7d3cdbddb4", x"98975c33b1bc7257", x"f7417e9684f8457c", x"d1680862ffa26de2", x"743d5028aa588a80", x"16f79ce8367ecee1", x"5dd0ef3162196eda");
            when 12882349 => data <= (x"1c9d9c8279ceea6f", x"b05e23fc7a687dc4", x"92a9e3cac60d3741", x"d8461bcf55bc3c6f", x"271f33de231ad52b", x"f4537f8ab6be76de", x"fca8c682f2cfafce", x"d5cf5ea0bd2a45cc");
            when 14734865 => data <= (x"09ea66f09dd24ce9", x"d39a3c3fca196dc7", x"357205270d1e401b", x"d6576c264bb418d0", x"afdc52c9ea02cd5c", x"710359df0988db44", x"592543016b08c1c0", x"3cf99c0ca5fd7874");
            when 24701500 => data <= (x"bc1f9315c532dd4f", x"f2602e44d446d20d", x"1400ab1cf9606182", x"b5296999232e70dc", x"83cbb381ed137522", x"56e9cf2eaf068724", x"bc73cab42e1f9dfd", x"b5684699a1f5a7d0");
            when 8999081 => data <= (x"bd56afb93029e98a", x"4a9b308aee30c992", x"66acb7ba4431d10f", x"de00bdc47f368275", x"8592ebb41a9627f1", x"5c04cfdc5742237d", x"70f0fc625c027d55", x"fca4079e68ab6f53");
            when 5612362 => data <= (x"7f263ca1d8d202a0", x"3fe63b1464ae4eda", x"1cdf841e0001e459", x"0c07bbda219d31cd", x"41b47cb8444ca939", x"b816683d242bd368", x"4afe6a6a639b21d7", x"228ce049735536ec");
            when 23118471 => data <= (x"8857453f689ac9da", x"9859d58276687c55", x"e8dca58e3b41ed59", x"72d69e9bdce7b177", x"6dc9d03f27d6de20", x"062f027d081978d0", x"6b56645263d83448", x"1d20ad52aca1e9f2");
            when 8433147 => data <= (x"dcd8146b5fe91ae9", x"094835c0b69927aa", x"74f6c9cc2b7cd89e", x"507bf184de046c60", x"3a7f67e501070c86", x"94ea895ad7ee37da", x"63ae82ca7c7e88bb", x"cbd7a468e17d3d7e");
            when 3533948 => data <= (x"bde91c6905811185", x"6530805e5d8d1e00", x"93ac2b20cf51c919", x"2685fef82ef3fd9d", x"a65c96eb7baa1e74", x"9285ba587696c612", x"808e80f7a9a20e59", x"c72b8186b8e5bb8f");
            when 9075953 => data <= (x"4c1eed9cf9bd5c39", x"da2200489392a684", x"bac46a1cb6aecaeb", x"d14b47c6bca10aaa", x"3b25a5dc4b44bc9a", x"fb2c6489bb96126d", x"c6fbf28a3e89b3d8", x"1961e90cab311efb");
            when 31438803 => data <= (x"d4f7540939e8cfeb", x"85026834473d7444", x"b0fd955f4d0f358a", x"4c647b74bcc89cba", x"3450367727fa079a", x"604211c6320dd7b1", x"6df1889ed1f1166a", x"11879460ce75ab7d");
            when 6019813 => data <= (x"5aab1cf9bd8f8315", x"72e55a4545e11811", x"9619995a2b5bd9e8", x"2fc4e6909b16a2fe", x"01d299c5530f3f5c", x"b7d7a4b72c8cfe5c", x"109d9b338206376b", x"a90d3d41d70d17ba");
            when 20741114 => data <= (x"532868385efd3721", x"e2978d2337fccaad", x"85949003ab213f41", x"b3447f580a9b8b4a", x"cb3eb26cad8c83ac", x"6eb7659c38cc79cf", x"5177eb540036dcd7", x"671f7d4a297c36e0");
            when 19932118 => data <= (x"858b92e76cd9ee6b", x"e8c216a9ae45c2f0", x"c2d9e7c3ab569b06", x"c84ab3ef140a6328", x"7e0f7bceb6bb935e", x"8b600feebfffcf50", x"9497d64246bc3898", x"ee490c5e00feddf5");
            when 22685449 => data <= (x"78b825708be0c3d5", x"de4ba465d0e3c449", x"6017094b28d7378c", x"03a59cd5fa478e5a", x"b80c5162b9a84ccd", x"ceecfbf0bfb6d367", x"12db5958991f7d02", x"ff30ea6bfa8805ee");
            when 13008924 => data <= (x"bf2fb0c7acaf317d", x"35296a071e0c849f", x"358f0c490e5dbc0c", x"c21a8e5020a8feff", x"c4d77a1e7e22af2e", x"2192bcf48d83ce7c", x"005ccef843ae819a", x"6fa0a9e5b4881b4d");
            when 5640131 => data <= (x"5618550a9351e349", x"b7cec9cbe6e5f102", x"f882a7bf7f0c427b", x"e3e42cdcd78dea28", x"0506c4e364dd7925", x"afbad76218f65490", x"b452a0a1885e1541", x"eb1cf98c70689b50");
            when 25382860 => data <= (x"63dd416568ff23a6", x"54e0328d9b0472cd", x"5ddb9275d06f6c57", x"cd2f218eb108dc8b", x"f459af2034754fe4", x"b4e5f60d2c83a30a", x"65444aabc6c39a81", x"eb4407e5304aa2a8");
            when 32803051 => data <= (x"b6e53dc84ff5e753", x"250c9957b276e8ce", x"83a9adc12f708a68", x"de152d1940741c0e", x"03617453524477fe", x"741ffe9f4f5751c5", x"6ef25e0dbde94ec8", x"513cc31be5343072");
            when 15469452 => data <= (x"4281d87099992ec0", x"9b0b61cc869a61c6", x"2250aa5521970971", x"35b407eb7337cb2c", x"e2406445a72be80d", x"b26ec69075f289fd", x"aef862bb523be0d7", x"6ecfa81c1dabc196");
            when 2394405 => data <= (x"53ecbba28c46b0c3", x"4cc619c0dbcab743", x"6a2855c8f0955629", x"195b67752e8036f5", x"3ff853eb51d34002", x"34319522dd9bdb4c", x"281febe7fd9ae5c1", x"a39d32d3aedeae0f");
            when 24478358 => data <= (x"c42cad01e224efc1", x"bba91e4f363b0e2f", x"4ef01db3d2dc8227", x"83492d38c255528b", x"3e1ca0681f16ceae", x"5133003dc8ecc936", x"5643f1693356683f", x"5acd67402867bca2");
            when 31125891 => data <= (x"92bf38dca367b61a", x"37b2e7f5e384748b", x"2d3a9f1dcfa3c53a", x"cf0b288a13c76de2", x"effadee1162e0b59", x"3ed42fe9288fe46a", x"43b8175e50b2c895", x"d8a7bed6109d39e4");
            when 21618800 => data <= (x"888b222627c5b2df", x"82edfbe810cb01fc", x"dc7bd02879a1d4aa", x"e5491ec0d44822d4", x"aa09c8a23b83ffe0", x"96d7f3d816ddc7d8", x"63dcea34936adc34", x"02e248557447b2fd");
            when 14614628 => data <= (x"3fba2904aa94f1bb", x"bddc8592bc826803", x"1d2ff84ee6a6d937", x"fc18597405dcbe97", x"2c0261a7ef1098c2", x"de8c3335c6e384e5", x"51e5f7fc932f356f", x"a71d930677af9c3e");
            when 18670221 => data <= (x"b9d41451c3b968b4", x"b6008a6c17a4db74", x"ab880f94671c78c3", x"13d5a605afd39d65", x"229f4ad1c7c7e89a", x"f0c6921e8c59c1ae", x"e46f4adf2631f3de", x"3bd53789b34a7f38");
            when 31180507 => data <= (x"28efc6749ddafb56", x"fad48ef07447c06b", x"14abecced4493908", x"c18bde6e3b7b4180", x"84ea8337a3741d16", x"24390060eae1c577", x"eba206a2b1892f8c", x"0d35b97d65f3d282");
            when 28516717 => data <= (x"cad72cd03be607a6", x"97fad72786e0a738", x"dda16c6b17a1da6f", x"3eede27873d17034", x"9f3395c34e0ea721", x"e48445f2efe2d680", x"601de0b50cfae9ee", x"aadb0b0b353ae02c");
            when 23395735 => data <= (x"ea085afea6505ea0", x"12df7c6f07a8d653", x"873ad6c8d64dfc06", x"298ed8d1f0b620c4", x"74ebd446cb80fd10", x"83e96a91142b507a", x"3f507d4f20cf7847", x"022e88265f28db5e");
            when 16673922 => data <= (x"0e8ebc386029e70d", x"4273cc144be2c904", x"06317473a77125d1", x"ddb4a68d30344856", x"d99d0d4823e29a48", x"e74cd58f11ce668b", x"da040b9ba7a91dcc", x"009a02b0208072b7");
            when 27525380 => data <= (x"b991e71f867b2a8f", x"d4315537ccc0281e", x"a4a954a3268eaee7", x"597ee69f64369986", x"36419d5a38d4fc6d", x"64f4a354b0043691", x"94b5e92c64d87cfd", x"58ee5ba668ad3bd2");
            when 11058323 => data <= (x"b98c73be21831757", x"b8ddd6ac870b1100", x"e23e41bc57466f3f", x"44097072417f24b1", x"b8c8ae53b4178625", x"016e4bc608912c36", x"d96a6982df151715", x"b904036c643b6563");
            when 10791233 => data <= (x"168c2e7baab49dab", x"e60899a9d8b67b94", x"7d91f24de43ff474", x"f26249a95f40d5ae", x"a32664d9965f9518", x"1a51c0ba666e5d70", x"8b2c4bd68d642199", x"82cec82bdd59d40b");
            when 1309031 => data <= (x"81f2c93bc2ab39b0", x"1d07251a80e7cd8f", x"0cf9516cdd8d008c", x"50482b5766114096", x"e74fd35f586fcd13", x"cbf543002d7b7e20", x"87721740bdb2ffe8", x"5dd6ff619316f701");
            when 28880243 => data <= (x"bc5e1e7f41273445", x"0d2f5bf43618e652", x"3d8abc4d9cf5b7c4", x"9696ba965dd79501", x"2c99ae54ba045d3e", x"d706c850e830e3d6", x"94bd79b7d87d648b", x"f5550d1ab2c96847");
            when 22054511 => data <= (x"201db8368d081074", x"69e87cccf48a3820", x"880a2197c657e8f7", x"8971e12a1bb7b4e9", x"c662d2bc969ddcc2", x"4f8aca22f2196a94", x"cabdc213e731bd98", x"58f4ab5d2c9a4dd9");
            when 14013561 => data <= (x"2be5d60a42c5c6db", x"b296115d0ce197f4", x"e8f3253a16579d0b", x"2b619aa9b0981e59", x"631d211b77cf0aca", x"d2c618fbcf08dd4a", x"d44e4855d742f8f1", x"da2bd557f5914e35");
            when 24999955 => data <= (x"9b3f6ad9c1040109", x"8225bcff37a027c8", x"7b3bd90b6c9100c9", x"156340cd43f2c1b6", x"42b1a126b79f6d7a", x"dad7fe2fa744cd02", x"df50865dede63598", x"a3d6297423aefe87");
            when 32915875 => data <= (x"76190fd048ba1076", x"c505ced5b4fbbb64", x"6d20a4555d867424", x"187996ab56315e80", x"4f9a260a884d699a", x"99da2dd922b51654", x"b4048cfeaeece29c", x"41e049fc6fe6d193");
            when 19588373 => data <= (x"bac3da5a3bd4bd1f", x"c4dc30e3032ee008", x"a7b387f2a36056d6", x"0fc3a7c0ca0ba0c8", x"1ce27e4c42ec8250", x"fe24a8b2bafce82a", x"d94173dc5d3d9ce4", x"8b746b319653b896");
            when 14716366 => data <= (x"6221e7429c9743b2", x"bcd9b7cb62f86243", x"2df681aec19b5906", x"81c726233de0d772", x"90d6d4b75abd4559", x"1dbed4a590cb4cb6", x"6c14c01427f3cb11", x"c792cd014f7deb6d");
            when 24443923 => data <= (x"7afcda8c8b11539a", x"ae819608f5d72d19", x"6ffa9b0262ff856a", x"81376b01a875588b", x"a66f05348db427e2", x"6104bb367110f232", x"08719d2472734a47", x"c3ad4858c202a838");
            when 15697533 => data <= (x"24b3f95f76c1e32a", x"423b9228c247f942", x"971df029c79e8529", x"eabcd381e1da0f13", x"2c1943563835753c", x"2bf0f8917afd195c", x"6e9c8d1c571d57c1", x"0b932d6582375fe2");
            when 17376696 => data <= (x"9762ff67aa0e085a", x"0dbe2cd52ffd1e34", x"afff989aa675b874", x"65f66676b43017ae", x"dab753c7a91b9643", x"74f715106295d280", x"a94dd068598b5994", x"c39841e0b616ffe4");
            when 26201693 => data <= (x"efb9f4e58edcdb12", x"bb848b7552405598", x"20af65454036f63b", x"8b65288c22c100c7", x"dd69402d94211f1d", x"814b766658b239f6", x"858d659b337efc53", x"739075419991ccf1");
            when 17363630 => data <= (x"6322546b11609c31", x"180862195574908b", x"e0e81dbed4a56859", x"465b756dc91ffaa7", x"854a388c01bbfd4b", x"af867fcf0627b75e", x"027fcb1229c1bce8", x"c7d474c4658134cb");
            when 20878970 => data <= (x"5f090bbb6ca1aa21", x"ccb06aa775b360f7", x"65062eef1b6da6e8", x"60fbc7692ba0ea5c", x"cf101cd275ff8c11", x"8072cbf3a45f169d", x"f36dc1bacd34f873", x"5c0d738e37810236");
            when 5881183 => data <= (x"7ab70427ea681c2f", x"875682edc6b252f0", x"9f859ee7c7b5c0c7", x"828feaa6ce6c57f9", x"857797d6a971b500", x"170a26761811be9c", x"38eeacd782fa627e", x"fbddac6541505fc4");
            when 24002842 => data <= (x"3146d471d98a5ce7", x"e821c39c0e70697f", x"349ce451deedd04a", x"7d21bf951f3698db", x"a3c7b6e476639c0e", x"a4dfa68bb180b0eb", x"c047003f14c0e7c3", x"afc3188262e24969");
            when 27561941 => data <= (x"d46415f9387b6ba4", x"3d7642052cf3f48b", x"2e430dd6c45db693", x"3717c1df4f54817e", x"41ce66a119212c4a", x"b98a8fda6a5ede6b", x"e6fb1616945e68bf", x"31137822f53e0f80");
            when 8042167 => data <= (x"035ead432461fdd0", x"002b93422eab03da", x"8e1f95e3f8d55ab2", x"9738dddea2003545", x"5594ab43c0f7d798", x"dfba46fb118c8411", x"46ce56867501b81d", x"e01f8146ec26c7b3");
            when 19025386 => data <= (x"2dbf82accd5ac2b0", x"7880d7ccb8abb250", x"33e5395a32996d8d", x"bf9eff2d26bf240d", x"96981658f2754531", x"c5563f21712cc946", x"d4be2e37a88c0249", x"7b989b8a8933a9f0");
            when 33007629 => data <= (x"bb94be93ca9047b3", x"69e1f371dfb1f12d", x"d02aac51a646ebda", x"598ca383f99fba3e", x"c0e7a1b8c57f97d4", x"b120ddaf755e3643", x"b5932518702415e1", x"af85561ee77466e2");
            when 29186425 => data <= (x"a2050f19a2d222c7", x"e226df72df928252", x"db6c71a82f88a5ab", x"24ccda0019fb66ad", x"66f08489ec77983a", x"85843a6528b113aa", x"446b12f198dbf301", x"2b0253c825f86047");
            when 30668589 => data <= (x"9e517091b69abff1", x"51dbf76098281028", x"887c8d8a4a496971", x"0ebeb09431c9f691", x"6b3423f603ccb61d", x"c0e5e62ae4925a82", x"1d2bb6459076befe", x"4f8368a9de09cc28");
            when 5425164 => data <= (x"af09d6d667fcf6ea", x"1da0db15282ba03b", x"675e839eab151d7e", x"3aa7ba4f92dd9dc5", x"31eb39b757ca4439", x"38f975947ee9a315", x"254b18703274224c", x"7073427f60b8e4d9");
            when 15655951 => data <= (x"c7cbb2321d794612", x"a81b367e42ff2649", x"c523cd617e598985", x"df8912eb9aa1e3e0", x"329b062a02e4f331", x"39942a14ed7a6f70", x"03d988ffcba794c0", x"0c94139f349531ad");
            when 8242799 => data <= (x"92192a5596b64748", x"d2e6f031f79066ae", x"cd4cc83229b2d77d", x"4e828214e91a56fb", x"a717ba9c532fd577", x"44703e267498d072", x"0157b8dca8bb3ee0", x"c33fec9689470be8");
            when 1005373 => data <= (x"e50a915e5fc51868", x"3c20cd2b8b239652", x"431a03b8616ab1af", x"56207c38cf48f374", x"7f7ebaf114fba09b", x"2ea32312e80364fb", x"de14e1adda602c41", x"4032431174c91872");
            when 27940323 => data <= (x"aabd5852e6159463", x"7bd5a7b79f5c1bb9", x"f752639062c45019", x"ba405dd07da45437", x"ee27084f53285fd0", x"bf43cbccb4bfd0a2", x"3257df577d142bd7", x"a4329f3e4b1abbaa");
            when 9629715 => data <= (x"abd586a726badb91", x"f6e5c5c6f0461086", x"9fcf0cf0c0512a2a", x"ce63b3dbf4fd42ee", x"d41501a098a07bc3", x"3fab77a9256fb720", x"e7dd71dce654032f", x"58242d5b384a262a");
            when 32906213 => data <= (x"41d3ff24f0d36aaf", x"5176206114d436a8", x"4199dd7e2c2e0487", x"a19c97af9dec686e", x"b0c2f55a03f01e9b", x"5a2072bded892dbb", x"72339b8ea30abfa7", x"72e848b809a43cb0");
            when 16185690 => data <= (x"b17f18a76d7ff402", x"a834624df724d1a5", x"a6f3408e41ca57ca", x"054b0a94625591b1", x"1f50501305f624d8", x"353db9df3386efb0", x"0e3001fa5f93e13d", x"49580e72af019531");
            when 33184223 => data <= (x"cb0f7679d2c19127", x"42e38db718cbcf12", x"e0a54370a0f8bb63", x"9807d2cefdb7ddde", x"e6ca805921e26c47", x"fc21af12613fb587", x"0fc85ea594278f4b", x"a7d9f3014ff4c3e6");
            when 20615254 => data <= (x"aebb156c302f6fdd", x"dcb37e4155225fcc", x"b33f08a1c1255efe", x"7816844dcc36ae14", x"a386acf5b0e5c05e", x"ecff73fd5fb6988e", x"d5e58454f65a5d8e", x"3f4af10bc88180b7");
            when 11578703 => data <= (x"5135c1f5eba8a173", x"5030ef8cd7e09504", x"87ba7083e3f22b44", x"c1e42bb7ce27ac0d", x"242b174030acfaac", x"687be6b68e0b90a9", x"1511a6a38a5f8201", x"b70f12954783bfac");
            when 28560914 => data <= (x"d79bc12066b92370", x"1d2ede9910939723", x"3a5315402de4cbce", x"94c30c11e7048d62", x"e10eadc0cc52d84a", x"c537a7edb87aba45", x"bf4c7487e884857b", x"c38a9d26e52f74cb");
            when 7607875 => data <= (x"99f0963243082e22", x"4c212bd7a50747ce", x"6444e404faf10990", x"ba8cd72fb89faad8", x"ed5847a141ae73a6", x"e5fea8349dd06e45", x"484f77426306ba40", x"9109b17d3f4caf82");
            when 2578550 => data <= (x"ee12353a3843f2b6", x"85561d912d904e5c", x"577af193ca091c86", x"3bac8805090ce82f", x"2b4f35022e33a3ad", x"8a52a90d17094591", x"ce1a8329a4480f33", x"9cca4b24a66e21a4");
            when 26130661 => data <= (x"88b7211ea0b13105", x"9fec01c99f6b7b63", x"ff05b855d0ccf8b0", x"e01d85725d41d18c", x"aaab47ddbbfb34f2", x"70ed9c0e0dbf504c", x"33fbfbcf69316a9d", x"60925f7bb7a04926");
            when 12178790 => data <= (x"629f7c042ab15dff", x"6746b433676bda2c", x"53e1a13b99d14870", x"3bf0f1ace3278189", x"2e97b958567ac3d7", x"d62edc2eaba12183", x"009118a170d78341", x"0847d9f5e1dd60f4");
            when 4180395 => data <= (x"5112970f090b54bc", x"dd5bea0e6b1b07a0", x"84b14e14871750ee", x"fa4f7818349571db", x"d968bf65e3d5a799", x"813646c2f53a1dbc", x"df5d08d8f8751cf9", x"10333d9af63025f5");
            when 3818321 => data <= (x"d6865fc555c9c860", x"285b5b317c006fed", x"27ab1df6db7699ef", x"07666334cf91327c", x"4fa2f69b649a3e91", x"1091b5a0a481df83", x"ad0f3f337af871eb", x"2e17927a21c83951");
            when 33896119 => data <= (x"4aacda7dfb9e90f8", x"ee70a315faf32713", x"413a9100f563b940", x"b3f82726e92aafec", x"cb7cd0b2db959dbb", x"862e0e7920762c21", x"47eb5728c637d3ba", x"74ca63e924248e2b");
            when 20292107 => data <= (x"5d942a750d36f05f", x"6d46742158a05dd3", x"1598b8ca418a0f28", x"bce84037ab38fafa", x"fe39062a2de029bf", x"db0705c9d7bf10eb", x"79915666bcad8073", x"f0c8393c287d7c03");
            when 12650701 => data <= (x"1fe31af4ad3dc19a", x"a66471d1e2d42b3a", x"523cd438e373cb55", x"ff7181d746bba984", x"bd30c08fb4a44cfd", x"cdd80c9e249c4135", x"cf9547c31460d818", x"3999df5807e40084");
            when 30129480 => data <= (x"be7290c60b38ac3f", x"b3b885da89154f04", x"024994eeb0f25156", x"fa8cddfb43ed4d7b", x"c4ebf6f921cf7274", x"d14dcdd80af71822", x"502a34504ce787fb", x"52bc1cc5eb9d52f9");
            when 806567 => data <= (x"78fc3e8a35ee3750", x"747b757476e30daf", x"a208dc5f589baaef", x"99510c1bfc469ff0", x"ff084984ab002e5a", x"d7200338fedbbbae", x"e168e57fd7d02e37", x"3648aceafe98c4bc");
            when 7946850 => data <= (x"a5acd95ea58fbb47", x"02adac7bf37200f2", x"68ebc129a1d61b67", x"7d0c417a738fba1c", x"123df78fd8b4b24f", x"4473e1229b9e57c1", x"2a23f3e1d1e5d706", x"f41e65c3aed83680");
            when 5053919 => data <= (x"d3eb4450c89e40b5", x"e6540458b6683b35", x"7ce808df1ba22eb6", x"0679a7e9e650f0a2", x"7a660e4a961fcc58", x"3edfcedb922d03f0", x"eb0600943a1a2b26", x"925b3659e7c83b3c");
            when 10248235 => data <= (x"2a70eeca280504ca", x"8afea734d96def49", x"5f150855424700ed", x"bfe6126c63a20896", x"35538500b8671d51", x"f85879b5bce8e790", x"e724b34d04c0b081", x"cff40951251e7769");
            when 7881921 => data <= (x"9a8f933f0b8e4e22", x"c18541f7e3dd9fb7", x"d5a7e6cfcea05ec1", x"d85b9cbbdc9700fe", x"22197551cabc04cc", x"4c886b122fd218b0", x"9b9f4b0b04da6c92", x"4bd36b560927597d");
            when 6937646 => data <= (x"8338fbf19d89aeb2", x"3ac25bbb0402398a", x"0e194068a647963f", x"f7cef4d0db1c374b", x"99a68915123d09df", x"550fa05a209cb1d6", x"38be5492ef45853f", x"f3b42907c7abf50d");
            when 26681581 => data <= (x"7d2eaef1acedd059", x"04470dcac826208b", x"c4e6df0db03af212", x"4fbd6a67218000fd", x"c05392131a3121bc", x"f880d3498fef2df7", x"6549e3078de45889", x"8138dbe66c4e41e8");
            when 7625785 => data <= (x"0303f51726b13191", x"cb4d6458b5fb4b87", x"e463da15a0fb7b5d", x"21d40a7d2c108be9", x"88ab88fbea5c3ca1", x"5e6abf698a10626f", x"811faa0e4d31c4f6", x"79dc2ce06aace2d5");
            when 9261118 => data <= (x"d97087cbf93b86b1", x"4b2cef8ffb82c241", x"53a66e5efc24dfd9", x"1751abf1323c1ed2", x"87602d1bd2dbc0a5", x"6084d7843148cabb", x"e004308d0199ff21", x"9aac0fa8c170823a");
            when 18300094 => data <= (x"6db807fcecb3911c", x"765f7255c2a17de4", x"9ecf0776e1979747", x"c336dddb715b9125", x"573e9724e87347f6", x"b5aa1c9706064928", x"6ac91a499cbd7606", x"1f062c168c668f04");
            when 4888257 => data <= (x"2193653438f780c1", x"464a18630356769a", x"da41b893d9853d67", x"a3b5c7569f7be16c", x"0ab5e6d43a2b1784", x"c9f56e0131731379", x"fe1bbd90d23089a2", x"658bedcb85a72cfa");
            when 10484333 => data <= (x"4d34851e2fb4ac2b", x"2689a37199bbae2b", x"29801af819d79e89", x"c3d444c44621b3f5", x"35e7adf400327ad5", x"3c3f2872a6ff699d", x"48ee72426402a48e", x"e6ccaa2972a85ef0");
            when 8099829 => data <= (x"b7758651d8d1c7ec", x"90a78292eb30dd8e", x"7e1b9f16958eb1f9", x"607b24eb2ff85ae7", x"499757241e73a5cb", x"fb5f5f07bed5b26b", x"e7f4f9e5cfc7d3ea", x"a72358e120125c9a");
            when 8076185 => data <= (x"e751758e70469637", x"dd2f70263fc67dee", x"ae6682c3a3664d12", x"3676d827121f24b4", x"eb5f1ef189214777", x"a33a5eef658ed422", x"725716cea5892efe", x"840fd6e50bdeb8eb");
            when 20798630 => data <= (x"6c0fe016b3b6e6b7", x"ea8f4073bd0f8e9f", x"194e39d28a73ed7f", x"882a6b1e2aaecdfa", x"3a000cb93da2a986", x"632e44fbeebce738", x"78e540996c935856", x"4bb2b2a2577351ec");
            when 10850000 => data <= (x"dba89ab7ddd1dbce", x"b7269e3a337fb0c5", x"807827fdee78efc9", x"d94f863d7f68a2c3", x"5164a1d31f6e7cd6", x"d65213675efa319e", x"24b3b7aa2f05997a", x"90434a3e8f5fb81c");
            when 33047323 => data <= (x"b1b5dabaf60b8f72", x"4deb279edcc47775", x"003aea8880b4a046", x"373cc96730888375", x"c84a051cd95b5cc9", x"8d1fcf9b54859e89", x"efff10760bbf6e77", x"2e0baae3be448699");
            when 12883363 => data <= (x"927f26d76d118c5e", x"c5757781b7a2266a", x"8442f90336cbc533", x"69d9279aee675a54", x"34139a8610196c6a", x"7721b68ba2d70d6b", x"9533cb9e4be19ce5", x"6bb1d16bce9cec4f");
            when 18152352 => data <= (x"1620208a70b7469d", x"d3eba9707bb27676", x"ae4bf9bdaabcab0f", x"01816f0195370fe3", x"091f959034812e65", x"414349eb20d32a96", x"312b13c7dfec42ef", x"fc46a4439bac2302");
            when 26387290 => data <= (x"2c32b40a67f8c453", x"1a7598297543fd6b", x"56953a2484d0c307", x"5ab2e60353a1b60d", x"f173c442f8e3ed01", x"0eb73b39a47c76ad", x"fc43ab63e03ae3b9", x"939837587b54966a");
            when 25132464 => data <= (x"2ca351004ae5432b", x"f63fad09e01fb2be", x"635423cd05bdfb0e", x"066dd9a8ffbd6f6a", x"0bea4f123a5223d2", x"0bc457a410c8d340", x"931eda300c486f6c", x"a5111fbbf727a82f");
            when 15797196 => data <= (x"de6297a1fe075b89", x"848ca8e883fe949b", x"3d2c78202f2dda41", x"4a0feec315885939", x"f96bc503416b3045", x"eeddf4cceffb1412", x"fc13460ccf5c0c77", x"c85f51b5952dc834");
            when 3583307 => data <= (x"199178c6b4b099ad", x"12e44ffbea691296", x"7ffe2f0f91ceafd5", x"629910490f75467d", x"9037739fd093ebde", x"693344372926310f", x"74d0db249ff7f53a", x"52874e44b4bbd84a");
            when 3132604 => data <= (x"c2ff9e4d55a101b0", x"069c9e0c30348e7a", x"3b852363f16fc801", x"c8946796404c4ff4", x"f5b5a569a4e8e588", x"3ee4423a4b0137f7", x"8a2ca830b846f34c", x"3d1d68301c4a7898");
            when 22695132 => data <= (x"8db4a2fd9fb91442", x"1cf032890d9bdfae", x"46d002b4823dfb65", x"3ede14d2221cca52", x"b08a043352a871f0", x"8e276eab9a96e5d5", x"c63e2a07d3b38bfb", x"c87f83aacecbe57c");
            when 8026425 => data <= (x"249f9e09bbece655", x"a23ee6e4bd1281b9", x"bbdf82421137a8ac", x"7ab83e9cced3f7db", x"2fd7de08c9890e8d", x"f9f885ab0dc5f606", x"40b704810af44c87", x"0be859e66ce61c91");
            when 21942612 => data <= (x"f63f32675f7ec021", x"fe3006b4ee853794", x"ba5548ae60c213ff", x"cb55912363692da2", x"8043581f507d8022", x"ab69c54fae9fcf14", x"a0371907175bc150", x"c0bf5e7191594002");
            when 5453489 => data <= (x"54a8f8cd01bbef1a", x"adaf4345584a2b79", x"61b4046656f000e4", x"7c065efa8c04ba20", x"559ae80db2f84e04", x"cd8c2a2014b9f452", x"b6b5ccd294612307", x"572fd426832d2041");
            when 25960882 => data <= (x"0582ef980334c035", x"9844669530a87d3d", x"826c1c7b88a91b78", x"5f01fff9a0c270ec", x"afa470f107d89881", x"ca6fc9be6e748388", x"9877636a92556a59", x"89f77a5faaacc059");
            when 8531921 => data <= (x"cbf7d4df78d47f46", x"3765be9466f29e98", x"456577047ee9e622", x"e4882397a279d184", x"227f1c3503fa3cbb", x"cd527ce18eb9cac7", x"49d160500c41568f", x"52531e885f034b40");
            when 12257474 => data <= (x"54dbe2e15ae789b7", x"bdbb119632444c78", x"4945db7f3a5aea9d", x"7943592be7b2fbe4", x"cab1aedf554e36f4", x"1d26affa24003321", x"c639dea1fe69ac33", x"9465461d2956ab57");
            when 3885069 => data <= (x"a0a4739f7a0ea9ba", x"ccb945773fd13bd0", x"a54d4c966c6d76b9", x"612bd68b47224d91", x"6ce6d7d56abe773b", x"cdd9ca7754c77969", x"78456139e856ffd1", x"28a9d3df5c95e9d0");
            when 27887500 => data <= (x"c82707454ae80d04", x"f1f6acc18eee6162", x"349a6813574cdc33", x"6ce0698164d44ff0", x"fc4011abd2dff2e7", x"8b5d89d38647d4f6", x"94171bf437c330d9", x"6b3852d96f2a99d0");
            when 2985018 => data <= (x"2460211862151094", x"bfc72d7e821a0f86", x"3fa4318dfc893cee", x"169ead1e86cc0e52", x"93c68c3353f099cd", x"7e12d232d2b780af", x"c7ca331ab4b2098d", x"5542699a6d84e6e0");
            when 10505142 => data <= (x"43e8a8a7320fefe2", x"e30b7932288943f0", x"448f6f4ed35afad1", x"094d9ec31ffce9db", x"a03742c883b50fbb", x"6bdcedd4db4ac648", x"1a9f7f2aa7c07d06", x"7e793ae735ddeb63");
            when 14992087 => data <= (x"5ecfe84e8dc421e0", x"4a66dbffe7eb2b35", x"84aa8f510755ec75", x"d6b425f03dc24470", x"0436f3e1d3813bf2", x"6bc503af9a653164", x"aa560f5c586ec8ea", x"eb07b0cdc13582c3");
            when 19548099 => data <= (x"740a3923bfd43dc9", x"d31ef75578694df8", x"c6717744d360d7be", x"2f3c56c26703f043", x"f47dbf2f339ebdfa", x"914e67addacea1b9", x"3cf5e8c119d0d45c", x"ba9d6ba73ddd5878");
            when 7069168 => data <= (x"8128254100804874", x"720c9f61131ab8a0", x"0c00034145589e52", x"f0205d8361f09302", x"17f8c91d7b8dae07", x"90d623c0be3cc7c4", x"9198e1aefdb790f5", x"ee4a4d30d764463c");
            when 9331052 => data <= (x"1258174f5f7cd072", x"6c16160a753ebfc8", x"3f3f5cac748c78ce", x"68855e3005e14b22", x"9da0b3c09ba9d09c", x"f8a5cfab924a9d02", x"fd082e8e83a2d946", x"1e60ff6223ba8566");
            when 28817751 => data <= (x"fd4029d8763d03b1", x"9acf6e1e7d627c94", x"0f1bc96cb39b1593", x"2b51efd81a64300e", x"6ea6aa4513841e98", x"122e159f6ccf2263", x"c73b8dc464db69f6", x"905a0af612b1b73f");
            when 27781069 => data <= (x"864b331d18c01ed5", x"d1dcc9651e77af5f", x"e8473825b31a24c0", x"63774051f1373582", x"e0d7e6f074001f79", x"84269c7743617fd7", x"53d56fa02b9d2aa9", x"c31aeae92b93f0be");
            when 33418024 => data <= (x"0fd7e39a72603a07", x"6139caf3030c0269", x"0d4ca4c48feae5b8", x"f6cbf798ba73d693", x"629ebf3062a994fb", x"efe7fb4037d7bae8", x"da00d362f03fcb43", x"312fa675bedae352");
            when 18706199 => data <= (x"a28868f9ccef1d3e", x"29f09eb921b28f64", x"4ca699720a71cbcb", x"754460363e9254a1", x"05400be28e537fd7", x"dd71e54ac3a524f5", x"1a71a3024c37fa2b", x"08ff4a45b4748791");
            when 25341091 => data <= (x"3104ec5d0257daf9", x"80708cbf56dd894e", x"9a53fe0697b63140", x"17538bee45642162", x"abad56d634f779b1", x"9099994caa7cc3a6", x"ac9d165bb5b04fa7", x"b226e9ba40254450");
            when 21299224 => data <= (x"d0d5148a93f2c53c", x"e7a22d6fa0e052b8", x"f3fc28026b39ded4", x"6655fc25f6787fc3", x"d1545180e1901617", x"1d6b0c2b728358b8", x"71dd9d754992ce6b", x"103dd14a67784ad5");
            when 2827611 => data <= (x"25c1c1abe4dae730", x"3eaf6da9608985ad", x"97903f01a079c49b", x"eabcd8750a412973", x"9fcd0d9b1d97519f", x"16332a702893cb1b", x"1ef97ac7340e7083", x"cea42cb6991115be");
            when 23345614 => data <= (x"effa36875d04a604", x"f692c7850adec49e", x"dadda109d390f6d8", x"fe51967d70e30db5", x"121228044ad5221c", x"4a742381560674d4", x"4c843f1cadfbbfac", x"37ee2f64d009c395");
            when 18471817 => data <= (x"c1d963e29c4a1b24", x"789a05774b8651e0", x"5f0d626aa8d35c53", x"405f5f70f0f4775d", x"47ba3e6a51d5d67a", x"95f995661eccb08a", x"54392b82f6f90799", x"1b4815a6345d4784");
            when 28110830 => data <= (x"45ae78170fedd838", x"4f9b304be576dd81", x"1e6105adc0a6519c", x"3f7e6e722f9c82d5", x"e9c88da5aa9d7277", x"c08318179ec9fa41", x"2bebf73a1d82cc5f", x"bbc1a27186aca64d");
            when 11716464 => data <= (x"e314b0e9167fab80", x"518507991bf30110", x"e93ce5b1b4e55a23", x"c2c1fc0b71906778", x"21a7903b8d449d57", x"443b79195165c4d3", x"4c0b651fdbdbae83", x"df51daf47d41ab5a");
            when 16206351 => data <= (x"7b3b5aa7fbdf5e8a", x"9d11975fc4bd03d4", x"a518bd0e12c56665", x"5b619d2cc7acb4f4", x"caf396fac1a9bec5", x"045e65410fe0b27a", x"2fdc14f6d42061a0", x"a1d92ac0a9197b8e");
            when 7426766 => data <= (x"304be01770f07df3", x"7360d18e3fd67cea", x"28f7aaf3650d6f93", x"278787ad524cd9bc", x"900621d54109b0f6", x"cd75c80576072f51", x"44a265c793d7c8ee", x"8bb4da66c953068b");
            when 28714448 => data <= (x"12f5a244dc336932", x"c1ba91c66a7e1b14", x"640de12b304d7f13", x"1e1ef2ee8768c8a3", x"d83ed5ad50cc74f5", x"7efaa0f8c5f59736", x"b529cdb43175d014", x"850b03d05f9aa626");
            when 23327415 => data <= (x"ff57a6c079600d23", x"fa781db9c2b91267", x"7f3dbd1eedd7489f", x"538ec59a2f24a5f7", x"027a2a7a03f39709", x"4111e6ef69a71086", x"b0a905b40276a6da", x"27fcd6c25955ed0a");
            when 24913490 => data <= (x"273abdeb567792a3", x"226718a8e479fe1c", x"4133af7832cadc84", x"177256038dc2813c", x"ecb48f71616d597b", x"349be0b92c5a539a", x"a1f6601257d907c2", x"dc223d217363a329");
            when 11360756 => data <= (x"1e50501318ac4ee5", x"1957be43ce701428", x"0f1115d88e32aa5e", x"09159c2f21c97188", x"401b0361e2a13e92", x"17e6f1eefca70ae3", x"6596507493f4d2b9", x"efce74f27643219b");
            when 25293335 => data <= (x"1122b3092f46c9de", x"edfa45a419e85204", x"f420e680757f51ca", x"4c907850fbdc69f7", x"5467f15dd531c72d", x"fba358293f36f7c4", x"c1f1b2ad27edb57c", x"67e95a0620b1976a");
            when 14119623 => data <= (x"1a6fe57f2ac289d6", x"e100cc92bc662998", x"fde84371a4f19f9c", x"7585d207ad407195", x"4302995e2de2380b", x"f418e6752f6a2f99", x"9ae8834d82aa949e", x"a3649f7400613c87");
            when 3086893 => data <= (x"7d465503042f2c3b", x"9b63e6455a99f1e4", x"8b49ab1ae02cfcee", x"fc4fa92cbc303e0f", x"3a546140f73d5c89", x"fcde0fcb3e7fd414", x"7c8ba6588b8b8cfe", x"c570a586ddccb003");
            when 24403831 => data <= (x"40a04246252512c9", x"b968a7cb11fa54ce", x"a3d2d9e4d01871ca", x"1bdac19d0014d0a3", x"8e801e8f9f64bff1", x"cae25ad900bcb5a9", x"38fd3440cfd3996e", x"ef4a21c66f792e1b");
            when 4494625 => data <= (x"9c3cbf258f110298", x"835a6107274bac6b", x"0f3ce29edb68b4b1", x"c5c8e5dde01d987d", x"73f0c6409a7abf17", x"33a7b9927eecde5e", x"e5c70cb72d3ed6d0", x"020041d5d93fc26a");
            when 12428775 => data <= (x"a9bce453df86852c", x"2529ad58e5b5d766", x"f191810b127fe492", x"7490c1c19488ce34", x"595409dcc403ad86", x"9e411cba4ffd77bf", x"2c54f7f463e20107", x"d839db457c62581e");
            when 4366413 => data <= (x"541279e9f984523a", x"57e445442dc8a313", x"0b8beed6c8b3c5c7", x"3ae216b2f954c43b", x"73c1e26409d9a8f2", x"0ebd356c50a5a702", x"75e9e2839bec2504", x"2c091452c1ac5201");
            when 22310233 => data <= (x"b3b393e2a149ce02", x"8a00446ec2b1dfc3", x"1754da7ff2fe7d72", x"f4c13f2cca74a0ea", x"c2b24fc293c1ae56", x"22896f880ac38fe1", x"1e380369e027fa9c", x"694ecbf17b41ee55");
            when 17545588 => data <= (x"c6a7acad7aa28934", x"aa3bcd1deb1d9be1", x"d48c4258c14b861b", x"20ce8c9f1977b204", x"06535c1abefcb39d", x"2c72080fa3cf8f6d", x"85784880139196bb", x"062b2b0691cad8d8");
            when 15258837 => data <= (x"1bf369911438db63", x"573b2c85c0e1bf36", x"8dd43459ef95eacc", x"a13c7f19bbe097e3", x"4d9578e969a65319", x"da715a8279f30ec3", x"1ab7b75dcdd52d2b", x"8404be130580501a");
            when 18706694 => data <= (x"96fb24bd62ef7f0d", x"2de98260de3f4c16", x"7e2db17ce5f21bb1", x"5475e64b3c0b9caf", x"14d1774fbebb69af", x"fafce6e02fbe0bd9", x"8ca61469aa12411e", x"761ffa7af6acc644");
            when 23097731 => data <= (x"bd4b5335f11b5717", x"2021a87c2886fa86", x"eddd8b99b88e0023", x"43a72c6b34627e6a", x"d6f2b83462a99350", x"39c949a0159a2bf6", x"de927b362489ebbe", x"61d7c2ff13535401");
            when 13550050 => data <= (x"cfc4e7e4448517ba", x"c8c3786b7f5b2a2d", x"888133136481820b", x"813794d9657d6434", x"9e9b2cd6a6fc7ad9", x"084240c212551dc6", x"cb79922bd3f0adcd", x"e660e55e83ac3179");
            when 32557827 => data <= (x"00292cb105bb59c0", x"9d528b715cc05dfe", x"86c228ae614f8dd1", x"f34a8fb35de18aee", x"c10d04a19b39c06e", x"d76dcdf211178545", x"6133c87f46082f64", x"cf1397835bb73148");
            when 16744886 => data <= (x"1430911599bfda07", x"3b8f9ba8f5366895", x"0b3fd12a25ba14d0", x"369d0a68750bb22f", x"a3c4e2240cc4ac50", x"3384970ad6f96e09", x"22e92785d76f928c", x"aaf18b08be07c806");
            when 6989600 => data <= (x"12492db03ffeca99", x"b79a0735952c5397", x"82efb2e8721d686b", x"13ae1e3ef9ff5722", x"51707ecd287f2c6c", x"2aba13daeadd5676", x"1df75a6f75026ec5", x"b2d36becdf8c65b7");
            when 5775296 => data <= (x"93d62c6534ea0504", x"be3045021f269976", x"cb60e85b727abead", x"cc67582ce60f10aa", x"430d051ce26b01c5", x"98e478a762dd0196", x"c0fec0bab76bf0b3", x"38a3fc54e79072bb");
            when 14171496 => data <= (x"d92c2f80312dbb8e", x"c6d5ed66376cd21e", x"b569f12a1b3dd827", x"3e5ed79da65ed4eb", x"07bda92ff852f4f2", x"c4a2164abb193a23", x"75b3eb1d27bf9dee", x"f4c20b8fe8cb8ebc");
            when 32237584 => data <= (x"1ef08a2b704ce403", x"95b2137eb549d69d", x"b28208007eed490b", x"50cdf4050c6b9b05", x"52baf2b3ed6bc36c", x"0dc15c28d2c9f6f8", x"66fba3af8a186903", x"24a6ccf4d06e6cf4");
            when 2569487 => data <= (x"da29c35bac532689", x"14c275999ee2c9ea", x"8d7cc5819f1489f0", x"39e8b3829cc37731", x"6a7ab9a940623313", x"1c8f4e7959dce8c0", x"c4d95102fe6b92e5", x"f361d014790919e5");
            when 29043879 => data <= (x"42aaec2f0fb94629", x"1c44073dbde7b804", x"b3ca78bf0fd80c09", x"783bdb8907a38704", x"66f646b0e4b60da3", x"eb7808498ce15033", x"cd7b1499b98b01de", x"1ca63c07a347ae8a");
            when 3414236 => data <= (x"ee57ea154719b0eb", x"911bd6b6c4020a6b", x"82d0906df94031c5", x"3b3ab89c4a0e4027", x"2395b477bbfabb66", x"c224856ac4bd23bb", x"411d041c96498c37", x"af5ec232fefc82d3");
            when 25439970 => data <= (x"cfe5bf484bc996e3", x"55860235c5d85939", x"177c9de75d397b8e", x"aa75282bceaa8de1", x"d9d9285f81e8e583", x"8db50c19b906bac1", x"e3d369defdb6f991", x"b13882c580ccc052");
            when 12887077 => data <= (x"629debff50b86299", x"31c424d3cf17e865", x"9305598d47f9aeb2", x"3f455f7e23e0ce2c", x"95f236caca7fb232", x"5f73fbb8a9e5f7d0", x"24491efc3140f829", x"7962a521f6345841");
            when 28874285 => data <= (x"6800573596e27625", x"9295a0bb089648fd", x"b84f8d0253063caf", x"7633924224cbbb0a", x"9a05076c58b1c10c", x"0238183778a529f7", x"e7419730b79fa6b1", x"a039e80f36fba37b");
            when 16778025 => data <= (x"a4c2b0ae38cd38ca", x"19a5052a44d56076", x"a4145ffd67fb9023", x"40f1f2b81b6efc1c", x"e2f9a597569a8ac1", x"c837aad1da05af39", x"92070092949cda7b", x"a469d21935529d6a");
            when 19846595 => data <= (x"23f7e146c2d9fd1d", x"cbc33dda6151575e", x"01ddac3cd8320271", x"1d52c2afdf0d3c71", x"351df71413fa27de", x"8603b28a235ec035", x"a2c2661d8d5965c2", x"9e6b3f948a8a2503");
            when 6326261 => data <= (x"dc85095bcd789280", x"8d7e5e8c581d0d2d", x"455778a7a4fc8e01", x"440fa1c57b4d995c", x"19e35064cd657ce2", x"44f85aad01120cb6", x"4aa2fd5132be4c71", x"a531a0586e9684bb");
            when 6402214 => data <= (x"dfb2a5c34be859ac", x"5f6814777d585af9", x"6fb0282316ce9da0", x"bde8d1d37e3f91f2", x"179f88016a7f403d", x"cd91355b231cc60d", x"271a69dde7a74044", x"f6dfc24474d40a4f");
            when 26463917 => data <= (x"15e54def8c9c350b", x"57608065c5d2e5e1", x"1e9ecc0e01f5160f", x"ed6b86a88b95a674", x"9479c4abf5cb6d1e", x"bad37fb2ac441c13", x"f7001e8b6280d675", x"f49f200f3ff59058");
            when 25411108 => data <= (x"6d28af2fe9296a7d", x"70f62c90d9204282", x"39a23598cb0b727b", x"bb1f93548cd69014", x"8d87a05db546fef5", x"0377883af47bb3be", x"f185e5ef7124ccf9", x"8b98cc00f96f5710");
            when 4443799 => data <= (x"03a6b1cfa523e15e", x"eeb5cbbd7ea36b83", x"fc14aa4c109b9b74", x"385176fdc47b78af", x"a6094382a9212a35", x"afebf7a0e9c4756b", x"31cbfe4ff6903b71", x"23991097344ad71d");
            when 31988766 => data <= (x"6183f117f7de633f", x"65a7214e753776e3", x"5bd2d9a5f72d5bc3", x"9e3991c4c4870368", x"f4fea124d2a59f5b", x"037e8565b019bf32", x"394472dfe2792f52", x"af31a5ddab035cea");
            when 501294 => data <= (x"b93b55deafc0b1c5", x"a5c07f0bb0a86cdc", x"125acfdaadb58280", x"733a5be1167244fb", x"b0ca3ae6667d7f6b", x"fb5c9176d40a2299", x"d9fd2d6d836167d7", x"69dff58255611755");
            when 4209791 => data <= (x"60e54e197594e27d", x"91f36e9108f8adc1", x"229eefff1ad2514f", x"e948c281e54bd7e8", x"f82223cd22989746", x"d4434fe253d262a0", x"334ef62539ab2ddf", x"80c55d920d750f36");
            when 32713099 => data <= (x"026ab3d1b7883ae7", x"4f14ecba98f3fec1", x"0800a3276879d5e0", x"3181966780474ff6", x"5ce06f8c569f509d", x"72803a97a33e7d70", x"5037d1ac8024e7b4", x"0d2f05837206575d");
            when 21539665 => data <= (x"1b7e09c6aed36754", x"6067aa44ab8f2b57", x"86478d0f1ecd9a36", x"7ba8d9c9c7cb680a", x"fd5717e36e3cf126", x"2583b7209e3d6dca", x"be65ed9029774034", x"f4da33e05c6c3757");
            when 5886924 => data <= (x"f27e1755905f0d33", x"5f5d3a1fc7d85016", x"a421f88e71419ab1", x"5a6c6f6f635eeafc", x"928a1a4b55f50e2d", x"c0358f8f79c1c5aa", x"9454c2fcb1a7d29d", x"567dc75212b62e09");
            when 30047792 => data <= (x"028891ed7ed31ea2", x"f5b148184659f8b3", x"359e1f41cf451ce1", x"54e86c41fa8b4fd0", x"ae8b3d88e02caf5d", x"b7721eaf5821796d", x"b3705ba26ed9bbac", x"6d6bd4e4a0faa636");
            when 1685851 => data <= (x"0e423f50b83e08e5", x"19502228514a94d4", x"0bc0d05f0a0c4e41", x"d3725d815d790e85", x"03c1f39e03bfb7e6", x"c5c81644146d2944", x"3ca583dc58f6740a", x"3e085f5d6e67b5d3");
            when 9491466 => data <= (x"4618dfca382f7df7", x"3b7d2afc88eb69c6", x"16ca7e913eaebc1b", x"e7b2bbe31449c51a", x"a01f715a6076542f", x"42560188e1eea05c", x"6c89668624698455", x"01cd2b0c26695d28");
            when 11608804 => data <= (x"7a0c78eae4f9f1d6", x"b8378f42aaaa415f", x"9f4c41296baf5756", x"4a80903f3afc9fcc", x"a63faefcc2b81d81", x"2a300d26c338687a", x"dd644f9172798837", x"9b4455791641544f");
            when 8871405 => data <= (x"f5a6986947124479", x"c1c44c408f338894", x"0f20408ea2803add", x"275420672e9390c8", x"b696575d19bab133", x"96c135a121eb1a77", x"4fcf0d7161dad9c4", x"cc7598472dfdc062");
            when 6257888 => data <= (x"e35e5e6d0c836aab", x"98e75380d4ce2d96", x"0d0223d0d2833e97", x"e56305fbbe7be8a1", x"a858d1bb90fde5ee", x"67332d9c3806543c", x"02ec6c8df1bc4fc9", x"0e80fb08cd839cbf");
            when 13107040 => data <= (x"d858b1e3cff45e98", x"d2bd4a6f010ecfd1", x"02da3b9a2c4b8b9a", x"cf1415da66f23426", x"e4010cc8a9a4e8c9", x"6814465b5f6afd40", x"dc2bbb8914433385", x"3d4260caf464c0b2");
            when 30852270 => data <= (x"0fe82d47433574d5", x"253cea618ea1599f", x"626df78d6e561d25", x"5abf9b8adde2d47a", x"d193d18d8f808a03", x"734f8817e8b636a0", x"b2a730953ae41d25", x"a0052994a0da3f42");
            when 4831437 => data <= (x"a8be044faead081c", x"c04a0460ffb9f10e", x"a2d858d9dca509eb", x"f0230f8e28100bc2", x"0639475a324e7961", x"3d3c8ac15f668465", x"85181085013e57a6", x"fb4397c719371d77");
            when 13211248 => data <= (x"79b580456874dc2d", x"0bc4df7c9562e4e0", x"10eae0cbc371ce62", x"108cac663888fb02", x"f121664999b20b90", x"1c1d898555f86f80", x"264bae71d46297a3", x"9b27d106fadfb765");
            when 31212846 => data <= (x"8ff00f00b04b22e2", x"1afe58857d5d9950", x"815690b2e32eeee5", x"cd4622cfcc236c2d", x"dd8a27fa5fe8a977", x"84ad454ed323f7c8", x"9f044810d85726ef", x"bb2688da9dcd2796");
            when 4998989 => data <= (x"24040b8df52c0731", x"c1e475fbe6d2fa06", x"1a46463306d210b3", x"f516fbbee2484b41", x"48eec78a7e4788cc", x"653785d4cd6f996c", x"0282be51dfb49b7a", x"8be71553358dd8fc");
            when 8402284 => data <= (x"515962700875d169", x"7a97e835cde4347f", x"7c032baaee5fc1a1", x"97928495e1c8a451", x"abed16ef3528fa51", x"eac7293c9bbbedb1", x"f3350f5c903c049a", x"4fe405bd10927067");
            when 31736251 => data <= (x"5b044f45f3edb8f0", x"4d245fb94aa627c0", x"2902219f68b9dde3", x"98ed69fa03ceaa50", x"7fd8a253c8b45330", x"cc06d1c0fd0dbf6f", x"be4903b8af400cff", x"5367d1bc8c8d9a86");
            when 28832395 => data <= (x"2e61b89fdd3e5b69", x"1b761f6144ef391b", x"ef907a48092bc5db", x"b828429139bbea1c", x"d454db2d9e7fa448", x"04ae960779c81b80", x"d010ba057cdbdf90", x"5141b6adc3729472");
            when 1435799 => data <= (x"0173101fbd0e1d69", x"ef88cc8c3064a1a9", x"2fc29e71310b9738", x"1d5f522269dbc3ca", x"79307868840e8db3", x"71ccfd726981d986", x"4f34326c111a468e", x"e88dd45f343c9456");
            when 11178840 => data <= (x"b6ed8670534aa943", x"5ad94c0f1075744d", x"043ef3c8881af4d3", x"4bfd570877345b63", x"19ae198df2f38184", x"3dd8af6b13917191", x"189c13a775a11411", x"a2d1a26a574b4499");
            when 19345305 => data <= (x"baa63f40c7667505", x"7c1669b98c381c75", x"9a6125996e4a3e9f", x"aa2a645e586f4d47", x"d74fe214415969ac", x"489c3c30d1881592", x"a3aa7a46b4d78a04", x"347e20c63e9341c5");
            when 24429135 => data <= (x"32d65e8cfecef187", x"730a42f335c4099f", x"076acfad1d8dc1f4", x"3d12f9836459244d", x"d0df7d3a1fcb6157", x"86830356e5081f38", x"70a41f06ddb6b77f", x"a095649969b13900");
            when 30425902 => data <= (x"d8a7d30369432203", x"1d1cf5080a8d8e8f", x"6bcc736bd4664128", x"509d8152b3363fff", x"3e1444688396d7ee", x"00b96ac3bf68c202", x"4a3f9ad016f061e3", x"f1bcb94ee6da3665");
            when 19900337 => data <= (x"3be0589b9037f545", x"5adefdcfaea73f0b", x"f2dfc34069b3f914", x"f743d903b30c2eb1", x"d4c1ed0f6340b132", x"cba6a53fc265dbc1", x"8b61493738c7e5d3", x"48c086f31395c926");
            when 29817974 => data <= (x"267f47b04b42ecb1", x"5b9146593622a5fd", x"72846e1e82391fdc", x"3b189e7cf851004a", x"e9c5f81ff0b5710b", x"68b42b56d7a85f12", x"6b14f5f7350d1542", x"0fa1450d5bbab005");
            when 28914633 => data <= (x"efc332634bb03b61", x"c1e37732af8dce69", x"7d2914adbdc63b4b", x"a850dd63fe6971c1", x"b4a2f08b9db583e7", x"7dab9e2ce202fe0f", x"2920cb44f5fa07a8", x"31bb1e3facf3a90d");
            when 13781922 => data <= (x"9c1aa107175d6d4b", x"09fca7482cfd954d", x"dcb667448fb6f69a", x"042e6010bc21a4a6", x"38c8c4e412e23a94", x"1f8402256df4554b", x"9a03601f5091cb14", x"16062654ef75b8c8");
            when 9279082 => data <= (x"2d4bcc2203392bd4", x"920084d8b1195483", x"18ab9c39658a2aee", x"a2ddaaa1ab78012a", x"029cd6d3ef31452a", x"4e31b6eae1d8758f", x"56cc6e13346c94ac", x"056de9d409db49c0");
            when 16389975 => data <= (x"5dba6709d155d472", x"a7f80f2fea21b1d9", x"92cb1eaab35145ad", x"0231d02c43b87f42", x"3e8f40062625e464", x"b854e939502c43b3", x"6b5952a644629e43", x"2cfb9c0a28b8d3d2");
            when 31203901 => data <= (x"08c621fc8983a5f6", x"d80377c635b2ef98", x"661b7f1d13e1cef0", x"1065a6b7453d4187", x"acbf80d9b0a2b106", x"e82bfabcb3eafd75", x"dd2843cf86eff452", x"47758ae15ef902c7");
            when 29403751 => data <= (x"27e9ede6b84b0bb6", x"aa100d798b5ff008", x"c52e2a01b51d8b0d", x"c8f3aabf7f039d77", x"85211557077afde1", x"5741ed71deb7daa3", x"b5e125d58349ac45", x"e62b967e04d90b1a");
            when 8411392 => data <= (x"f7c3523cae22897e", x"9a00b79e4a4d34d4", x"1f40e1a25f47c3f1", x"fa6f360e0d8e8e83", x"9575eb8b975930e7", x"632fc711fbad7e1d", x"5539ab1bbf9f3c30", x"241e4ee2b9b56abf");
            when 2117254 => data <= (x"e8919f37c5b9a6c4", x"a30d81bf3b3bc79a", x"8ff15b72916c95ec", x"31dd7b71eb26173d", x"7ae4dda70ba6a1fe", x"27810162500e54cb", x"888e5ed2f50a2b41", x"79246c3f3a298ceb");
            when 7551240 => data <= (x"100b47dc18d7ca22", x"05e41d93bbc11f8d", x"e5bc18dc54760e73", x"2dbb5c342b8a88ff", x"40a659b890becb2a", x"c4486805b6cc8a90", x"6105bf71a9525937", x"b930ff05cd887fcd");
            when 7471460 => data <= (x"4d3d62c42df8c1ad", x"52ed94da61c838b2", x"e82bb3e16283a3a5", x"af69457423fe1ea0", x"5df7b04005f131ca", x"b79a0c1e93018c4b", x"4bd9c4aee95cb3d0", x"17f14b2b92305b7c");
            when 2357252 => data <= (x"0d334e654bb192d9", x"3c42b4e68c707aac", x"3674e860c8fd17fd", x"a0887288e2ac87aa", x"d0db74edaffa088d", x"2caeae8fdaf7ab14", x"66461908617f2313", x"ba2fe91a7b34b119");
            when 2439123 => data <= (x"d93d9722e652f777", x"13fb93829cd3a86f", x"6f7d88543b97b534", x"fa318be621bf90dd", x"0016793da0300c1d", x"3920c7d94cae5c55", x"7f075fcf44677add", x"8b17c69046d35cb2");
            when 19800094 => data <= (x"9407d8abda2547d0", x"cae5cb13615a3076", x"4a749260efc38a36", x"937c0828d6d5730d", x"1e90a82b514e1c48", x"86d1b3f216cb8261", x"77463f479f2c8810", x"f563cc8dfde34909");
            when 11324346 => data <= (x"ebfce456a2e9f706", x"320f41bdc1392556", x"9e9d62b8e3f15e5a", x"2f854545787d34b8", x"c571050ba14df417", x"2d2cff52a3f5f2b1", x"41b7abd6edf7b195", x"aa2a7d84851905c3");
            when 5240840 => data <= (x"f8ec8e660e615e22", x"78a3dcb886b18e62", x"508ea094a2eb6a86", x"5cb6b5153d4be030", x"be3bae3f6a5bb745", x"2b1508a1e07747c2", x"59a22c634c6a751a", x"276c89ac17601f52");
            when 18306814 => data <= (x"081705b57f693ab8", x"39c1a601fea3ef13", x"d90f6ffc09f00c81", x"2a85b8fa0d625d8e", x"0616f131b7a1ab77", x"3fa3e0c35cd67106", x"104ee6ec91b7a6ef", x"6fa3e6a3f0349735");
            when 32081824 => data <= (x"180f46760a6272cb", x"e574095855ae5524", x"c2a249b030e02499", x"0cbc777e2b38f79c", x"567689d6242f83ed", x"4bd489596d3ab14b", x"3ba3527235a6d1a7", x"b7fcf8f317ece948");
            when 21832672 => data <= (x"96c37a9a1e174c09", x"f97f8eda958fc24c", x"fc300cb099289bb9", x"b8c508bc8088e064", x"b4ae15ae91ef2bf7", x"195b9cc169c50a87", x"15bdfcc69473f37b", x"2f69b501c1e57c28");
            when 7258141 => data <= (x"3fefafa905585368", x"fdd9b8c22e577eb2", x"efea8bd9a48abdac", x"630d6cfc5838d657", x"84b066bd00a307cd", x"be2ea6ebd8236877", x"d26824430f3109ac", x"eadf9de884ed790c");
            when 5811178 => data <= (x"4c036657d9fd3abb", x"f774964f10ad84a4", x"3c9e767ff6092d0c", x"8e375993cc9f1ac6", x"846f62a3521f834c", x"a1863407273b2cac", x"5c7a5c35d53ed170", x"d8427b2b96187a0e");
            when 26303300 => data <= (x"8676dfaf89d6132e", x"55d913f8be3f75ba", x"8502579a3699f210", x"bcc9061df424f752", x"b6a84134a240be73", x"95856ecc024e983a", x"c98760c74251699c", x"1eb8722be06b59c0");
            when 28677037 => data <= (x"9c4c0fc9f54aa86d", x"a32d84ba44d5b9fc", x"c7e2366bccc4b471", x"f92d23e3b4de3410", x"55a374f98c46ffd8", x"fb29131af99c4550", x"2e98ce4f2389f4cf", x"f172ccda96265b55");
            when 18806380 => data <= (x"d0554d8f3d4dbe7e", x"8f3cea4048aa411b", x"fbb317ede94140ab", x"f2cdc3f2d1c97fec", x"3b1aa8c281366b8a", x"ee0e0a22dd8c3ae7", x"6f241ec93a7a308a", x"111d66dcd6ab5c8d");
            when 12426355 => data <= (x"46d679d6e1282548", x"f4b43a9405347938", x"c174920851085598", x"c6306c4bc7dd0490", x"a6f66a1bdad29a6e", x"225d4d97d6f2623d", x"b53632382692cc93", x"a776ea85b7409b0c");
            when 16698266 => data <= (x"381c2ee0f3356356", x"72a7097d45faaf51", x"df6d7e0b8db99ca0", x"79a40e8b6f09defb", x"65166a8ab9196c8b", x"1544e28cf3962991", x"e59a9480c7c444c6", x"4106e5ef5aa9023d");
            when 4187972 => data <= (x"436bc24dc548d2b2", x"6f378f4c085b8b85", x"cfd99b31dd3f882d", x"0325bac5df9e96bc", x"f332e3fb6a6dda75", x"f7a1026d51beab0c", x"1c42150b2ffbbb62", x"487385a9873bcb63");
            when 13469398 => data <= (x"d0d00c136d649d72", x"ce115089662f60dd", x"460b59bcd80abd84", x"0f8d1ab13575b295", x"87e8aea7aad1a751", x"4b33b1f46f820185", x"6ef7bf26f9fa2a21", x"29733137b42f0664");
            when 3025402 => data <= (x"9feb311246710197", x"107cb3c8e6630bc9", x"889118c09c4fc7a7", x"01dfbdac312568fb", x"d943dd05e276709a", x"103c9fd3a7018bf7", x"fc64e4ac4801b892", x"7c72d2dc0526f52a");
            when 25570437 => data <= (x"241f1c14ef7151d2", x"24ccb790f3dfb237", x"e0db62298a1f3549", x"c7dba3412649d48c", x"6ba31d3c2e6ddc29", x"14151630bf478a3a", x"722711341edd79f7", x"b3e85e7484fdf4a7");
            when 2264802 => data <= (x"f73f3fd8fe14d01d", x"77b22aed6ad01f69", x"23019c5a362ef60c", x"b54d7ddcbf4f2143", x"6cbbd25cce0bf51a", x"3dcfea1230a9b975", x"56d2a62ab82e70a0", x"2c1768dc230f476c");
            when 19949805 => data <= (x"a1e06956d25ca54b", x"e3c61361823adb9d", x"e3c64bc5523fe83e", x"e1d1313edf070bf8", x"364c957fe4b3f361", x"35fd1a8ca02b3dcb", x"79049e2ea6946543", x"78bef89f77274b29");
            when 5538710 => data <= (x"518d493ffe118229", x"11da2cb2ccfcc4fe", x"97ba62b8d390df89", x"0ad64e57af83df07", x"3d68a092442c07d4", x"2662857eb9ea04a0", x"232463a96d7d74f7", x"f06853c1229e5f39");
            when 10065018 => data <= (x"be2a1278159ccce7", x"24b83b3b3bf29cb7", x"0c3c296a9bd9387e", x"ce454e0977542ca9", x"c9738cb7993db577", x"ad26ed4f73ccead0", x"50771f5d02729306", x"94330b1d1ba66562");
            when 4203702 => data <= (x"7971b0048cb63af9", x"9d383458d68aefda", x"7bd8ea9b4a3dc757", x"6181e14306eabf50", x"b60c109a689a1d77", x"6e228cf3a7d3a964", x"1b10b9743f192994", x"b1a42361ac14326a");
            when 6660483 => data <= (x"91160ac75807193d", x"291d3d00618c570c", x"4bed6fac7d79b7c9", x"d6618e847e2d6f1d", x"e01be482d1f3282f", x"b342c70e197a5d92", x"6cc9db7951f57e24", x"07f5c602b0159033");
            when 5350936 => data <= (x"92d162f2b43bb870", x"da3b6bf48182957c", x"eccf11d51052dcdb", x"e1d0f078d4613dd7", x"563f604ad708046b", x"00cf62f1efa2cd5c", x"9951ce5390872cba", x"1af953e601573efa");
            when 3893824 => data <= (x"2e32743369b4b86d", x"422743bb3fdfce1c", x"3c4793dccc5fe209", x"01d43d2339c4ecda", x"df601f56c1b68a54", x"f3e57b8a451a21b1", x"5f073612c90205ee", x"14ec24d149684482");
            when 13360946 => data <= (x"e2136cb0b9400088", x"c1b0bbd7899a0eb8", x"f004e7d38da886c4", x"991f81eff77f4138", x"0448cdcd4f44728a", x"b3f589725975b9f1", x"3bc4c4cb3fbecf3a", x"fe74deef3b9bc37c");
            when 28849435 => data <= (x"7ac99e3f2fbcd03a", x"566933276fbadf56", x"84c0ed5193b6154a", x"bcfee3e8882bd4cb", x"33a624258f7df612", x"20eae7565a2ecb44", x"a794738ac0890d6c", x"d02e2e9f555efba9");
            when 2677161 => data <= (x"13f010e5a2a61935", x"331fa8cc4611402d", x"57f4153810d23e94", x"2b36a4cedb026fe3", x"58f2f9b22e3d9dd4", x"b444628880fcc8d4", x"ba0d647e38cc04d7", x"edf9afcf8ec9a542");
            when 28695693 => data <= (x"3af8453ffc6b794f", x"0256e40e44eab78d", x"9d7ff9686458e2fb", x"a6eec864e05088da", x"9db2755329a9f698", x"525e4d33330aa546", x"5342852afb869884", x"e43b0b9c3db39ec2");
            when 29716586 => data <= (x"620a50b84a080e67", x"bce2fab563b2ff36", x"ff41d85e2f004cd0", x"a971f242fa2de4bc", x"30834d10d2603753", x"2319e7ec06f7fb59", x"76aaee0b29cdad67", x"f7d710989bea45b8");
            when 17955508 => data <= (x"e86aa15809730207", x"18606c2da25d346c", x"5217d0bb63c36c3c", x"b3ee23531c428487", x"5265a08a41a67b4d", x"328d71ff91bbd561", x"7808d2678c5da63b", x"506ecba190287d74");
            when 8830847 => data <= (x"005c5ad839ebf9f7", x"67b8fe0fc159e83d", x"84c1f74661a325ae", x"cba979f8a449dbac", x"9f540352d96254e5", x"9311e66ef7ad3d85", x"88918083bc606a70", x"a49ea33babafa2e4");
            when 17462405 => data <= (x"2231f07a913c9d9b", x"1f80f13155f896d3", x"5bc7f9abf9acafa8", x"67d1ae6698da4e6c", x"5172c0f3457d3d98", x"a6078ad385f6196a", x"ae045f8d6b4ae5d2", x"0f1914a3c07f82b9");
            when 30262350 => data <= (x"4c509b9b517befa3", x"89406edb87bc3522", x"519adc8cc0f34379", x"8f1ffdb634240f97", x"da489c1f9e0a0b18", x"0b7ab9c831524c9f", x"6d42f0bf137a45c6", x"e8f3de6397ab5f39");
            when 4471364 => data <= (x"d99fe7fd620f1a96", x"7a9bc0c2ba4757ef", x"91cda65b730a93e5", x"1c2be5d5019eaf28", x"c278e32220ba5ea1", x"990fe439a0892abf", x"5ac9a4a1608e50a5", x"d6d0b2430fe5e563");
            when 6272962 => data <= (x"7de8b4f748ee1ce3", x"0879669a2de050f3", x"f75446e1af1593e5", x"2d0829f451ca4f32", x"5f006c5893eca59a", x"1aeb1cc9aad39018", x"7854e0fac7344827", x"915552de557f692b");
            when 30947788 => data <= (x"1dd17c1d9bbd6947", x"4c06e8c816c0694c", x"958c9a636808eeed", x"44dcd18b0098ece8", x"fd1d694bb7494027", x"170f2fda8dac7bbd", x"fb70d27d21ca8fcb", x"c8c0be4ba8281906");
            when 25231545 => data <= (x"66e930c517bdb148", x"0004b0ad8095aa26", x"6daac7430dac2a04", x"a35eb28fa57956f3", x"a8c3da37d6363ad3", x"a7d5a231afc45acf", x"67f7a1e92120ee41", x"1bebe0a8998bee9b");
            when 12215015 => data <= (x"f55dd5a7c69e1aec", x"6fc20d99e46c00d0", x"e553f9363eb230c6", x"b1dc825ec8ffd3aa", x"9244ee64dadfee03", x"5a240c85ee0f3da7", x"6789da0cd3429e51", x"f92557069c73688c");
            when 10263643 => data <= (x"9eece1c2eb062993", x"8e9e5b2287d5ff0b", x"01f15e68b2a0db7a", x"434ba2bdc700240b", x"a6bb86f8f1b37c67", x"c2c1e23696b53581", x"8f373ef0fcf70ad2", x"c963048760782500");
            when 13382245 => data <= (x"f850b3fdecba21c5", x"3c865068aacd56fd", x"0459375835dbea03", x"364139fb70294acc", x"9f202a8afade6789", x"e9108d40332f156f", x"3b39edf706c4f644", x"0fb87f9af62b7455");
            when 8875128 => data <= (x"1e1b00ff2b2a6cb1", x"7d1d1a856a61b426", x"ecc324cfc6eaac05", x"e86c715a77085588", x"c70ba154c50f7c06", x"198fe913547117fa", x"4da927cf19ff3d2b", x"2f62fa03c0f1665a");
            when 7580458 => data <= (x"f21a6b61a8958b9d", x"4b5d8617dba4be40", x"3959aad25924841c", x"c42c9f1260a2e1e8", x"5d524d26d6dfdf1e", x"a850128db15a2190", x"34f1c8b728fc4079", x"39c1142958f17b66");
            when 8029355 => data <= (x"0f7019dfbd522456", x"057a359339280beb", x"6c7ba391a0e801b9", x"d3559e57bf8aedaf", x"0b9145b6d81632ed", x"608de1a811aba64f", x"9002b16d331985e0", x"9268d6eb9d010250");
            when 12493101 => data <= (x"e337e61a91a77b43", x"6127b928cf26000c", x"1a80239ef71e7b63", x"dc9d3fb1044c8380", x"8a543c1fa3af6d67", x"77558de6972c9f09", x"486213a5c6234f68", x"d5ed0618e3a63c6f");
            when 10254450 => data <= (x"30c39b84a548dfe1", x"5df4685d7d9a8e0d", x"7a29722968ecac59", x"a37017b6c9fa77a7", x"8908193dd1604029", x"0a70ba51f9465629", x"697c3e9d0f171802", x"455e164b2dd766bb");
            when 13778843 => data <= (x"dd94a563c089e053", x"f2d798f20a98e6be", x"d00b24259ff4708f", x"a9b189f42148d9f6", x"36b086dc1a9a131f", x"ac3525525079143e", x"b9e61b6c3a3e6c93", x"7fba9ff31abdec02");
            when 5703935 => data <= (x"d74024c7c1b7ab61", x"463e221d8a2c5dc7", x"86bd20bcddfdc664", x"547b02283a526023", x"59390339db0e5f0d", x"f586cb422c426d5f", x"072e65255e942f34", x"f7a5612bf34f00c2");
            when 786661 => data <= (x"f970430d2b63e3fe", x"fc549459218bf8cb", x"bc06c9575fbd9433", x"a86d41dbfe7966f9", x"17d17c3b6a0d33fa", x"d86601791c2be492", x"52e20bb8fbd96416", x"846dc0746120964a");
            when 24920736 => data <= (x"904b5eb137f4f59e", x"3977e24ad71b8bf3", x"6fe429168291d270", x"7cb2fec7962bccd6", x"508685d6cadfbe80", x"871e2610335a6884", x"e94eeee621c6d3c2", x"385a4f70c55cfe94");
            when 25936657 => data <= (x"560179c78e3f69e4", x"a2aab4026a50e5b3", x"5a46f40ddea205db", x"7d22b69ae5d87c07", x"e484e79cdaff38bc", x"b3f9713e2599c544", x"850c52abf5d86f90", x"d243f3343d35e65d");
            when 23644353 => data <= (x"0dd51baab4c41ea6", x"d282b6de0d78c867", x"bb94e16472ace325", x"19563e1156f6b5e1", x"5f5c4c3f2e657846", x"6343bf018a80a77b", x"4c39224ea264f1a9", x"252b2bda3fec1957");
            when 24516633 => data <= (x"02539cebeac60bf8", x"4b457ad8e42e1865", x"4bf386e6f75e9ac1", x"465f7e4084f021c0", x"ef38297cd986ef02", x"d5e18563227edaa3", x"a2c83989ee370ba6", x"0b099a56156343c7");
            when 1346048 => data <= (x"2c7db56d4406dc2e", x"dbf826b07fd2b5d3", x"e557ff6727e6eff7", x"c705d1d0e58b7f02", x"b10566e84dc8e855", x"6da4c0f1db29b961", x"54e65ccae54581a1", x"bc42097dcab4a68e");
            when 25652770 => data <= (x"111b7c72410f20b4", x"87e4b36207939517", x"d6ba8fd1336931d4", x"b0e01d641d707ef3", x"6881d4eb96804952", x"79d83d9b71ab3a4a", x"414223b2071559f8", x"aa179e7feeb2a4c3");
            when 33010052 => data <= (x"d87e3c4ac714329f", x"f8b0a7dcff5cc21e", x"886dd5ff256005b1", x"dee812c2a02fefdd", x"7079b859557514cf", x"72272b4a11054f3d", x"acb51f7d2d0b5a16", x"b3ebf335fdcaba12");
            when 26969812 => data <= (x"f1ed65b0b1eab800", x"c0f97c9014e2e413", x"1073b80c0cf97048", x"86fbdceba74e2ea0", x"5680465999386e02", x"caf7a86eec4c0951", x"89048634fab50ad3", x"665f81bb0a29e68d");
            when 8975390 => data <= (x"77b66bad459c4b72", x"386a3c01d7c1610c", x"1dcf8be667f73a45", x"4d3ae8b354b94c32", x"2066a68dc1f7fb50", x"2316806a9ab80b35", x"28f8c4b7aee2e368", x"619e8bad8c10bbb8");
            when 32752226 => data <= (x"caa6bd6d3ef668df", x"23ce4753f7071064", x"d3814a2fc5450350", x"b84ea15ec90c2bba", x"435dbd571795f595", x"44f3ae4ee1ca2e03", x"64a7c575cb7f47ea", x"cc8658f6bda56f89");
            when 16245071 => data <= (x"60edc0024c72a1e1", x"f8adf7911b97044a", x"1ca47e44bf009990", x"fb8a119aeea8dd42", x"10d47e3561b23015", x"a194348c47e2b75f", x"e8d6ae1d16cfb390", x"ebdcc0fc1965e712");
            when 28210841 => data <= (x"4579468ec484388e", x"bef4b77adb0d6f63", x"5e5d436f5d11d13c", x"402fd33cdc9c9505", x"8dfbebfb3555c99e", x"bd7e264cefa45b06", x"4211d48f60b754cf", x"caf8e9b47c19939f");
            when 9034382 => data <= (x"26863de66682a53b", x"4283215715245fdd", x"ebab9cb44f312609", x"bf582e532bc6c2b0", x"71a93e899449de00", x"3c2b2bf249c0e747", x"53e6bf5941b488e7", x"28971af87c1e9d21");
            when 24098537 => data <= (x"33c9ad8bd25df3b0", x"8ddf947e7b675987", x"b66af37050dcf808", x"7f0686981350c7bd", x"006751e08d1cf0e2", x"fc02dd4e84a94762", x"9493a76f8c80770c", x"a59cce3b7d7e248a");
            when 26059918 => data <= (x"cd7148f9c854b627", x"16155a0081485e7e", x"91678b5b4fea0f71", x"74813c4934a900f9", x"f030997e02e625c4", x"faa6b9bed6219355", x"614f38023b0684d2", x"f0ecb43bcbfd1d5e");
            when 14799638 => data <= (x"4dcd71d7b52c4400", x"97bbe778d78d3663", x"343ba4c79f3f2f23", x"3904adcadad447e8", x"0acb5e76a39971af", x"10283be313f7875c", x"19cb417e0eb97da9", x"826da15128c232ef");
            when 18225192 => data <= (x"7d70603d123386a9", x"3559dced1faef285", x"e9a6a89a0f78c5e0", x"40179c6fab885761", x"a02d363cd4d79be2", x"952608055ffc9c75", x"fe49fc6592ca345e", x"d8e4057550c8f610");
            when 8181330 => data <= (x"f24d843a6ccfe1ca", x"258ae860171a21f5", x"56532a06677714dc", x"f17d61089f834959", x"1f8765632ed6fcda", x"4d480bfcd27b82bc", x"0b14b68fca154bb2", x"9513e0de9efc334f");
            when 20775042 => data <= (x"a0fff62a45d83d02", x"2f9ce19c0c698b06", x"ed095c003404f121", x"398c933e17659949", x"9fd77e22e3a93819", x"a44a338138a758b1", x"6fe612d26d0f650a", x"b5efd2df2e4ed58b");
            when 31521035 => data <= (x"e2fb0949aba4974e", x"7e5d0345228b97da", x"7b39349fdbee9b7c", x"8034bc01e4e68dc5", x"b9d2a9ce9202b993", x"d1ec2a8ef9940352", x"a5fd142683373edf", x"e92492eec87061fc");
            when 19017676 => data <= (x"2ab11dc0498162c9", x"15febede1c2b7af6", x"9f20ce5fabdc870a", x"296472ee3edfc3fd", x"0b09be4f1dcecf96", x"a9f6efc586b39d96", x"ab391b094af87b9a", x"2eeb7c8f6f1939c7");
            when 3341657 => data <= (x"63225bd9074ea15a", x"ff7f36944c69612d", x"3fd3ce37ea16d7f9", x"9b1de26248562adf", x"7567d2a4e9e5e52d", x"d6158f1afdee8050", x"5ab7d14faecbe68c", x"1e70bfb24b078732");
            when 27659598 => data <= (x"6911ec5d02401682", x"62c760fa55b1c133", x"49d1b4a22f9ad9a2", x"3de9a5042878fafa", x"c4c0124667e4c59b", x"867c751706a6c016", x"35b682e6020a1062", x"f63d3f7efb0e1b83");
            when 19499048 => data <= (x"5a08fa8ba3aa2fd7", x"228debfd28f1a700", x"4dfd0b389d869781", x"7f431bd3a113e05d", x"18f26d76a881834b", x"d5c0fb45ce50debf", x"2854cd53cc340c8b", x"53da0db51425f1cb");
            when 1686499 => data <= (x"ff2f24b5a026559a", x"d944ec55b92c7e99", x"255e08b291592791", x"e0c03acbab2168f8", x"c4eaa7bb82c5e523", x"2612fe5633eaf500", x"ff1ecbc43056f0ec", x"cea3905461c29398");
            when 21250924 => data <= (x"089671010e025f7f", x"6ec3acf7cfdee539", x"85f87a8220615d0f", x"57ed70661744ba95", x"fdd8c77518a16476", x"d0bbef19e6132ce9", x"56b084b53ddabefd", x"841020e1bd0d9377");
            when 12125823 => data <= (x"bed41698ec65adcf", x"e592a9fe742984de", x"bfb825903ccf31d7", x"e5e499524107414b", x"b6781f5cf3de584a", x"3d988404bda85d9c", x"59975a9bae96f95c", x"2a8de3450f4aaab3");
            when 14665014 => data <= (x"03ff889989aa6fd8", x"8c85cf93d26e00c8", x"c0c3e9dd29c0ecae", x"ad2202d5582f303e", x"f580867766f68ce6", x"47645a8a10c7d5eb", x"6e1abac963c308b4", x"17b74acdde6cd4d5");
            when 17266979 => data <= (x"5b51d589be3bfe79", x"7711100584b64995", x"1387a72dcf5d034c", x"81de0e3dd4076dbd", x"ee1e01883664dba3", x"7b6aaf13a674815b", x"05a2e77488b6cab7", x"e9f9c63148f042ce");
            when 7320381 => data <= (x"e3778a6d6de65a35", x"24f82c5291b3dbd5", x"e7de07914a1e21b9", x"91d194756720e846", x"b2c711d248448428", x"a6a3bc9c7ecda84e", x"d56c53d29215fd89", x"29f0348293f547e5");
            when 5801681 => data <= (x"851665d796d595f1", x"ac8d4557f681a25e", x"6362d3986d567b4c", x"835c275dd74e3dca", x"d784a1073990ab16", x"c899007799c336b2", x"048802c7e065c837", x"32a7d14967b6bd66");
            when 27608398 => data <= (x"09036964a40a3364", x"5fa3170b48054b8c", x"67b5757cdbc02de7", x"872033102307955a", x"3d57eeac202f1417", x"d684c54da885d0f1", x"2cbab47ccb4aac50", x"e6b9e758774d4693");
            when 31216211 => data <= (x"256e19e8e1b1810d", x"7de6552ff08a69a5", x"013fcc56b9fe0c15", x"26b8249e7e3f75fc", x"78c963e9b6b617a3", x"7c8f89f38741e814", x"b81bbe3f91d07f91", x"d952d1ec33431808");
            when 33431870 => data <= (x"65b6d32aa192c5a4", x"09daa1ba2ab2ced8", x"08f2828365fc93cd", x"5fa4a3a26c02e0e3", x"613a38bba31765d9", x"038fc5693a4eb69f", x"0cb7a7161ddafc1d", x"0459635f1f481084");
            when 13248874 => data <= (x"878cfd25e4ccc2cf", x"3e2767df0d3e2ced", x"64905a39402108b5", x"d5506f994b99e10c", x"f06d974c2c8140e9", x"10348d505f2e6858", x"8023a32d65aa03a2", x"8e8c9f910caf0947");
            when 3636783 => data <= (x"72f85feb33ecd600", x"bc271eb140330f5a", x"6ed1e508cb103812", x"9e756b76f24718f7", x"c87428f1bb3c7920", x"b4329ade28af09f4", x"a36a09e684052d79", x"8843dd29709636fb");
            when 28664418 => data <= (x"ec5050e5292e7813", x"5deb305dc403e97e", x"81ac67f81b94d973", x"fd68a891ece28eea", x"babbfbb04df3732b", x"a7aca602887c2368", x"87401ae33c4a6118", x"fae29faca3d8d91d");
            when 8636856 => data <= (x"f1abdfe062f9125b", x"a930dad09cadc8f1", x"3a9164c7cddc3a9a", x"1a3b842b117ea805", x"339353f67c9ac800", x"cdf134a04c55278c", x"6c954c4acfe33757", x"68f7fae48cebef53");
            when 11139417 => data <= (x"0044ea48831893ce", x"739f1144ceeaee46", x"8d8f17d1fc7c25f0", x"b3dfef9709fd6144", x"06674604dc67a18f", x"c6c1acb4a14e878a", x"a63c8478f239b64c", x"169d744aaacf65db");
            when 14399389 => data <= (x"bded2068ef716ae1", x"1cb81ff746e48388", x"5f36f6b2448cb2d8", x"f9d0ebcaeb6f17b8", x"bd499278315126a4", x"da7216d8e49ac6cb", x"122e6a1e85552ffb", x"072e130aa449e831");
            when 31566088 => data <= (x"88f19605f7a2ad77", x"58e0a50338e8bfd5", x"6cdb3d3de05d3e13", x"16a1c764b9b09407", x"16599d79d6c78472", x"84344c1e59eeacee", x"74c23ffd060c56b1", x"12601e6b1cffcbed");
            when 30015757 => data <= (x"fe838ffc43f4dbb9", x"5e0a6aaa90ebfc2c", x"9432dff2464bf9f6", x"6dcbf8cdb9a4a01b", x"0a80225db1acb6e7", x"b66365da8540eb3a", x"d1e8cccd2afdeab0", x"a0a4013c927d0aa9");
            when 30754482 => data <= (x"c9793b684d5986bf", x"944278de634e82f2", x"dabff7d4fed6ec72", x"fd98a6de6daf621d", x"2ed38fe76ac62bdb", x"c7a84972e9d233cc", x"615bbdc793978f2b", x"3f7bfe54cd92b3f1");
            when 16699517 => data <= (x"38c8176f027fc31d", x"fc4634f183a6d6c5", x"579583eaeb096829", x"e1af5298d10515a7", x"52efaa7213766ee3", x"e7e98f08393b2866", x"a1c3f858938690ea", x"ddad89cee70f2c30");
            when 7260927 => data <= (x"15384ab188042f9f", x"d0014eb9a6946666", x"f098cb75a3d378ec", x"dd6c4832da3b06d0", x"9d06f90a8457149e", x"191a037714f8ee76", x"ca8dd0ebdcbe8c1b", x"816be2ece7890b42");
            when 26920475 => data <= (x"f056e1a351a76007", x"b113e3a5ab3b272a", x"e8665b8f1cd2023f", x"a9ca541df26d40a8", x"996777fb4b81de3b", x"2af0fe771397ef7f", x"ea2cca7ac321c51e", x"aff40e168893680f");
            when 12176172 => data <= (x"27a5b1cc218db39c", x"d62cedf36f6dec77", x"ee0a86c3724dc4e1", x"aebe90bf532636c8", x"0ced12222fca397f", x"b4da917c26606aac", x"c545d3e74ca0ed43", x"60f63f5c67f7ce9c");
            when 14169896 => data <= (x"909c6f529084ad6f", x"899a095950691d31", x"09681997a5d9809e", x"685b945d7e926b40", x"db8c58df778428ac", x"07a585b9ca65cff8", x"2ab8fb2fbf6524fa", x"aeb6e6396d72d430");
            when 16260105 => data <= (x"6dca7dda68f10d54", x"9168528ced55afd1", x"5b2a8040764a2c8f", x"a10a4a440cd49899", x"36f4cf883c2964cb", x"05d8e4562926a45d", x"e1deb3d8f4c4c527", x"8edd7fe7223629b8");
            when 28835225 => data <= (x"452422680eb30a99", x"b8f49fe8eb18602d", x"cde6c580b2f32bfe", x"1c883a344303165b", x"c928c74554444daf", x"60e50e3e94006801", x"1d2f7396e1ebc577", x"767d8620cd465028");
            when 23702488 => data <= (x"266571c615e4fad0", x"d14d8d669a32c60b", x"d90983519ee5f41c", x"d6b968aadd9f7c3e", x"02342dcdab4e39a2", x"f8128e0591b3cb05", x"dc28cd62c332668b", x"161b0e3f206257b3");
            when 30374645 => data <= (x"0830358e5b4a7936", x"febe841a455b4540", x"17a3b057853f2aba", x"3aa871511d0e7df2", x"7cbe239cd2f96629", x"1a74eaf838a5d5b8", x"7843be57f9d2be21", x"6e47027f016ddafd");
            when 30803993 => data <= (x"d39b963785e10ce0", x"e60ced91d0c4521f", x"047bd8ea4c69e007", x"0a658e315243d5a0", x"7e4d36b011744cac", x"c0a4b77a3889142a", x"a1066ebf99ef7254", x"3342670f1936c7a4");
            when 24274657 => data <= (x"c0772bb5d331da87", x"df4df973201c84db", x"4fdc0ec6ffd47844", x"7f407f0eacbb49d6", x"5e5699a247865269", x"2d4972e72e725f76", x"4bcfd58d39a838c0", x"be1349ec5ad43045");
            when 32946695 => data <= (x"48df5a6bcfa48f40", x"e4441003c62886a9", x"5dcacf3d587d70a3", x"6a5b46b1d11d9fc3", x"df1f4e01e1eb0d0b", x"110df5b38afa2ace", x"258f8a8f2112753c", x"17a2c108c68787a0");
            when 20483703 => data <= (x"e3c4e46b7d71a418", x"3de88984b149d94f", x"104cf31c9a2523b1", x"bdd44aa02c57f7aa", x"9ceaf001d1cacdd8", x"681ad3860cd3ed65", x"79ecf15426e77da7", x"e3bbde6af83ba3a5");
            when 28798150 => data <= (x"1ca3764f7628b424", x"3c333d39b09d8460", x"27fb0f8be61dceac", x"0b918e0cd31d2521", x"51636d75255ca815", x"de793d8ebb326f87", x"fb5557d6c0f57210", x"8481188b2970a38e");
            when 7837414 => data <= (x"0d7f612b55a89a87", x"0292941af56de897", x"4eaa45f5cabd1c5a", x"3a4834b8b52db568", x"6256c032100453f3", x"40c756591bce570a", x"59ee454ab2997f4e", x"44bff5759dfa58d5");
            when 7081729 => data <= (x"2a48e2d25d333326", x"d920662a4907e513", x"ef20229f0ba2ac10", x"ae2bd92ef2025852", x"bf9cdfcdb2f78fca", x"9ba7f2011b9eb16d", x"a7ae676800ae691d", x"1dc1acaad5a05bc6");
            when 22351380 => data <= (x"865134c05947267e", x"6eaa77ceeba6f948", x"cf4a1f5b5408aba4", x"bd2a58724a3ab3c4", x"dd10c0dd13a2bc4e", x"5abd9f5c208bb837", x"b77dc05e5f092838", x"94b5e846d7975757");
            when 12491562 => data <= (x"a06527132f04ba04", x"5bc58f56a9fa556a", x"d656162d59ba4523", x"d4e3e6ad236cb6da", x"9f661fed8caf2403", x"df68a800a8a7ccdd", x"f07c7a1297889648", x"840a2284b7081460");
            when 19478212 => data <= (x"7b9301a960035a75", x"615b8135a7482428", x"3b5b599fa86e443e", x"d152066d01123ebf", x"c03f22a0d15282e4", x"40963fa27244849c", x"489fdbc78eb3962e", x"7db275e69c1fee05");
            when 15840372 => data <= (x"3a26bd351a2699e5", x"afcea8b6d3e3c8a6", x"8a96b65155d25280", x"c910003b08f233d5", x"8e23ce9642bd9970", x"009e3d13f471bd39", x"852b380cad764370", x"518f082f8bcd725c");
            when 11637296 => data <= (x"2176ccfcefb19780", x"e139f60fcbe969fb", x"9527d1d8bee448e6", x"681ffc81084582b0", x"011c90d50228b127", x"246b61304b311613", x"9f028c7c3f9e7896", x"4f865bb4f28396e4");
            when 17005177 => data <= (x"cdfaa549dfd2589c", x"b83e6b41f13a27ec", x"25c946f2ae6dbee1", x"49dac18a69dc8af3", x"094dffbf5bc91f34", x"dda93af1d00f879d", x"a2dd6511a4e9f785", x"5cd73ffc6b6a969a");
            when 22155419 => data <= (x"928fc6f6a7a616fe", x"d4a4a18763f0adcf", x"4b3d7b32ceb990b3", x"4737b58ab9b6d91e", x"4d9a53ca957a0fe3", x"ab4a6c9bc003f09a", x"9078109384c19bc8", x"3cfb1413a4f242d1");
            when 15925852 => data <= (x"0593f92c37272c89", x"60208105d15632d5", x"e4759cf804d38e19", x"95cae38f80cbff7d", x"258a17ffa6a80a55", x"278f143f26a9a514", x"ddd77159dc9aa2a4", x"22abd5539d2dcd19");
            when 12636301 => data <= (x"f8b3d7e7b01c3b97", x"361376c472b2ec9e", x"b22c2b94f5c23f2a", x"d323c2bae719264c", x"9d26097e18bf5f40", x"b76c47070cd74c67", x"1dc47fd4b4473a9c", x"6a980a155b082abb");
            when 22519871 => data <= (x"4199887485f4d790", x"22f593d7bd995878", x"36d772236d624f0b", x"df9e84fc15824025", x"212aae8a15e6bfc7", x"275cd5dc77f1a878", x"3ae97f001f4f6f80", x"645a598addb1a670");
            when 30729285 => data <= (x"6698df5bab9e7a1a", x"9cacef600507b015", x"db9ed1cb7b4356a7", x"676e5f7780a44538", x"aa90a9b8feaa5bf7", x"762b05ab65952283", x"62214b99f8ce6fc6", x"99ae672c77525f51");
            when 11769399 => data <= (x"c7cc69bbff64828c", x"bc77b5fd7e5afd2a", x"f3e1c50488036874", x"d3d5bcca49b62f7b", x"f1c9e65ee85ab8b9", x"ceee66f2afc1a1bd", x"9979df487d3bc815", x"12cf5d81a47da850");
            when 4794762 => data <= (x"668ddd4ebbb9894c", x"58a3d881bb2c6289", x"60776d192e400aa7", x"fd0b375f672e49ff", x"d803fb4133de5e28", x"6f99063f4f672895", x"2120fcd442ab7ccc", x"604f1a3b6e254ae8");
            when 15758711 => data <= (x"c10bfe2a39811494", x"43e8978cf9f2a33e", x"43038277d8984887", x"63343760de949f84", x"66f608eec5cc97fe", x"d56ad08129857d95", x"df26050ba53439bc", x"82749ddbe962f63c");
            when 7763802 => data <= (x"931a87b68f00e9bb", x"f0c93a4d7ca5f4d3", x"7989a4f951d30959", x"00fc4e728bb5c4b9", x"4ced527795c5b165", x"50d56792dc524985", x"44ee39b9a659e90b", x"0ce6916fedfbfb10");
            when 17986879 => data <= (x"ffa6cbe8f29051c7", x"c87ce9e02b7fa4c5", x"575a2078d5749551", x"9d397c15018fab69", x"1edf17de838fa2dc", x"9e73d1eeecb0f3ae", x"5faf45c58bfc62f6", x"41efeca5259964fe");
            when 15911217 => data <= (x"bd7d19dda6247704", x"9730cd504ef956aa", x"3f1951b273494c78", x"042565bff7f65f3d", x"4a6bfb9dd8eef4d2", x"ef62045612f414a2", x"15323b22a762502d", x"248e6fe98b52d63c");
            when 4100815 => data <= (x"3e9f7bf75b21d097", x"6f6a213e4e376705", x"e379346cac9f2803", x"ad2441e80059a8e1", x"ddc7656f99ac1c09", x"005850a39d70338d", x"bed07e8d9e95d147", x"7cf9446e2e0d2426");
            when 30332931 => data <= (x"31ba1ff199832eae", x"f6e4ef4153ec0149", x"90d64857d3e18038", x"eb18d499162f7b6a", x"bd4fba20513f44c8", x"5a0cce042e905786", x"5196c334eb5c1be7", x"9956671c997478ae");
            when 26512005 => data <= (x"a9d5d6d306cb44af", x"f068120d082a3dea", x"d85b069df9349d54", x"9b8e6ef052ad4c4c", x"0de067da739c2554", x"5af854321ebd017b", x"6aac2e9ab8d49ef7", x"7ef6e39d559a4180");
            when 12006542 => data <= (x"0d6f0c90c453cb8d", x"e8d9abcabab66a8c", x"1e22ba7ae1612771", x"44fb4c1a4c153168", x"abfd4d1c257178d2", x"52a129f2b6d7e16f", x"d1b243cd8f2121d3", x"80cf59371445526d");
            when 22160636 => data <= (x"deea98c431d89fb3", x"9cb6f56fee269b33", x"0f8281406bb8bee8", x"0e2af037c36363af", x"e92b9ce9f76dd0f2", x"6fe29d9d74cb1fe2", x"400ee911d54d6434", x"a52d25a799b87baf");
            when 31903280 => data <= (x"31b0bc126b0afaee", x"5ab7cc86b013cacd", x"4612890a12a6f6b1", x"611a16e25a197df1", x"6f4dda8b6cdd4b77", x"77d8c5bb04d4ecb3", x"837e08f2e635908c", x"0b4166f3e51c519b");
            when 8526514 => data <= (x"5a187e6654e2fe3a", x"ee85f359bdc8740c", x"7fee1f0963b8465d", x"2742df9b0a2f2b9f", x"8450176a99a14242", x"f18f9fa2f5aa753f", x"3d69f49c56e0eab9", x"a27fa4ee55bc1c34");
            when 8882975 => data <= (x"d370860babeb7166", x"e05141785b6e1086", x"51455cb37cca1bfe", x"3ffe7ea21a285e3d", x"4cb2f7e15ccbb114", x"49c342802016c5de", x"4603f6e8569adcd1", x"26ddf5a5fe990aef");
            when 1604963 => data <= (x"b2212d9c79b4d5d9", x"3f95274d0f45dca8", x"c5a574a969f605e2", x"b6db2fec976d3ce4", x"4051f18b833b0369", x"c3de7b7ccac947c9", x"afbf1ba5c5f2a66d", x"c056cd3b158cdb5a");
            when 14985334 => data <= (x"434213bbad23c4df", x"b1143266b5406e01", x"6bec2d97405f93f3", x"d81e1d1e6ceb787a", x"31ee769d5d6ae887", x"531481619c167d9a", x"50dd11683e5b5120", x"23afddb1f1fa80f3");
            when 28109828 => data <= (x"5459707a90d70991", x"dcb1dbfbe4e1ed56", x"4635059035b59e09", x"e3ce68c5c4902bc4", x"bf54041ebd02f577", x"68aa53d36cd2e240", x"3822e430335c31b7", x"e24f4fc6435304c6");
            when 299054 => data <= (x"94d4f17aaca0a14f", x"eaa4744945aca8c8", x"d4501a26106c9848", x"49f7555b078680df", x"39fc51a8a689c799", x"aabc9fd9ac035041", x"f8a24fe83b4aa716", x"e9a97ce04753e892");
            when 734642 => data <= (x"0996e0d068315ac3", x"c77a8b2a91e479b8", x"59e734b12c3441ff", x"02609e2dd1a3bced", x"533312152a6cf466", x"9831fc9d7ca9c74c", x"48db19db1c7a592d", x"f83a478fbb6f0678");
            when 3746222 => data <= (x"7cd5c6c7bc329993", x"3f2ac0b6d0564e55", x"cb7ad7d85c110f71", x"7e0cb66dad979987", x"897440003749583c", x"97f5f8bc91e81ffd", x"0dc2934e6cdc9ed0", x"5757a461e2d11d96");
            when 4509265 => data <= (x"b20ac670d1c4a61f", x"4fd04871e66eea8d", x"a6b4a9aec2a0be2f", x"3a5bf6f1a59d9026", x"f9e162a0453e5462", x"a7e6e1ffc772f888", x"fc40f8a72dc246a6", x"93f0e7e4d519ad64");
            when 12340171 => data <= (x"58e38067c45256e2", x"e363c58de96d8e5a", x"74bb5257f5789df6", x"f7d1e4e61dfa19df", x"3e1509ffe37e6a4b", x"da938e1f18fa79a5", x"62a08ae8c2da7f2b", x"764077dc50547700");
            when 12764992 => data <= (x"fa6a6ed682e8120f", x"6a53293e285b823d", x"17a1f1d495041aee", x"dac2297c305bcd78", x"9c9e42560b98f296", x"f81833e0ef8ef636", x"6a0ff4119e777c78", x"4230d0ea6f297b35");
            when 31790422 => data <= (x"c9808b94150cd3ba", x"a343e775cba3bd92", x"007fab9c78736322", x"af94f3b879ff6988", x"1f04b19d11f6c2af", x"066d676d7920be5e", x"9dc477303d518f82", x"a1e128cfda7aa3a5");
            when 26491072 => data <= (x"39054ec2b8c6deba", x"5847fe45cfe3054b", x"00731c0b9d3df11a", x"0f3c04d675d2cc5d", x"7c4513ebee268f12", x"89379206897b0c2c", x"eb10f78db83c56a1", x"a6f0e907eb21b0df");
            when 2528905 => data <= (x"fb7680b6170b7f07", x"59800ee9fd4e9687", x"824ccb7ebb0763c9", x"540370b2f925148b", x"7836480fc2dd0d9c", x"cf51fb455e202454", x"d0466c75f4970ff9", x"eea3a3447990d8af");
            when 7295782 => data <= (x"ee7892f11273c8ba", x"0f3b236d983c0e4a", x"0efca88a41615df0", x"db1b7e2dd83c9177", x"eaa2da936a4af643", x"ad89ee7ee7b04de8", x"5744ee4e23634aae", x"e58fdbce189e1435");
            when 23568810 => data <= (x"12fd7ce078dd0eaf", x"60d1adb62dd442ed", x"bbd12604ef0e2f89", x"e79472d113d60853", x"d6cd9b89ef9a3ddd", x"b1982eb5bd33ae63", x"08c396faa1259ced", x"514c6c69cf215802");
            when 14463737 => data <= (x"50c34984214b0435", x"98f0042b12828db7", x"741d7ce21ca6c4ea", x"60f40ba03ae4640c", x"a6ce294758910ef5", x"4dc029544c917a5d", x"74a2e83450bbd74b", x"6d9fa1f4eb23efc7");
            when 24724436 => data <= (x"b0513cef8c27133a", x"220b27fec702d5b3", x"91fb3525c3eeff71", x"4525aa3ce43b7139", x"d98092a5ae8563a5", x"6d614d2810ff135d", x"212aba5515bd0524", x"eb077ffbb8f1b946");
            when 18117901 => data <= (x"cc6c44049ac14585", x"8f8e003d4bca5c70", x"2e3ab1048a00c895", x"e03ed4ef67dcaf5b", x"bb9d464952ce0096", x"aa6c8c265b5b25f9", x"9bbce2337b46b5fc", x"d06328608355bf4b");
            when 6675644 => data <= (x"839291c2280ffedb", x"1d5846de9c6fad1c", x"878d9ac07852d8fb", x"55995d1d7aeca7dd", x"04fe55365f1882da", x"e0c016e2156ec9cc", x"c416643e0c228c06", x"68325fd7d53d1d3b");
            when 6654438 => data <= (x"1f1dba00794e2971", x"3596141e28d259fb", x"dc02c861982d3979", x"4b101e23536d8840", x"a83ef5d8b2ddd01e", x"6945e96e841935f9", x"8394ddb283989367", x"5935787d5f8b6568");
            when 10975483 => data <= (x"1a2fe42112bf494b", x"3e93d296fe0f4d92", x"0246a311b040efb3", x"bae4b93a15af54fa", x"e63ea57af9fac38d", x"9307c6573d68900f", x"0cc8983616a8f464", x"a849b18bbb57fcd7");
            when 16907878 => data <= (x"bf47ad3953cb4f60", x"6bdc6b088610705d", x"e555d978bdadb680", x"6065cea916293c82", x"a76cb08c70893484", x"bbd93282570f8cc8", x"b8cb18a0592f85cc", x"57f2768466518c0d");
            when 32329485 => data <= (x"77198899edb54063", x"a6af43592e65403f", x"602ddcd891450749", x"250e1eedaacd8719", x"5c07b4e52da4c1cc", x"1686363a8c68dea9", x"45f56cbe566f3782", x"15f2c7b413830370");
            when 14091605 => data <= (x"e059fda45dda2ccc", x"57ab8747d4022286", x"69bf58c40190c99d", x"dac08fa9e295d5ca", x"508bf908f1ce2d09", x"9a625e34f771bf18", x"9b970342151b34ec", x"c11b11a3e9173d48");
            when 17685951 => data <= (x"37b87a051de5110e", x"30a5fa2fbbb54043", x"c63b98afc3d30ddb", x"fb0a2b75ebfa70ca", x"625438449c0c485e", x"62302579159536f8", x"d49e0e3ba961c23e", x"bd61b570bde30cde");
            when 3335136 => data <= (x"5dc06f5a0c467201", x"cc5506c7cf87e857", x"48ad3941afa89c14", x"e5c59540e8e97a82", x"1c1332dcf56352d2", x"e47b7cdcc4989960", x"a5961d31824d8ef5", x"233e3aef2f3a697d");
            when 11495583 => data <= (x"a0f893b40e17bfe9", x"c2fbaa5d21781698", x"c176c1ef6a5e7abd", x"acac9c4f646a92c7", x"3ecf48ae4f057e9a", x"980a27290b9259e8", x"e5849eba443095cf", x"b5932499fadc6f08");
            when 21487095 => data <= (x"7469786e243abbfc", x"ccdb9c9dcc930315", x"9bc7c0018a912d5e", x"c07b56120cbe44ea", x"0836c63b3cbd4934", x"c0deeb8891e5cab1", x"87764238adf8ce1e", x"80e7b972ec19e74f");
            when 3726330 => data <= (x"fa4dbe1571730e49", x"8aa7198e7d50dfd2", x"83d9f40010656599", x"a5b5a2166f7d85e6", x"8a05c188913eeb27", x"4958e36ffd30caea", x"68b25f5c441bf6ed", x"933b930d279fd6a6");
            when 17408540 => data <= (x"40ed11abbf51c0b0", x"b03b59e37be51009", x"5a64050266d4eefa", x"deb84ceb3f4b3b87", x"2d43a4e45d0ec36a", x"b2574015eb2adc7d", x"0a4509cb329013dc", x"3a8ce7ecbf159599");
            when 20544018 => data <= (x"b1845b11cced3b6c", x"fcad00fa497ba965", x"88c7e8cf0f1c8392", x"eec4c6137c9628ce", x"fdb86af958549698", x"3c24570757697078", x"3a96304991e0836d", x"e9324ed0d7c5a6f6");
            when 2074276 => data <= (x"7f6a3b607e1d7867", x"12b1152272d70018", x"6e7dee881c3be567", x"6620f31044b1666c", x"40dd93554f7c6793", x"032f827d9a0b9414", x"0bf2d77d5d9e00f0", x"091683457634a21a");
            when 12908187 => data <= (x"75d85565d98876ec", x"dab1e66c52ece7de", x"d873f442d2877704", x"2745810ed7b90432", x"ca7f575cfbca84f6", x"fec2c5ba7484cd73", x"a5262cd19207425e", x"327d0aaf08a65526");
            when 29547584 => data <= (x"c6020a1193c9d064", x"07ae6096cf90d7c8", x"caa71f2de5ffe842", x"569def37c7bdba85", x"54e77cdc5a6cee34", x"7df5dbd8c15fbd5f", x"eaf4cc0a03bda895", x"46716862e5a3181b");
            when 26024841 => data <= (x"61d7cf3b54b71397", x"ca87a26c61cd1c90", x"822467d24813d461", x"e6a29a3c7a378588", x"a465ee49ee3eee0c", x"1726c4e0835af74a", x"9142874749dc406c", x"7a8a6f68b1e0d1fe");
            when 13645373 => data <= (x"7ba647adf8280226", x"09839fa92384740e", x"c46095e3415bbcc6", x"3e5cf3e0eabff5f3", x"4432266596ca4d61", x"c44586a1c8047883", x"01185dc5167b0135", x"84501b8b7900b5fb");
            when 5706344 => data <= (x"6725eb43ebb959f3", x"917c80d64de1f3c3", x"361f4dbc77d5d9d4", x"1eef153e8a85adb1", x"215a9ed4353a5018", x"cb545095d75bdb1a", x"d36283cc67cf935d", x"a5f5f364afd15bd7");
            when 27177707 => data <= (x"0bbb54898ffb9757", x"778f8067e5e4836b", x"2e81b4b6baef47a4", x"e1f9854867f2a4b9", x"e3d665f3229c4f9e", x"b27ecd90bc5002af", x"05dfb95ef08e7ef5", x"cf73516ed755e03c");
            when 10839798 => data <= (x"703b11d2fd853284", x"29106a7a37fa8dd9", x"80787d423dfb01bf", x"876e73a7847c5a4e", x"92615e5adf6a645a", x"cc82acdf58d85f8a", x"b3a90d76e35bd05b", x"429e7112a85dc707");
            when 5533999 => data <= (x"89cd2698d7b9f8b8", x"3cdf9dcfdc1ff3ba", x"153cc30a82f4fb96", x"3267dbc3c4ce9fbe", x"8a34adb244de4961", x"4a574de41ab8922c", x"047cdab109cf6210", x"c41e55509c157dfb");
            when 20757807 => data <= (x"d3bf7c399406ae16", x"337e9dd907be90dc", x"61e58bd105761a89", x"9d8cc6e6533cac5f", x"d01bb88c91f238f2", x"a14849381b04c59f", x"debb97935acab938", x"437ff884b7d5b2a7");
            when 29668725 => data <= (x"514b9b82bfb45ca2", x"7ae578ba04999839", x"784210345dbd1eef", x"5e5910d2ac14778b", x"ec3e42e8404ec356", x"9aca80c59e9cd798", x"9f3e794c7188bd77", x"99173635ab04d4aa");
            when 29458944 => data <= (x"494657512a11305e", x"3f11240cb0a1dafe", x"bde8a8a406c73a41", x"65bf106537b8902d", x"ca541dd547f6c70e", x"87ae9d36c51fe013", x"007ca7ec9d5dec4e", x"34bd52804c872cb9");
            when 25229827 => data <= (x"cbf3cb6810c32a26", x"a605054b5ed0bb86", x"9a9a5f76c16da083", x"0883a2d5c5b93730", x"583485ac42a25a73", x"6f7c8b91ef511e00", x"b3f37b53b0fd3944", x"0c0623a680bdd6e8");
            when 11816461 => data <= (x"60be943959143e82", x"b47905a397e3c907", x"463158666f504ab2", x"6c526b47fbd22e7d", x"548ff666085cfc0f", x"6adfa35468c78b6c", x"07bf3847a530915f", x"7033430bad7ca97c");
            when 29723730 => data <= (x"0bd99f497204d52d", x"dc69ff5f2fea5da0", x"42817d08563d4500", x"8197ee79ba23dcf2", x"51b4bcbbd102090a", x"a7b116b99d038609", x"54e3d4ccf7ccc661", x"69fb2d7723ec5633");
            when 7342494 => data <= (x"e25625ea43045b27", x"a50278a4e4d25939", x"b928383351208b24", x"a20d72e30eddea34", x"a5afab0c9b73e8d9", x"9c7e6129853fb6ee", x"11d384408d6a3c63", x"434fe7714329cbe4");
            when 12227216 => data <= (x"0eef24cf2dc03008", x"da59f4aeda3f5793", x"ec166376116d1590", x"8ea49933f8f74556", x"813ba1980006e258", x"5d9ef45fe1293d41", x"b29e74042078cea7", x"eb78180d97eb822e");
            when 28571095 => data <= (x"be09aa165348cafc", x"5da9952eb57a6519", x"c7ed38b9ec4ae420", x"a9d880663c28d691", x"19b2eb85ef2ce031", x"c9676275504d19ad", x"8c8d9841e209ba71", x"717e68981012651c");
            when 29123706 => data <= (x"eac3fc32f61d290d", x"2f05fab1ceb5ac24", x"badaa979b5b6b6ee", x"265ebb57aa174970", x"82c327cf01e60242", x"a6475528a285f864", x"5c1c4c17342ec324", x"f28f9f9da8e7eb69");
            when 22231815 => data <= (x"cdcd004d6621d826", x"ac73df90e0bb7e2a", x"58ba636be119aea8", x"64075adb49239e48", x"76a3f22f79e9578c", x"2bedb20c7d7c6eea", x"af155fa6465fc997", x"6a3a2fc9d9b9fb42");
            when 17292162 => data <= (x"9c4ec63a4083261b", x"d2238e5a26227492", x"b3367ac605c35223", x"5ef2d033988ebd46", x"a003b65b5d45f280", x"146e4fd1b0845948", x"dddc48026992348c", x"29cc923e496e38fb");
            when 1751307 => data <= (x"4dc9bf27f5b6c01e", x"144f687f8fa0f8ab", x"fa3296249d4bb7b7", x"9d88db572d63333b", x"9011347e07c3a5af", x"e19c9419c63faf58", x"85b935c50a147597", x"5acf1a0a5e77add2");
            when 12529397 => data <= (x"07a02b4bf8e25cbe", x"5940c5ce26017534", x"68693b95d9ec3a4b", x"a07aed2ddc5aca2f", x"dab1f808c1831150", x"f1c4544a2b2c0ffd", x"68361cff143d102f", x"5b9dcf0b310cdea9");
            when 22425339 => data <= (x"f8864d2f1a730a6f", x"fbb8758066509bbf", x"0f6724461453f73d", x"cef0dc6fcfbf8353", x"bd5b7b7fdcf35d91", x"033b03c88fb0b0b1", x"07cee395e2716252", x"159a95d56dcbd769");
            when 6996865 => data <= (x"b5708f4040586559", x"985022c6ec9f6067", x"bebb26f71ddb4cc1", x"d1cf77176378ebe4", x"c4cf0cc8bd11d6ca", x"6009b205dd6a9a64", x"6f48959179d9e87c", x"b7bf84734b52b683");
            when 4128267 => data <= (x"ddcede78876b8964", x"a2cbd2307ef41272", x"d890a8073ff4baee", x"40d767e722ebb561", x"6d3c8929abe96a50", x"790794a242d84d75", x"bcaf5de1815c5fed", x"f77669eeb9177f22");
            when 6713133 => data <= (x"4f8e71dbca10d8df", x"69e4cffebdca85b0", x"6fcb124666055742", x"0960330a9e703410", x"7cdf94e9705e81dd", x"d1d230d5304d9014", x"c5a935b08fbdb578", x"59c47ba7e77da88b");
            when 1582405 => data <= (x"dd26ccf2114ddc70", x"02f894e9bf373f8c", x"c929e618d768d93b", x"07a368e97b79b0d6", x"46f718525bbe1d38", x"c0c1d296b6bc893f", x"b8e2b7fea2ec8cc9", x"012677a66438eacf");
            when 3406673 => data <= (x"75ea6b5c28eb188b", x"40dcd8b2849e5304", x"4f28d8fe36cf8c03", x"42f600c1b31b4a22", x"8b51a1f632956760", x"5686776d1a947d83", x"655b70766950d53e", x"e5f647ccc0b863fc");
            when 4920508 => data <= (x"3a9950add473908c", x"562590a9401d6ae3", x"47056012f776fe59", x"66bb963f99d7ac7b", x"c20e5abe24d0b7c6", x"e368fb160756b690", x"c26c8ed035af4ce9", x"9b061b29d9049320");
            when 1363275 => data <= (x"2a70ec9b6349d783", x"8363f4c7f4f3be82", x"bda2b45dc75029b6", x"05ebebd119f58bc6", x"dc7791bf05cfdf43", x"eaaba4d15ab823e8", x"aa41b9efc5bc8fac", x"51befcb8fabe07e7");
            when 16217229 => data <= (x"8e5bd2f2a4fe8d1d", x"76cba14a59fa8f0e", x"9fcdf6e905d5b107", x"15835b8b27f5e8bc", x"4a56a47cc7caa6aa", x"2748212b179a9ebe", x"45a5ea4ca66114aa", x"9dba745ef74ce4b9");
            when 29353114 => data <= (x"20d75dd75989f4ce", x"6251608c93933480", x"04c42fb5af52f40c", x"ff0f5bda4909f53a", x"f6bfcc5907747472", x"96768dc59805fc48", x"c8b8f7d8a01ed2aa", x"4720477dbe3b7164");
            when 19158086 => data <= (x"91ebb0a34a4959fb", x"6b3cff8cf9b938ef", x"410a4afdab20c262", x"b86027e25977a8ea", x"4b09ef036f8755c5", x"2d118bc8e5a380b6", x"89adf0aa1b2ef140", x"c5beed668d24c28d");
            when 23060422 => data <= (x"6c29f92d336c9b0d", x"a501a5403d136097", x"86381b6d4fc51bbd", x"08f08c3329113ffe", x"2dc8fd333e721735", x"43e0e17cbd96b6fa", x"1850b6b3f2be0a44", x"958fe573e160958f");
            when 6708434 => data <= (x"dbefa684ce6c5a0a", x"43f0027924b62d34", x"1dd5c02cdf831dc0", x"52e481ba49100770", x"abfe040ed2742d89", x"bd426db8f93c430c", x"94ca50aa7dc00db5", x"9a9cd492880f8d7d");
            when 14201378 => data <= (x"d038775f2f4c146b", x"50d89b910edd491a", x"796f5234ebe82032", x"f0991226169cdaa1", x"91bc7f206423ae3a", x"5407f81413485f55", x"d1da786d778d69a9", x"464c216c62358c3b");
            when 5915458 => data <= (x"dec1168371129af2", x"123297eae1b118ab", x"793c72f625cd4709", x"483fb0e9935efa06", x"a859c29fc217109f", x"e3d0b745100db44b", x"4072a2973051cf06", x"3ae4e492917da18c");
            when 19834334 => data <= (x"92ba186f7cbde3b8", x"5989a7bdea572ff9", x"ae8c6f4e916368ef", x"9438dec2fb3681c9", x"30dac00d99e9d83f", x"ec745b3d8b2d4e7f", x"deea9a609c4315ef", x"c2a90321b5c01587");
            when 7493223 => data <= (x"9c15098e4f4dd4cb", x"b458e44512810aaf", x"bad190a489ec3719", x"e72d8643ef95da68", x"9a6b8eac8b6e6086", x"0b57df262b56b7c6", x"5f15749572bdd6d1", x"3b48dd047a26177d");
            when 16162545 => data <= (x"595349d47ebef838", x"ab01420782c76a70", x"565b6b42434e38fe", x"414b50835abe03e8", x"6b0ff9364e9bb4a5", x"18d8103f388418a4", x"e93a80bf29fabbb8", x"6087b5644e3906b0");
            when 23572428 => data <= (x"25a608b5e22d327d", x"6cb7ff82421ad5e2", x"9f522ce19fcb3a81", x"dfd986f3679cf43b", x"abe358b7846347f5", x"64e5e9c3db13d070", x"9b2d2edf12bd6816", x"96d42f1d73fad17d");
            when 24910366 => data <= (x"b43182eed64c708c", x"1da99e41feb089be", x"95935068ee6bddc2", x"d7d20af4a50871ce", x"1d37a688fe2f7534", x"a0ac97f6a88f9e74", x"73d041f3789987c7", x"af72a64beb458f65");
            when 14905992 => data <= (x"4f2ffd9946e24d45", x"112c7f5e48506b2f", x"fd84c6f7bbff146d", x"236ecbc60676bceb", x"8fd216b4144f265e", x"ee3563844543fd12", x"8e11727f60d8854b", x"a6dcbd244af68eb0");
            when 1606564 => data <= (x"23a0aa0d7e1d396a", x"1aaede40c3086212", x"9629e26670a3bcdb", x"d5399d29b1acd9be", x"0184c95fc5d8a291", x"78d2525143d69cb8", x"dbba77f9a4eaa8ca", x"de0b624bfcd4c107");
            when 17506740 => data <= (x"3e64c7232cbae698", x"9f56003e47288eca", x"c3969a2d8663dc11", x"e0d29f7c583b8a18", x"713a9099377f0f95", x"2f255b4075c360f8", x"e0c67d09339798ac", x"d154a30bd2d4f0aa");
            when 7211057 => data <= (x"811e412c7a7e0788", x"a25d1f70fde4fdc7", x"7ec95c6639bdc46c", x"a644b907498f1272", x"621642b41708a25e", x"b46fed1e39499ab4", x"e4e0b911e07f6591", x"94528825eca8d4c7");
            when 15247434 => data <= (x"e0c43eaa8b60f9fd", x"dfb5ea33300a58af", x"e68ba23d2cd96c5e", x"d35f2fcb0f948dee", x"e62590096dc9ff0b", x"5bca2c75880e04fc", x"ce0e8458035f081d", x"5cfa96cefb4d0618");
            when 9310574 => data <= (x"50907e9f47ccc925", x"8fb6bbf702aa1980", x"61fcab10ea9814c3", x"05e1f5c88ffc8f02", x"ed8515edc3105b49", x"92e50ab50d8a24a5", x"fbe4f4165f6f1171", x"46804e6175e9ecf9");
            when 12213900 => data <= (x"97d21635b85c282d", x"2d09dd6fd9ee65ce", x"e4442b17500e14a7", x"a066309b25d05aba", x"6b9a578ddba61078", x"fdb89be5c6b12030", x"9f91fc1af12b4c1e", x"8d61900f0082eb92");
            when 1401583 => data <= (x"9ff66f78bc1f9f57", x"2eb2c6dc5eb2bb78", x"9a7c85b691b92ddc", x"d634f5e534b332e0", x"ff135653593209e9", x"0638047e1091c7f0", x"4ba782442359a457", x"8a7e2dfebe2ec214");
            when 24535417 => data <= (x"4b8007c822c3f88c", x"559ae7ecb755cc47", x"5fb37f6a6d54107f", x"1236536030d88c98", x"56e425da5a501690", x"8169e864507dcc96", x"781c19ecb021dda0", x"c0ee03f21d1efe83");
            when 11989945 => data <= (x"b5509164cbc2910a", x"0b7fe027aed143c2", x"ee2d45c74bd047c7", x"bff7251799714eaa", x"39d8e6d60e8c1528", x"18c73070c45a5f39", x"4de0cbeaff5c9446", x"c2ac62449d40ae03");
            when 224849 => data <= (x"0972595d4e15847a", x"a81777214a1805ac", x"3e1daed18453789b", x"846a308236192275", x"f67830c64fd0ce5b", x"5e6612406b6af126", x"b56d7f9ae248a5c4", x"b38af09f5e5f939b");
            when 20108576 => data <= (x"2d65e405101dcaa5", x"a0bdbf52722184e3", x"705eb3a7e222003e", x"65a11b85ed5a3dc4", x"1604257bb89ca401", x"33f39e2476654d5e", x"d043d5be80d12baf", x"72bc6879a10edac7");
            when 29292413 => data <= (x"65b289be7419a1ff", x"f3e0288f66de61a6", x"98ec69d8e7a744e8", x"8ec0d167932e18ab", x"f45721dbbb000b79", x"2c590719b14d8144", x"27eb0031ca721fc2", x"184a35b8ab486c32");
            when 4842533 => data <= (x"a2f06a5341392877", x"9b0425588c62b296", x"e31e57f80fe56a7e", x"f5c4b742c56605e9", x"908d13bb10702ed1", x"ede8217929666521", x"6b15e2b3a3d9c6b0", x"7b17dd556a525434");
            when 22156639 => data <= (x"a75fbb5b851ad610", x"8a4d1b0bee1fc4b6", x"fef5b5b195188ee5", x"af643b65a2bd286f", x"1e15d8eb66dd7379", x"0d81af9a2accc2a0", x"386b1bcd8f447499", x"789fd8f6c19edc7d");
            when 23596713 => data <= (x"cd03ffd16e2e2ff5", x"b63bb29409f450c3", x"95ac4371d930881b", x"e1440832403aed79", x"216d19b40b793cdc", x"ddc9e96981e296ea", x"04af4c01799bb4c2", x"fa663e1cf16d6281");
            when 5166059 => data <= (x"d46ff610cb963fb0", x"e859dce30dacd5ab", x"99395220fc0f2a28", x"dacd72405eb159c3", x"66398d36fa5b6f10", x"f13b9e24beb0bfff", x"0fd3e51d8021ad68", x"6962259202e70612");
            when 29949824 => data <= (x"e63a719693d0e57d", x"128ca52136b6fd43", x"bd9c9c39a1342547", x"04e8562340d339af", x"d55f627b40148a2a", x"b87da6142748c775", x"45086b149ba4046d", x"060e51660da40018");
            when 2574983 => data <= (x"dfe920fb6a64203a", x"83e6119c04e19581", x"823ef1bee5930ac3", x"f2a4af8e05b5d375", x"61b13d98791d08a8", x"382186f8b2c7e85c", x"a4ca3c42a2364943", x"683f63bea4d18c58");
            when 21630565 => data <= (x"ce2ef223ac0caf76", x"e7b21ecf4f6bcfb9", x"9e44f38d39ff7ce0", x"29fba4185ec3bdd1", x"5177f2b2c9819ac6", x"0ae6fcc8be57ed14", x"2216aa217a18bafa", x"b9a5555ba94b5cef");
            when 10372875 => data <= (x"360dc0cffe5b21f6", x"513350e456bbe994", x"65cfc582f12e1b32", x"15fad0e7ca297560", x"5d1eccc5a4761a11", x"85cefccc245da7a2", x"9ffb1e4503d6e3de", x"84bba738a829b7c1");
            when 17521915 => data <= (x"66beab4d6b9baf9d", x"3d141519eda140b1", x"47e7aaa65b316eb3", x"8bf6b5a01782bd8e", x"44cd00730125a8c1", x"23e4046a924420bb", x"45f2f4c2f1679ab8", x"90fb76e3833375cd");
            when 23415561 => data <= (x"e90d40673b15cdec", x"531be6a594868ddf", x"2cc883c5e4481d46", x"375e80d61e0fe6e1", x"ca3977a3ada6d1e0", x"3928654ca8f852b9", x"0ab8e3f9b39ceeb8", x"ccc908dd9e4b7b5b");
            when 486926 => data <= (x"f41a1b98dd40cb13", x"5c5a0e0ec40ef73b", x"e6611b01e5dea42b", x"c9e983bf931a944d", x"f5644d04e46d69ad", x"4b1cfeca91ff59c9", x"b1d0600f11ab37c8", x"e96f5ae78ee7ecf6");
            when 3212534 => data <= (x"2fdc033d29a762c8", x"b27d1bb03f397419", x"872e63ea87d132e3", x"0edce1ee1d4e99c5", x"0ed4458d7ed5adf4", x"ad3200f393299b25", x"d47fdc369159d3bb", x"07587dadd1fe1c83");
            when 9035840 => data <= (x"3dcc8b9c2dcf4a24", x"e9df098a98d813b5", x"0fefe8e3c38f1656", x"73c2cba7d666f104", x"0488fdb5e4ea38e7", x"5f17eeb6b911fcc4", x"f729a83d151676ce", x"ea6ab7a9787225f6");
            when 26726946 => data <= (x"9420205ca69d3f9c", x"297206bd6f069a78", x"8fef2a5fb744e7de", x"d1667d0adbd8f70e", x"3e4adbf96efb9147", x"327ec352e3165a8f", x"9f9efbed1d4a99fd", x"5326517da48356aa");
            when 6061618 => data <= (x"f7f421fcae81e64d", x"c7fea6a744f5ab88", x"1150b159c29e50b4", x"e905d65963bf3a35", x"0e53a9572493be11", x"39ee062146b231fc", x"0ac12d91358303bf", x"7e480d5e67d1bc4a");
            when 12932860 => data <= (x"861ae945b004606d", x"dd81a0824631d334", x"00dd0fd4edf74006", x"003d6a83c03f33dd", x"1e3e14a87982294a", x"e37921690ce37881", x"4bdc04285e276452", x"85bcf0e133783155");
            when 20018722 => data <= (x"85400d01483596bf", x"c3d542c014e65e71", x"969a4e8a895575a2", x"cc3a31f3c55bea06", x"29275843cb0ff388", x"d3e59d43248b4725", x"01fd53120b0fd20f", x"2b171bbd7951a21b");
            when 5042521 => data <= (x"6ed5eb501103756b", x"23783f886a1ea3de", x"131f36dfbb06b3d8", x"9b7809106b116e30", x"0efeb3a5fe8134bb", x"217333ab0017e6f7", x"2cabf8daf914cd29", x"e9b72526e05ab062");
            when 32399833 => data <= (x"0d895a2f845b208c", x"5d781675371f1e4e", x"6889a3dd0a6d4cd5", x"7d41dd0482760dc1", x"8df59379d17a12a4", x"a6ebdb58385d5972", x"c46dd77e3a57d876", x"bd66793a27077350");
            when 14890077 => data <= (x"944f3df13b0ec878", x"e24afd47e3f021e8", x"372234f99d8dfcb0", x"358975c245574f77", x"62bbc9c9562524cb", x"77ad24dc3561c77f", x"50ff42dce4a37695", x"c2764706d26fa054");
            when 26400100 => data <= (x"1b8492cb57abddff", x"a2ad6db7e53a03fc", x"aa1b3488f42d9be3", x"ddf71453002ac229", x"afaff53a43b8de6b", x"4ef5e1feb540732a", x"d763beb5b5ac61cb", x"130ba4416a19dfa7");
            when 20817174 => data <= (x"2c996107ff4cccb0", x"2ef7340dd3d2a52b", x"5a842bd33e519aba", x"dfa98af9f34759a7", x"720e8192c60dd3bb", x"20e432777da58cdb", x"550423a5a58a1fa1", x"cfcdf9a821894548");
            when 23066760 => data <= (x"c169d641d80c8cdd", x"c068f4a1a83310d7", x"fa16665e1cb5d4a3", x"248c26987043c4a4", x"bde783c7f1b5e6bd", x"60ca117464178bf8", x"16edd80f0f675896", x"8e65924610f603aa");
            when 8539004 => data <= (x"1723ff82e2d03002", x"5a79bc72b8d5d82d", x"f2382340b0a33ade", x"ba5e378945e91a31", x"180f375ff27ba54d", x"92ae602e45e2fb63", x"05637755c924211a", x"e66739fca1d78323");
            when 7136853 => data <= (x"04b8dc8596d377d0", x"8a4670b6bd5d9a68", x"26837edba7e11fd5", x"910a5204cde0077e", x"f2d0a9d9cced5b14", x"3bec423b96984fa3", x"291d23d5bcb68493", x"5c4b7db7896a243f");
            when 12140673 => data <= (x"9487e79618e46e10", x"98901e34aac3372c", x"56e59653ba27219c", x"4d541a47194a2852", x"64ea28df47d2fe47", x"fcf07d0c073c8d29", x"df0f6f32a2715483", x"a511990bb81c4adf");
            when 18252411 => data <= (x"317d39ce6f659720", x"e05a3168afd661e3", x"d72455132f14bb38", x"9ad523fe34069a2b", x"9c62cbd1015b3774", x"c67bc9aa8c1004ff", x"cee227c5a7f2a2ff", x"6775d0dc61483c28");
            when 26983323 => data <= (x"35784003ac42be6e", x"1ce18c45fd6be357", x"c547c5011b496654", x"6ace99c43a2ebd81", x"c77ca791e27c007f", x"e17c1e6547b5a2cc", x"66cc91ca155b66cb", x"acf8c9e8a925d323");
            when 33511971 => data <= (x"f3d99146240ec81a", x"5c4e3af663f971c5", x"376ecbfab9db3653", x"cd721554188a4644", x"a95ae36a16b8371b", x"3c04592db597c956", x"ce6ed92399abed2b", x"aa55c8a818c7a0d6");
            when 29828151 => data <= (x"55b111a2a5179b75", x"555189f2a8daedce", x"7eb942487f115cde", x"73d8bad33c723ed9", x"6cb8f306a03b8d1c", x"dc67437683b323fe", x"ea01ce8d574f7a82", x"8dfcd8c8fb47d208");
            when 18436164 => data <= (x"352fb2795bc5cac3", x"b9e0581c130fa077", x"cfccd7b5932aa45f", x"25bd13d2ce1ad77d", x"c0fbbb13a7ee246c", x"a77ff9f3fc0c37e9", x"30380a798880cef5", x"4aa681ee98a3273b");
            when 28834879 => data <= (x"b07fec3b17ee971f", x"3f0fd2540544f1ae", x"ba74c572e31dcf92", x"aa571ac6912c82d0", x"a4563eadd96d1967", x"f7f41f75d3c47a05", x"ea77550853dc44ae", x"cdb22f526a8fe424");
            when 9048760 => data <= (x"1fd63bfde8e48a9a", x"606d471fad8b0361", x"c92b902d8ab4f968", x"9b19d21507ffaa07", x"339f777ef5cd4467", x"b862b0468bd133c6", x"663f5c712eab45d0", x"3e935fd426176ade");
            when 8241314 => data <= (x"74822032dbb5c536", x"60b6a7fd5b447bfe", x"4c0ed0fe25c8174d", x"a4ad84a44030b8af", x"2ba094914e0f167c", x"e0ef33743faa7471", x"3561ae3dbf3375c0", x"c19aeb913f7bbff8");
            when 9059648 => data <= (x"cbd11cbcdd2092d4", x"84535cfb047aff45", x"d312a07e6a4da766", x"9836c4d2d7a02ef7", x"07a3c0305bfa085b", x"5c96b9b4e0bfa118", x"8ba35921fc274659", x"de2853575d32e47f");
            when 32422983 => data <= (x"8cca007c5081384e", x"91230d59ec97d9fb", x"0147cdec62740879", x"fbdda7ce2cb5ee19", x"a6cc8b0761ce463f", x"78f085d6c1405382", x"5a009fc9e191806e", x"d0f2e482da9e4ca7");
            when 20840630 => data <= (x"e6d2e33940ae1439", x"e45139daf27e4bf5", x"a53068dda01b15a3", x"6633d586574f2f06", x"a6cef6b5f50a1d18", x"d1e1128342c33e4d", x"bc215e806f082d60", x"e660c7030ca217df");
            when 14748371 => data <= (x"a7f34e7b465b51d6", x"7a4cf59bcd0e855a", x"ba981152cd2565bf", x"3c8109c7a8a6ca9f", x"b308a6d5dbfbcdaa", x"1ffdfab70c83fb5e", x"d3d632db1f0084f4", x"c0cad534b79c33a0");
            when 24144516 => data <= (x"42aaaf201c037f02", x"ede7aff254e62525", x"157b55938ebf3d5f", x"3e01148ee20c9d05", x"a5faab2efd933f23", x"0a2a7e347c7564be", x"bbf6701f6f3d9b71", x"55f75846a997ea57");
            when 9627044 => data <= (x"65875c9cb43c9f23", x"0ff473946d124e19", x"4ea4f043c86f9fc2", x"600e5b853d2f0e79", x"77b57e4ef23aa72e", x"bdefc071db54c386", x"c046473cf29acc73", x"47a785d6487bc4af");
            when 9173693 => data <= (x"1f1f5f30ec5f0d93", x"38d6f484c8ae1423", x"3868731da4e8011b", x"10744fce92b8cc0f", x"bc5e826238a0cfe6", x"4d7d87acc232eaba", x"3f9af9e58e587aa1", x"7f0390611476efa2");
            when 28037436 => data <= (x"24c710cea3d0ea29", x"c9ff04ad9cb1e699", x"ff1290f67cf2e209", x"0f8b190a86a412b9", x"5dcf51b85d545c7d", x"5e1652ba03cc26b1", x"89db57045ac7f2b7", x"395be83b3bc736ea");
            when 27308132 => data <= (x"15d693f5855a3158", x"ddc3d647974a18da", x"a4f3392fc52240aa", x"0bfb91fb4dee5a5f", x"55ba13e089a365a4", x"97ee921d886bb6bd", x"ff49966a8064c88f", x"918aae7c9c24828c");
            when 9215314 => data <= (x"77674e8f60c5d9bf", x"d0319fab5765e5f3", x"acdc2404b3b06564", x"b1d6ca944b2a01e8", x"583ff6cd8ada7fc0", x"83235a8330d56b44", x"51826ab6353b1193", x"99bc629370376163");
            when 9981966 => data <= (x"ca20b13a760e4e2c", x"d7c428ef2163226c", x"4892862d53bd27d6", x"ccdfd8c8764ecb00", x"5c1d65af344f3437", x"31daa7778908f47b", x"2224e4398be350ae", x"38636967c094f071");
            when 25382478 => data <= (x"51e44e7b30c04d80", x"04bb638b666ed977", x"2d785f628685ce28", x"4a30a4bf5d935918", x"a5317370dc0f637e", x"092ad12573ee0ad2", x"ccb8ade087dd9bc8", x"420a793d2102dd81");
            when 14911032 => data <= (x"06ee6f3c3500a800", x"d568b01be9e5e0f7", x"a4a433e56e238033", x"f25daef1cac915a2", x"f778f2f03cdab454", x"86e0acd36bb9b8b0", x"f81a99fb59e6e875", x"28add2efcefe132a");
            when 19178067 => data <= (x"2d508ecb9fb6ff8f", x"7684b0fd645fb4ba", x"fdd5986abcd25a99", x"f3676a9a4eda0ee9", x"0bfde7819eac2eb2", x"752bb139dac0dc78", x"c1331b293d7baf8a", x"cf18c0e39bab7525");
            when 14202757 => data <= (x"81a630975f39ab1a", x"1888d589319626e2", x"12c6114f059deb59", x"b51e7f7e24deb737", x"377fdf818f58f635", x"79b3f34751cb6c7e", x"5ae485efdc9c07c3", x"c9484d0342a7d321");
            when 14720703 => data <= (x"0104226cd760a1f0", x"16c0a527f0531663", x"ba445118bc40cf7d", x"16d1ce5ea70b280c", x"a11e49d3dbf0ac25", x"d969853d003de85e", x"42708ff8a44f6150", x"1c8ad514969a0064");
            when 27310758 => data <= (x"1c7507f8dfa01ff2", x"7c68f420e99ff6a3", x"165aced535547d85", x"5e05cd360e34bd5e", x"3ff3043ec64c2744", x"bcc927f63a1b2b49", x"1f7014c9a80bc216", x"8e3e9a74f9a1738d");
            when 15661145 => data <= (x"d6a67309e0e8b7c0", x"284db697facc4daf", x"e5ff1e1ad491d151", x"a7e79db291ed0554", x"e5f4aebc67d3c347", x"0c764cac24b0629d", x"48e28c3f612ad017", x"95f4dca345f8cf54");
            when 15015504 => data <= (x"9d73ea4d01bc9b6b", x"86b7aa41986b1995", x"f80cd9981b03e814", x"2e73e93a4d26986c", x"813c89311174b1d2", x"d03ecedd5d45c21e", x"7d558e566d7378e3", x"b87d674d3448e536");
            when 20111935 => data <= (x"72bbe9d0bd0876fa", x"f7726477587e6668", x"124debfd40ea8dec", x"27745bade921b440", x"87e91c7343524b36", x"a8ec34de27a7fd04", x"d0afbce08ae1dfde", x"b29fd5429f34ec9d");
            when 4327320 => data <= (x"d4a678d2b4ce05fe", x"78717dd4f7bdf28f", x"7b2c1ef0dd1dd53b", x"9ec9f479ad053629", x"3dc549014a59d8e0", x"dd57b4fac09a6ce3", x"80f119575a629909", x"fe6b853545ea76b9");
            when 18796672 => data <= (x"728293f3fbe242ea", x"0b2508069da1d2bf", x"ab80e28aafac8e93", x"42403679d3290d7c", x"6f22c78b0c1219c6", x"264fdedfe0c13565", x"45b08940731d4d95", x"a1d02d5652c2254a");
            when 32034640 => data <= (x"ff4d46f6443c274c", x"6c0f191ddef66ea0", x"493c58973161223e", x"2d7b387bb5ff7f33", x"e1783ccc9f8ff48e", x"1a5144f84b58b4b2", x"08ea0e379a3c91cd", x"d0add8828c20f050");
            when 8154247 => data <= (x"59bc33c2597c3fc5", x"364fae951a34fb75", x"9a9b7687a6f7e4b4", x"6d0210a57e0868e1", x"014d02ba80de6e5c", x"5ce0d2e606ce001e", x"f813e97f020215ca", x"ae586a2e5ea59eba");
            when 26556269 => data <= (x"e59f6a359b35ae2f", x"61f717099d05c652", x"a49e16604be89505", x"ebfed473c67bbe79", x"4a8d76f06612b50c", x"675acad4cf371805", x"28c7a8afaff3f642", x"22f6c3fde66b9ee1");
            when 33247689 => data <= (x"0aa1916c3981e979", x"dc804067d15d2d5c", x"d2783c7296e6bbc0", x"2e8020dc2d486ff8", x"dee752eb360ba357", x"70dad4001c866cf9", x"d1f0661a4045efba", x"1870011921deff6d");
            when 1484804 => data <= (x"564f40c3d72b0991", x"48385dc383df153e", x"b06ad9fa96d2fa47", x"1e61297fdacf186d", x"51a21f9fa83987c6", x"f37fead6d4796197", x"c1924b310722e1a6", x"3c1de4aa038fe238");
            when 31427016 => data <= (x"29e55fa3aab739cc", x"b6e879de8c123119", x"64267b89bfad5104", x"788f508dba377db2", x"471f1d43d3bffb5d", x"ec4302b827e6c8a8", x"a10b35a0083b263a", x"2dba463c776ebeb9");
            when 23672532 => data <= (x"b7471e8c6bd12fbd", x"25b77526ea179c88", x"8ee7f09263eaa7dd", x"a15869a7ae80b38f", x"a2ba3e27c6c1ed94", x"a2b9439c6e9115e3", x"3bfb194f3a847f95", x"3ea23482ed27b2f0");
            when 22855995 => data <= (x"f972f1e6db51875c", x"cdc713623747d758", x"da36477aa6a7909a", x"eb9a726484269e61", x"7cc31f642948ffc2", x"5535c8c70a889229", x"6ab5ea76b5af0a02", x"fc8086aa36311cff");
            when 12577815 => data <= (x"9c5070961aeee161", x"53f661ed8981fba2", x"92efcf2b5988369a", x"b7bc91424904319b", x"31b486aa0060c496", x"1cbcbb8f39f8c10a", x"0b3520bf386a0fd6", x"bcfcd3517d72024d");
            when 5823670 => data <= (x"8d511114b4f1041c", x"1e5612bc96bd3b7c", x"d51c1796937a3587", x"4e0a082c74d8c412", x"74a1f90daa1e03a5", x"eebcd2682349532c", x"a4feb26f898e0587", x"b9f11ed6fbda9ff4");
            when 16572951 => data <= (x"cff60923a2e922d3", x"ecca5e77bb3ad925", x"8e1730b810623f75", x"42ddbf691d9cc042", x"b13c4f2d67120301", x"7befa7f70e1b3c78", x"4949de423f4e6076", x"6079d29386da0087");
            when 18765894 => data <= (x"7767f78e3b6dbd9b", x"baa2182fbf45d02d", x"faba5977f4c7b827", x"e683ac247ca29a39", x"2a2f1ce2896beb8e", x"21c410f17f2e9ba8", x"dec61ef5743272e8", x"6e00e2358e035d0e");
            when 20481284 => data <= (x"65ef525081f7c381", x"54420c79e61825f2", x"07e8c57bd4d9c52f", x"c2520aba80525cc2", x"21fce9722694c1aa", x"d4885f2929c0befb", x"7e747b09f8993d81", x"e70502998e769ea7");
            when 1996197 => data <= (x"830251c557c98b7a", x"1e14b168d0285be3", x"c0f4f4ba75521e6d", x"a656c609cf5ef8cf", x"3f2175891f08c440", x"78ce5d684af02666", x"d6a350e2f26f3da8", x"1e591f1ff3483d55");
            when 32696346 => data <= (x"094b0f06cb5fa7e6", x"32613ddc55834a1c", x"cca812295d2d1197", x"d36dcf6ce77d3a06", x"d2557d2145d1dedd", x"a399d6f377c65555", x"9ae3882088a959e0", x"f28df65c521435ba");
            when 17943679 => data <= (x"d364169f0ebc5b3c", x"e4a8fdab326b5b7f", x"df1628f18165a065", x"f87c228031693478", x"86c51697a5d441b7", x"08ce706630e27376", x"3694d46ea32fc0ce", x"2c032a05a88f7acf");
            when 26793138 => data <= (x"4b62e5090d5c791e", x"1b530e78305a6031", x"d7dd9d4f99f5374c", x"a7d5f62011bec2ab", x"0c4a4f9d60ce0345", x"0d75e524888b6593", x"156d0660008de1d5", x"e4d4aed213d7eaf3");
            when 15308716 => data <= (x"a4844937b5042fa7", x"0a83cb78de381583", x"bdaa75010bf5d828", x"c7ed4b037bd13fdd", x"2730e09e362f6250", x"e6b1782e1aef50b0", x"e0b12f371f110a58", x"c52949503edab3fd");
            when 28873324 => data <= (x"992ac6740342744b", x"374a937345f2b897", x"414b9cc81ca7aa13", x"f30e3cdb4dbbd8ab", x"30ab3469d158baaf", x"913b50bae2da9154", x"a9544e5b5106a85a", x"a04023caa1750b8a");
            when 32579985 => data <= (x"5b7c39457cf625fe", x"940e461c6b28a639", x"721d82129a75a1f2", x"99935aa9369cdee8", x"d888a894afaf46f3", x"f6dbf88271e58d00", x"dbe9bea66e932023", x"0cfe5fc4f62a8097");
            when 16596173 => data <= (x"15563efb405772e9", x"66fbe2c9d7caac3d", x"00fef680f01d643b", x"74d645c2dc2087fe", x"0bf86676809dbc96", x"287469d7adde6920", x"c72347a817eab152", x"8144fecece2857bc");
            when 19834603 => data <= (x"71a5259788d4c24d", x"5b3d28d0ba67d75e", x"bea1b2de672fc018", x"c65371efe7ee3ba0", x"a18877a0b6368d34", x"8220f84300e38dba", x"c148fdcd1bee916f", x"201b7d5a1fdd8989");
            when 30867371 => data <= (x"1803133e0edc3cdb", x"72e3cc02fdb528ff", x"a7c860cc7efe2b19", x"1841c72cd4bc4227", x"9f41743fb22bba27", x"9c17c11a9cfb66cd", x"bb1f407321b6aed3", x"fb2037a9f82d9fde");
            when 5119820 => data <= (x"5c4807ee7e6c8201", x"52cde7e569358524", x"5e05362e47263e83", x"8823784492b44ab2", x"6b6fed6f6b260e8a", x"12e492768b33fba8", x"ed796d6734fa9135", x"54bef71526dd6788");
            when 31318804 => data <= (x"cca67998510a944e", x"a0f2b11d00a45d5e", x"6e01a044d7222925", x"061b2da2f2f71cad", x"a0c43b2aaec02249", x"bf92eef211398de2", x"9575fa7cdcea3fab", x"fa24b02f4c50ded1");
            when 4732129 => data <= (x"1ff77353081bf7bb", x"4c13c78be9f86d50", x"4cf297fd8d2d1bd0", x"3a5f0abc603d5331", x"64902df386caa463", x"c2d37479f1d84467", x"feeccd6aa409c069", x"44c4ec75b7afd682");
            when 17526341 => data <= (x"61b10302299b6cce", x"31a92db2061bebae", x"460622514c62a3e5", x"9d438848eb7e212a", x"23cfe10e2a4bb569", x"8b482aee728fcf63", x"020d3f36f87d5c4f", x"ac1b2b341284b489");
            when 343160 => data <= (x"6f9ff1c0cbc44421", x"126eef8e69085989", x"352e72697ca5ec93", x"009286cf72134fc1", x"310a4d56de23fbf5", x"1c3e6bfe08d312ef", x"7f266e764711e2d1", x"9487365ab5f19d6c");
            when 25922952 => data <= (x"9b1f5043487cdd75", x"e4aa654967937114", x"b2282d8c0f683dfa", x"00092528ec4d6241", x"dec58d158147ee11", x"fdc81200bbea5a54", x"6cbe322f139d9e6f", x"2c5895f2fce13b2b");
            when 12181117 => data <= (x"a64389f58e00f4ca", x"a04ca4a1acab0f9d", x"05ced02a8b3a2237", x"224d19fb7468730c", x"f8c0fa984618f7c6", x"8c434ff76f2f15bf", x"9c9e8539a3abd891", x"7171ee02367e80dd");
            when 2261312 => data <= (x"daba9b2867ebcda4", x"e01c444485bb1509", x"e06288eeff44d70b", x"ef8348a49e2c7ef7", x"4463939bfa87aad9", x"afde91f53bb79bc3", x"4b28f0ab6301d030", x"489912c4adb171cd");
            when 23879526 => data <= (x"b2e5d82396ff040b", x"86bc3b7d5a2bae81", x"267759fbfbe09c7c", x"32acbf1c84ccb62b", x"d47f8676700b054e", x"f676536d4561d721", x"05f8f1e2b725af59", x"a7828e62046359d7");
            when 1619413 => data <= (x"c6e79d1375b51536", x"12fc1fd869e8a5bd", x"ccd19268fbf5e53a", x"36399a8935f60318", x"1b6b1ff17f23d18e", x"c42f7c0a9f88f682", x"0e6e497008b5b8db", x"e329e965e819b293");
            when 2464004 => data <= (x"941606e98ba25cb3", x"235d5cfa8885d73e", x"ae7e8fbb291234c8", x"417a5e110e2a9884", x"3b4d18f94fa0c87c", x"3b47ea22e548955f", x"0555dd4e454914fa", x"99313b10baaa9f9a");
            when 13558793 => data <= (x"9b46fae530979e5b", x"8b8f6df8d02580fb", x"c27a31c2e48fa504", x"4dbda16b8430d71c", x"2885f1b04aa87512", x"e409a7467cc87dd9", x"fdc21297121267d9", x"ab7dbeec0a2ad987");
            when 9265095 => data <= (x"3382efa76aa18901", x"6a2ec558ad0102fe", x"038d624fced59492", x"08e99c889ee59148", x"eabe764dbe10a55e", x"b514f879a2ec6f5a", x"a3dc4673c402adc5", x"8e8d1f2022048db9");
            when 9840066 => data <= (x"bf4b28872d7849ce", x"fcf5cbf100fc29e9", x"72a9796b80eb30b7", x"3a5b3c37d055e521", x"b5b4b56c5562eaf1", x"0e7ef356bf4afd9a", x"c6f3bf344accbdea", x"0a5f9bb1b6289dd8");
            when 27072381 => data <= (x"689b08dccbcc8747", x"9f1b6b2fa0a9bb2d", x"85627e8395597013", x"1ce6eb77b8ca696c", x"e081006ff494b0f2", x"9eae559f4bfecba8", x"56c0661652b9f8ad", x"617127a7ca37e394");
            when 17321656 => data <= (x"16fad2cd011e8fa3", x"aaf890ff7bb1c6c5", x"5daf25034e91ff56", x"d2510c3e5712fa7c", x"129ce13d97df8ca7", x"319e584ef7f88193", x"8e93fa0fc88b527b", x"415074caef77a21e");
            when 30211446 => data <= (x"68a0056584d76449", x"ef041d9d8ba1d61d", x"ca75dce65439eff5", x"8989021712120973", x"2e01334e38d4c98f", x"f1be482f81d92e2f", x"c19bc3a06f1bd6dc", x"bbb6ddefd4564ea0");
            when 23170963 => data <= (x"ba1898fa588b501f", x"75071975dec6f407", x"a88d90b9475d544d", x"cad7581dc7c018dd", x"3fbb5e721a2251dd", x"dcfd6e9773d861b3", x"21fb58e974917679", x"29fb568244a20c39");
            when 24506135 => data <= (x"8c25f19a16c72be6", x"d3696d334074ea9f", x"244d8a21a0ae73da", x"caf1246d613866e2", x"c2932fe264b25e33", x"d9dc7f9e545acfe6", x"1104d71172f3e6d7", x"e025241353b5f7d1");
            when 22456679 => data <= (x"22e74c18e77a2c4d", x"7deb13ed75e425a4", x"50ac39b269498fcb", x"4a390d42330c067f", x"482c2263a90ae5ed", x"ad33edad37396d8d", x"1734b42c2810f758", x"d03ac2056565209c");
            when 27098200 => data <= (x"848904b1faee4058", x"98dd2b26967843d2", x"ff09d6013309d057", x"12c196aba9320d2e", x"e324303f324e91ae", x"672595b7a1f7b80e", x"4b85ab33c8343392", x"357018e6ebb664fc");
            when 7191860 => data <= (x"da8122bc9f95d050", x"e9c8fea6f9ed5e3d", x"3139ee5885b77eb5", x"1fd887d8783e1497", x"c88272ca713fefd9", x"2f91dab5209981ff", x"c8f5942e50a94395", x"1f419fe56ab0cf08");
            when 21907722 => data <= (x"30a8f652fdc689d1", x"47706703d702a87b", x"076bf294ff1b2a2c", x"2af1c96dc04c3c83", x"82aaf67939b762f5", x"e2ae9f353975cc57", x"7d1e3587404cf657", x"a90097dc3069fc4e");
            when 15204899 => data <= (x"fdba495ae9dc5d9e", x"847aa7aa3220b2ab", x"9d764f0ee04746dd", x"bc8effb8209342fd", x"101a7b91beece3b3", x"d5a91ea93fb3ad5f", x"1b061ce99edbdeff", x"c4197ad2a30c62f9");
            when 16916731 => data <= (x"70da0ae34baa19aa", x"dbd9e0d35ff0f13e", x"c9459994e7cd4c01", x"b195f522d6130eac", x"5242e3c0025e943e", x"b76b802d83287ca0", x"90c33c36c11c7c91", x"578f71a8889caf93");
            when 30572414 => data <= (x"a706e4ba755c3ed8", x"3acb348feb3ba505", x"f8cbbac356f309d0", x"0745e12e9f86be8d", x"69885baa1f07c993", x"1d90b44524e7ce59", x"39268360fab93247", x"7e6d735cfaad7eeb");
            when 28954175 => data <= (x"ea1c7d968d95b3d4", x"b7469f9bb8d53289", x"9515fe90ca6d4f4e", x"bdd298c80d592ee1", x"a9cb2cd704a04666", x"6373b1a268b71001", x"a3133803703edc0f", x"a12833bb5306a5a4");
            when 31114540 => data <= (x"255b75e5cd6b32fd", x"af52c41919ac3622", x"e94822f8e2fa518d", x"d533ca952b900914", x"e32a7f809ea9de24", x"f5a441900a02bb42", x"8ee7b061bbf36793", x"e97ef1b26e070b2a");
            when 4200276 => data <= (x"bd28e306a0704c43", x"a467f8478b1768a4", x"1023ee98b0a187df", x"d280957c5148c7a7", x"e3df5fc773cdaf62", x"8311527e8c1cefea", x"6d922f716a6ae140", x"e206cad88a9b9db9");
            when 25447028 => data <= (x"5b9dcd2585aacba5", x"320b29ff12025314", x"979515d10caf3cd8", x"77258ea828919527", x"bd76632ce507c58d", x"169bd35e48b3f9b1", x"25668b3a78e9642e", x"86fa5923708b0813");
            when 11235368 => data <= (x"6335744eac243d3b", x"e4ec6e050aec1c51", x"8c80a8cbc99c3dc0", x"e49cfe6a39288fb8", x"17af0aee994e5bdd", x"bff7917e5f713b51", x"f38f832a412b157f", x"96270a5e4d8a8513");
            when 19581433 => data <= (x"7c7d15c857976dc0", x"09d918d50d0275ca", x"ef2056f36e9d364c", x"ee1a4a19126aa366", x"0b67a43094623117", x"52f79bb931a35ac7", x"59741b02b75524c8", x"34eda9c6ba41e06a");
            when 12701742 => data <= (x"b5e1d7faff92948e", x"b5bfee790e0c11dd", x"8cc21b2c0eab049d", x"4705b35ace456de1", x"e2947ef362ced1e8", x"7e6de9eb4a7edfb5", x"a5a916b3d5dbfe91", x"8c9bc684c50f5577");
            when 8751728 => data <= (x"7532650aaadfcccf", x"a83776c61131417b", x"00d93559eb13e2e4", x"3cbc96cc096fdf0e", x"e31197fca369f142", x"f618876c74a1eb5b", x"a0de15dfc811b419", x"8e2e007eb933b10a");
            when 5687307 => data <= (x"d32b0dead636e0cb", x"ea3230ed6f435d40", x"f87603f4bee3a508", x"441de40a241f6d5e", x"38d08306225f4d54", x"882ecdb88b6dca26", x"197f02ae22cfec0d", x"8cf4c50a0a85bbc4");
            when 7066678 => data <= (x"a9b1e5c57ac5466f", x"dc9cb96fbae37914", x"8a430ede3393a842", x"a1a55c9fa4187e0f", x"f96922b785f2d31e", x"bae1647a4a47f9d0", x"894021ab40b16b95", x"4cf27d7ecd1d9561");
            when 4719475 => data <= (x"47d7cf087883af48", x"49a20f327c29f776", x"0f2839343e3e3dc6", x"c02f09946da498d1", x"bcd87f5275d26ed3", x"c763fc4f04512be0", x"4ad3d2c7f7d14763", x"4c3c5a40f9db5e18");
            when 650912 => data <= (x"cd179f53f1efeaad", x"248cf9787b875948", x"552e2cc4a84c0fdf", x"8934ebffe5963faa", x"3c64c4e0e2cf81cf", x"49aa882629da6bf8", x"a92644ad162a793b", x"66cc0b975efbe7ca");
            when 1022184 => data <= (x"ba64f55696c07742", x"08d0c72af7170379", x"274dee21919832c5", x"3daa442fd6b8d595", x"c6df5bd913adda29", x"e7d8f4d40c60faec", x"7800e6b51a106c8a", x"4d95bec684c36245");
            when 33516570 => data <= (x"d33dcfea02102e3d", x"b10f86a3f14bf125", x"cd823f236d1c9eca", x"1d15a4d6c349dde3", x"b8493bffb0744f81", x"6fad0e72e028d65f", x"b21f51c397ddf835", x"7b99516b00585ca9");
            when 2086560 => data <= (x"78570fbc27c14566", x"0884aefb826a3889", x"86300bc94df78213", x"a7eef60533ddde93", x"38fbf7719b84ae42", x"256c9fa574c193ed", x"47cb391a1b59c9e2", x"6ba3fb048644de73");
            when 32800891 => data <= (x"ee7ffd85448ad819", x"c8f6d392143a3839", x"7383c02633de82f0", x"4ee4edebb3559e9e", x"48c6cef5a88d390e", x"9ef4e0ac67683f00", x"6e06707434d16311", x"fc58f12315061541");
            when 32423744 => data <= (x"792fd98958fec18b", x"0db795259df25610", x"3c61c65be57a4461", x"f202cabe74f97e90", x"c067b8bb527c624a", x"b86e18f99048376e", x"4dd09af05dac5d76", x"48c5d1954dbea82d");
            when 33214493 => data <= (x"c009e155c5c367e5", x"eba4024536af7df3", x"3efef9d80a9b2c3d", x"997ad5604e67c693", x"9f07c166f2fc250c", x"99d34b5b830acb22", x"f59794c5475c7fc6", x"885216ce563032ec");
            when 6046882 => data <= (x"04c491716fdf0c1c", x"56c1b2ee8f0e6e15", x"e4f3214ab9ae43b0", x"29c094718c57da09", x"e515b2596638f095", x"8d5300d586078dac", x"1276f4e0b57357b3", x"c935799430c42fca");
            when 30942637 => data <= (x"02e7240ff9abc64c", x"be8b343ea220819b", x"230064728e9c9ea6", x"a7449beb24184302", x"d8ef7805221be18d", x"e8ff0d2bcb9a93d3", x"6d017d050ad09e6c", x"fff86a0487f7f458");
            when 25279910 => data <= (x"6acd364f779c2328", x"46c696eb95e04db0", x"05da186665248f0c", x"306331f3b275f83f", x"bf54d1c4d2305466", x"ee7fdc4bef0de1e1", x"107563a227fc0e85", x"2dd2cc6823bc5b83");
            when 5719631 => data <= (x"39b4575e1b5ea884", x"5e563f7da02d63ab", x"2398065775d77bba", x"0aa79680faf0b878", x"98d12d39a66c0fdc", x"67a94ce1101840ba", x"3043597e8cc528c9", x"1d9ba80e47cf9159");
            when 20687155 => data <= (x"609ece808bd401da", x"eff1e4b8aa8be703", x"19490688f2537618", x"420a29ac22389c30", x"9f785297f1205841", x"8a93c3263abb7743", x"06d9a15f7997c4a0", x"0c1add9c95b53d1b");
            when 29992672 => data <= (x"33614ee0bdd45ed8", x"53375a906f9fef77", x"61d0926c13f0dc26", x"3a42a4f73e3920d5", x"a803633c73040aa0", x"ffe2ec4e27576d27", x"7a093a68b05f783e", x"5cf346efa8dece58");
            when 21565098 => data <= (x"0b0ef6fe3e27cd14", x"4cfa5b3b8e2b9efc", x"a96bab932e5f59e0", x"3882835ec66149ab", x"670cfb55d0d907d5", x"1158e29bde07e83f", x"97416220428a33b0", x"55c184e2b0d55a1c");
            when 7109345 => data <= (x"162bb63fd2c62510", x"8921834572375448", x"832a9e66d5b9df4a", x"f528a57899fe7a35", x"df1ec9869d3000a3", x"a80e8bf5c3c8b20d", x"8793444eee51e213", x"f4b4903ed2abbeb4");
            when 32466022 => data <= (x"418b22581c28f81a", x"eeae587fdba1b2cb", x"c87ab1e4a144d2ff", x"498eaa90ba354545", x"39c4e4a7f6be3737", x"163cd7a2ed33fa0e", x"56a4cb22931bb4af", x"e122f370bc826875");
            when 21312966 => data <= (x"54d50918dff5433c", x"ca5a2a95f0c182e4", x"649d6b1c94cd53f9", x"e649fd3010f80f5a", x"db32567a0d19ddc4", x"78c0cd6ff9cb253a", x"303722007ea0e937", x"47eac6d7dce25485");
            when 6411142 => data <= (x"96c15a29d398236b", x"215545afe2a49f41", x"47d671b073fc378a", x"95703d6b7ed603e2", x"7f42d342766847fe", x"53917fcc8a0b0a27", x"a420d33d1a1f4d8f", x"8e6117efcd5149c5");
            when 28232041 => data <= (x"e2493c4ead8476b3", x"aeab41cf5be89b7e", x"065d6d514634a95f", x"5d6f6c10ea5f512b", x"68d0bba80cd51d39", x"402c7c0d7290f576", x"774e5e10ee985b71", x"b746ae81b979fe11");
            when 28942891 => data <= (x"646cfe28ac320886", x"b4bbd490608daa1d", x"ca28573f7eba1048", x"dda35bc169c314d8", x"559922ea29ec6f9f", x"e780ea7d00a9b946", x"f3a0e3d6119ad57f", x"e1b6bfb52bc81132");
            when 6098804 => data <= (x"2b75337d90fcddb7", x"ac99e74ee0783df3", x"1d4b462cdb9c194e", x"fd57c1362a5e9827", x"a4a838cc16f3d240", x"ed8df35e2d01f168", x"006a200eb7ef97f9", x"eb5a0422a33433ad");
            when 6916841 => data <= (x"ea76a9319ccfd780", x"7586b409fada56e1", x"bc2e61397ea5d3d3", x"07db689892437586", x"587f2042e014d208", x"abf6b96266fe174b", x"1becbf6f98ef9b29", x"84ce63e4ec1800bb");
            when 12604954 => data <= (x"59a6bf1a7810ba61", x"53703960796e1d11", x"88eb5d315c3fe456", x"e71fc63d5b2b69e8", x"9a0d0e94a637847c", x"f95c5ab487c773ca", x"74e0c1717548adc0", x"9696b9fe050aa5c8");
            when 28622364 => data <= (x"358afea5762c512d", x"d82a8661ae939925", x"355bb17d3f1e828f", x"4b964f76b015bede", x"12354c5aa758e1c2", x"7263801ad2f7e724", x"69ab72e8ee9fc6e5", x"8f5ddbfaae781e5d");
            when 28466287 => data <= (x"b93d5bdd65f90a5e", x"f8b43f0a686d0734", x"e8d04057f7712d30", x"c39c3400da701a68", x"a0d9a0f008f137c2", x"4ad4745053e8cb5a", x"acd75144bf732e0b", x"2b1bfeaee35a762e");
            when 31859753 => data <= (x"2a706d6e6cf57b4c", x"f2ac6ab70556895a", x"e11a358cb9172719", x"3aca9d0c98e073d2", x"0d1d3b396502eb62", x"9c8d5407de39fba3", x"d0d5c397717a38d2", x"10c3a21244bf20fc");
            when 159064 => data <= (x"1a8fad43c7a139d2", x"772aa322444d2899", x"50de62eace23b12b", x"66fa287cd2cb8a4e", x"ad0078304bf33208", x"85742e1eb87bed0c", x"1dab0fc9d1379d2e", x"5b511d8f135c32f7");
            when 4847221 => data <= (x"88fd3ccc94137df4", x"b4f897c5d2cbd9e8", x"6a95d3ab65551161", x"0b7fe4c63a29f358", x"ba484bc16dab0f14", x"e35d2bdb1925653f", x"132f33d8025e6c71", x"a4e4c90d5374828a");
            when 26045205 => data <= (x"5feb94c71e9c0e78", x"005d01225dcd6cac", x"0c86e130d755589a", x"dfbb748d40380599", x"8407354ecd59a227", x"896781f0ddfa1041", x"571645503e857b8a", x"3f0b6a5dcabcb5ca");
            when 14565870 => data <= (x"a4b294492fa06489", x"a136439bddcb850f", x"5533b45f438f7cc4", x"eb1cd210e73cce6d", x"7f720833ec767d7f", x"6b2135e740795d02", x"727ffde3f14d71f2", x"59ebb897836e22f1");
            when 30834102 => data <= (x"45d78f550721e285", x"fa2e269e6646d5f3", x"6fdf0d5a2714ec10", x"d8aa84af1c842635", x"119d2486a2b8ee92", x"446151659a1bcd80", x"7c10cdadcbe41e74", x"c67dd7d567529179");
            when 11018895 => data <= (x"984335ed94105097", x"7a351acc90aa1c30", x"8a97060dfb94658a", x"5ac1cff7966b385a", x"1a7cf57396b286f9", x"2a6da05b157d3736", x"276e574223a91913", x"e11b8b8257c5c309");
            when 2230742 => data <= (x"d3b40a5747fbb78d", x"07a299f512a8d6af", x"99337046a147bdc5", x"2e176eebe987ee90", x"332bd7d28af1f449", x"e0a2d91a0c7d01bd", x"2db95917080a7792", x"e6a6867c3b5ec1b7");
            when 1495307 => data <= (x"f97c023f1d60b88b", x"f58f4262b21c63f3", x"89f8651aa483726e", x"fc5008a7b19c069f", x"5cee82684f8c0b3b", x"471b1d4bef57b41f", x"cd63f947aaebc927", x"b1a7909036941d6e");
            when 11777159 => data <= (x"f575efda530b194c", x"be65bd71fb49f3ea", x"2a07ad27b1c3938b", x"5ce8a3a88a7c5004", x"86f279746572397d", x"1a42c06bb4e77390", x"23f1dae9b1ec3399", x"00d38739472d3a42");
            when 18667769 => data <= (x"8f0738aa8724f969", x"e876187c8f25b0ba", x"c5dc8f2c7d7d80de", x"fec1574347e5c33f", x"b6f958bdaff976f0", x"a2ebb194204b8ebf", x"2b2f8e50ec7e0b4e", x"0a2411723e5af5dc");
            when 6277778 => data <= (x"2c257d35896a60f0", x"b0e5e1aa4674e7e9", x"09a21951464ad4ac", x"0966530e8d3f5e56", x"89c8a07aba555a24", x"484ad8228e042173", x"4522828c13cc63e3", x"ccb9eff2ca019599");
            when 25947603 => data <= (x"d3b9b5f5a04de18e", x"cc01c16a353d868d", x"9e99df7a2378c1b8", x"2c23a12682b06775", x"9fe1b469c2b8176c", x"f3a284b84ad1fdc1", x"446a99ef9f824fbd", x"d0fbb3482bbca51a");
            when 21341267 => data <= (x"1b5af7cc5c1c8333", x"17b3a6c4258bccb4", x"ba8a42d2513b923b", x"e7cd99f708cacf18", x"04c4ee23fd8f8a2d", x"dd000095c2631c90", x"30749e0f65ba59b6", x"5abbca3fdcec1aae");
            when 11984343 => data <= (x"52fbf79737f8bc70", x"3c01c8eefcd9fea1", x"068c3af9e5fd4444", x"1aadc1b98b274ef8", x"f65f5e3780dc1ac4", x"3e4789a45a1d83f7", x"f595282bf7b3c9f3", x"373cd7649f4070da");
            when 23922020 => data <= (x"9786748fca0b82d3", x"a06a56cdbd6a4660", x"55f643addc5b0244", x"5c6e495f4259eff9", x"eb64dc40a677937b", x"6259f9f6ef389e13", x"64a04a29718d92ee", x"04d4c0265c1c4d55");
            when 1762049 => data <= (x"73b30c62bee654da", x"89ee62d0824e32d1", x"332cb754e9a62ba0", x"e3cb690053a2791a", x"40246f7ec6000f4f", x"3ddf170e7fb8625b", x"e6304d3af3034f0a", x"23d66bc73285c38e");
            when 26574638 => data <= (x"8e54836bd572623c", x"d711da0a0528facc", x"4bc32f92ecc8e16a", x"a0e821e85d633f06", x"5f3566d0364d3431", x"cfd1fe6e4faa90b0", x"a9b7ee325f0eaa76", x"4967cfe3ea287483");
            when 369327 => data <= (x"e02d4167368fc061", x"b908e22710904999", x"81fb7c1486c8e75b", x"2f36f24361b5b120", x"8084afb1f9650327", x"8a0617c47e7d7035", x"af2fb322e9a672e3", x"e26d654b407782da");
            when 30308734 => data <= (x"878de691c6dfa3f2", x"16351e7181875742", x"f308f9e2f30f223c", x"4d9e738d481a6b0b", x"164804e17151a43f", x"1a26aa874bb14c9f", x"76fdbbeef310871c", x"c1b62f9f16c90a38");
            when 27077825 => data <= (x"2ebbe54773019fa3", x"738009cdc5688422", x"f70af039c22bf93d", x"8e1e81e81c7b7d73", x"8b2b701d869c97f9", x"4bd1eeb9ce1ddb1b", x"03dee3c74834bcc7", x"b990d0237f90dda1");
            when 11013451 => data <= (x"05296f22fcd6dbed", x"02acdb8e2b1442a3", x"5c3f0b30a57cac39", x"5f0af224fd464a03", x"d2b2fa600487e24f", x"8779ca3b2c13febf", x"fcabc5abfb6bb4f2", x"7ae2a4b1447149f0");
            when 17796139 => data <= (x"b1631f83634f58ec", x"da2117a40403beac", x"d5d9355f7d991fb0", x"d3f76616cd3daefb", x"467869a8fa2bea2f", x"1cd5a8238fd1bd82", x"6fb4729cb5c8addd", x"97ef461a8d0ce6f1");
            when 32230349 => data <= (x"86884f328feb05d7", x"c27d140fcca955f3", x"18a27007f45fc43d", x"93b1e2ce00cfc66d", x"2de91113151862b6", x"2ee4cc8b0cfe1b25", x"2ecdc2705245601e", x"18a4ad2510e9138d");
            when 12743934 => data <= (x"f6bcbb5284727f3c", x"ba506825d0a83ed0", x"5835920a06fd4cc1", x"67a9c427881fb136", x"6d09f5c86af60b80", x"e1a7a41c1449727b", x"db2fa42cb9b00127", x"a6a0bc0ce5daffdf");
            when 19578839 => data <= (x"c954e988e1e229ea", x"b71b6fd9553950dd", x"923d99c4675a985b", x"480d42ed38673299", x"8d25c0c28b66243b", x"a247f1c87c962ddb", x"f6fa7faf01ff0bb9", x"16f213f7fbac8a9d");
            when 2321884 => data <= (x"b364296d59da6a5c", x"a2047a8c0af2ed37", x"54b6505466774e48", x"ed3377f0d2a13185", x"12c2e246821d6cfb", x"4612e8c5becad55b", x"c8e89b81a20f1df5", x"374f75cfee254bd6");
            when 22322512 => data <= (x"4db11d43578aeff1", x"b738a9f7d78632f2", x"536a7e58ac4c4db0", x"c5875e96cee3fed2", x"2df79c9564dc57b6", x"bfd416c6ed57ca2b", x"6d959c7b28cc5c91", x"2474c7b89d164fa5");
            when 27451865 => data <= (x"cd9086c621a3cb01", x"831d33ad739e3b4f", x"fa07274491959aa8", x"c58b974adbc5bb00", x"8baf0bfff8aabac5", x"13e37e5aa37204ef", x"3b616894319e5d39", x"099b3535ebf6cb46");
            when 13973799 => data <= (x"889370d9694cef51", x"a5542bfb6276ab86", x"33af449e408ab14f", x"8f33566fb3ec82d0", x"476133401f7606d6", x"aac684a409dc4cb9", x"eb84946c3effcf4f", x"f0f9b0c02f313f9e");
            when 7641922 => data <= (x"20c73c20d99d4407", x"7cde64578bd59389", x"696a6ed7dce6bd5b", x"8976ac9ccff5389b", x"173e9869e9b38a71", x"f0c4b4d5ab7df78b", x"32d52232ad975f82", x"00dfaa0f014efe2a");
            when 29491199 => data <= (x"2c230c7f72308d8d", x"421b531146fed57f", x"571f61c6e3e49f6e", x"2fffdd8c66e9dbd8", x"32f2a6e5323d0d2e", x"e99ac0f9f5ba6a03", x"388407c8353bccbd", x"0e6251989e17f9ec");
            when 19194991 => data <= (x"f175e724967b26ea", x"524f115ccfec708b", x"5e3528e8076ad2eb", x"4943ea5d0a7ca42a", x"375b81ac3c77d996", x"508e73745219f37e", x"ad7c4cbe9f921da3", x"271b94f2082b8ee3");
            when 19030845 => data <= (x"82368bcb11c317b8", x"052666e1c1e566a0", x"95f0e8cedbfd0792", x"945b5d2830392e52", x"7e9004747faadb8b", x"a22c2295c848da71", x"8a14ebeaee896a5a", x"987f8bd50a451732");
            when 22299727 => data <= (x"a8448e31eed93beb", x"2ca8546756739b23", x"6ff49d8388bc1e91", x"b16119a4ecf968c5", x"c6da5b44e0ff5168", x"67c360790af6c97a", x"bc086470cd88a3c4", x"c7e32c258001968e");
            when 14113622 => data <= (x"77e8caab0e953021", x"fe91f1148b96efb5", x"b97f4e16b59791e8", x"437db379625b3e19", x"0f8c5930d36e8e46", x"4ef692c7113a9c73", x"32e84fe4f115b702", x"c1e80708e368243e");
            when 25819067 => data <= (x"13e4ab95c27326d5", x"a172ca575b16d3f5", x"80ea3e089dca6902", x"7c989af17255d2cb", x"d148e47756215116", x"e4dce2248cf67287", x"49e9986e0cf4174c", x"3563ba9122fb4a93");
            when 15343466 => data <= (x"08e62b795c031f50", x"1d2e692c1cd0f1ea", x"c4584493eee04f61", x"dee987b2e353d7c9", x"4d05e375df9c68c9", x"d2929e59d3374bca", x"e27aed81c63eb267", x"4d7df8a64fab5321");
            when 19643313 => data <= (x"e9ae629cbe715306", x"c6337c91351f9fa5", x"ee21d6353b0bd2ff", x"d9bcdcb73e3adc53", x"b1920baa4948e954", x"ed75e8cb29281e36", x"ca46b66929588e35", x"e22091b0994abcc1");
            when 847029 => data <= (x"8e6771a811c0037c", x"fcdc80207af6ab67", x"492811630063d8d8", x"ac28f2b058b13f56", x"94723af1f8b2bf26", x"f7ec74e31604ba39", x"36d38c78a40f5f46", x"00a161a18de0e39f");
            when 4212023 => data <= (x"39ea6bd99d40badc", x"abe3fa0ce8fcb563", x"779467614c0574d1", x"86e233d90290907f", x"474297fe86f62529", x"f9002b36bf619172", x"2562f05e46569e42", x"87607813c52c02db");
            when 2176831 => data <= (x"2215c433b9eb893b", x"a208e7e2ab38fce6", x"b469efe06641faea", x"9896124c99c110c0", x"5409386ae5ff6b68", x"080ede4dc9e54dd5", x"b55235f0fa69acd6", x"d9468a80ef536dd4");
            when 27043435 => data <= (x"62d4d80da9e3ce95", x"3430d25c1bd81f43", x"75b395d2bbf2284c", x"ad9cd965f07cf3ac", x"a1f2f05a7f1355d7", x"41054f3da8feca06", x"d2c659988a6b1967", x"852b27d2a4c300a9");
            when 13060725 => data <= (x"2ca6c67dfcd68b3d", x"6d04d2591279ae79", x"655b6df93133d1a4", x"af43015894cd92ae", x"0d9e694971cca38a", x"125f5b0cebd530b4", x"abc3b5edfbe801a2", x"e1021e8404b9598e");
            when 14287608 => data <= (x"d48ae616fe6b5e28", x"f3ecd203b003215a", x"7bf43437e99f8400", x"09d5cc7277ce0c75", x"1ea0bd4041d2d31b", x"07dbd07e09a40541", x"2f7c39d1b4671529", x"6fdc5f0164455b4f");
            when 8939568 => data <= (x"db7c978caa11b24d", x"fb22fe3eec477153", x"4d28933d0e0d1deb", x"a4839eb5fd2bec24", x"0a21f8f6b151e418", x"d3a5912bca6138ce", x"f999af695e6eafcf", x"9bd956b9788a3fe7");
            when 28094343 => data <= (x"4385df98f3bc1d57", x"232f720e365203db", x"d90841d517c789c8", x"d22fd1e5d247fed3", x"b231e5e81eaa47fa", x"a4d2bb4d05dc80ae", x"78ece730f15f7d43", x"679f7014c814a6ce");
            when 13192102 => data <= (x"7f6168270af6b4e0", x"2d34685dcd64ef7e", x"732bc59e1607e995", x"d49dfdb2c857d27c", x"5c88bd72a825d49c", x"b14d0f009e91d9d0", x"e185674c73eea958", x"11caa45bb3f7afe3");
            when 22022163 => data <= (x"2ea21f0aee0fa3bb", x"0a43cc3a90148688", x"88f859b96552406e", x"680d31322efb6226", x"48c9506a5433f6a1", x"0f19a4df2461b662", x"64b12ff4e4204980", x"d03784a78ea6239e");
            when 4652000 => data <= (x"3f63369be46167da", x"51d25b8daecf991c", x"4a35adf0a213d595", x"dc3c29d46080caf8", x"f4068888ebebc374", x"586c7121fcd79ddf", x"3e13d18bae4801de", x"2aed0de5b46ac60c");
            when 5477283 => data <= (x"9fd66e58f7b28f89", x"d1f614b897620647", x"b8308c99a7d200ee", x"4d0cf355928aee6f", x"ef01e43fe489b190", x"36ed5ac03f90fc37", x"a599d37e7ba628f7", x"609b4553fa89cf6b");
            when 3826753 => data <= (x"c1377fc8903ee241", x"0f1d1541e0baaee8", x"8f981428a2829b14", x"b1e2a63238f0bf71", x"35b4e01c6585ab0a", x"a3e74767d389d1fb", x"bf0a47a9d88b3c1b", x"57138154ef02450e");
            when 23969596 => data <= (x"03e81e41ce7f9182", x"dcdd7f0d47a13c82", x"a36516ffef56462f", x"44825bfd0dd5c1d9", x"8ebaf4e5504c55f6", x"5cdc5b7198d80507", x"e7a349e6b2620b75", x"0484739d3510b362");
            when 5745374 => data <= (x"c64988238d4734cc", x"ce9bfac21bed9370", x"6a901e45a5672e54", x"68ff24daf526ad27", x"ebc31fa81761ee43", x"15d07c861a1a4c59", x"3538c762265ddde3", x"26ff7e83516d582f");
            when 7690584 => data <= (x"c074b51f4f586945", x"5bb3d6d666b37dc5", x"34f01855d9248d36", x"9c56b2c7e4485cc1", x"f51bcd7929c832c7", x"14a898f643af8b2e", x"8ac62fe222287842", x"ec99782e17f1af35");
            when 19325426 => data <= (x"ba419d988e04d6e0", x"14a1bd9d9dbc43ed", x"e3f2be4d48becb24", x"ee0ae59d789a30ec", x"4e9a9869d13a7b92", x"eb91a0d718f3b976", x"9d0f2be5dd1ff047", x"a581d95138048635");
            when 22503508 => data <= (x"ec3cd119198645fa", x"dbaa4d125cda4318", x"55f02d493a6df8ce", x"eb712b294bc27232", x"435d9657b702220b", x"b81f9df54764afee", x"19d8731209582054", x"5484fe0aff00146a");
            when 31152063 => data <= (x"6bad0f018b5459b6", x"212c9615258cb81e", x"89d18f7ae7645c56", x"9496c15d6af34b51", x"e189cfd7529f4061", x"39c76dc43585fcde", x"44c44b9082f13392", x"4a7e355108df71e7");
            when 20998677 => data <= (x"95afacae55f77434", x"34dbee029a5d9f22", x"79d74d4e7a2afe57", x"065ba7ef44f374c8", x"18d6bdfc803c624f", x"cdf7d72d7bc8ffe2", x"047d1f62e27b8975", x"e5fc5c414c5c6cf9");
            when 33164248 => data <= (x"28d5b57ac24923da", x"233af04584bb457a", x"93488b04d0c67e95", x"b2f1021bdfad637b", x"652b81b5ccb1167e", x"3aa7ddec10ed0c80", x"a49830d7a86417a3", x"7cd83021578e6174");
            when 14776529 => data <= (x"bd2cc2b0ea0c6d46", x"8e543e6f12d80be0", x"e6f1f3030a568287", x"d43402ff7223b7d4", x"3aea37bf915bc0e9", x"177d8e1202424c1c", x"9681f40bbe212dc5", x"d25013233360eb63");
            when 11945625 => data <= (x"6ca06e393fdb447f", x"b26ef46df4990095", x"a85bd61598650581", x"06b8d144a4a678b7", x"f46bca728f6fde62", x"dae3972950dca2d8", x"8c5e0fb3f155471d", x"e64a5f04bbbbedbf");
            when 25077332 => data <= (x"8114245facb99612", x"18a0d771d6d0ef2a", x"151b3e94550a4c7d", x"fc9fbd82288c44c1", x"cfc01a6dfb4dbfaa", x"22ee515455aa24d9", x"81cea20f5917e9e3", x"5161bf1db07f178a");
            when 11572017 => data <= (x"ccaeab9ce06a3e15", x"9dc58a6a95a10c4f", x"a3c5f1c892f82d32", x"e95ca01debf6cca1", x"418dbb4c8ee76834", x"ef53b1138012f5da", x"d6bd6949139987f7", x"6a0e83858ea71107");
            when 3426571 => data <= (x"e75358f2333275c6", x"684cb538cf93b92b", x"cdc4210908439024", x"ad865815ebd51911", x"93235ab7f2442b08", x"2255abf7286dd145", x"fb713d4e21e3c142", x"45e66a3610006229");
            when 16956272 => data <= (x"78c94419fa9d105c", x"744f8561dd3d9de6", x"b9e7ae2c74701de6", x"1a2849e5cf00815e", x"be3ee40a413713fa", x"796647fb2c760899", x"7d778ca664b765c9", x"055dde73000c12ae");
            when 3274070 => data <= (x"39cb141b4a14debe", x"b988b9364631bc43", x"abb97680b73a8f28", x"9546f9e2d5e82a22", x"48a94bcd66ed95e4", x"47c8f22014f3b593", x"c81a2f10213a7eae", x"61222bf8e690e98a");
            when 10422066 => data <= (x"faa4af86a918594b", x"c85fd48546bf0c9e", x"ad2bd1ab0d623c2d", x"749240bc633ff595", x"359eb94a8c999181", x"aafb9d16890cb049", x"f33ec7ea04c71784", x"8d24ea5eff0dd851");
            when 2850957 => data <= (x"b0a0da24191eb38f", x"37857e5ff85e6061", x"780f8ede705b1ba2", x"71afd83b63fd5f25", x"c0076628642d0422", x"ab92ea1c994a7043", x"a0a6f9b61d83fc06", x"23a4ee7e25907ca3");
            when 23786539 => data <= (x"c765214479f8012f", x"feccdccb4fc4063f", x"3dbefc43e0a1d1eb", x"c2ea2ac57ff0e506", x"ce29fdc0f5535778", x"8f345a120b47418f", x"7291cbee29e64c46", x"a3d58cb5c9e711ea");
            when 3539532 => data <= (x"8e62c688464bee3b", x"4de2b206844b215c", x"34390decf64a762a", x"af00399ecb672d6f", x"c93eeee54582ca5c", x"d4c1a45e30f12969", x"057289cedcac9fdd", x"bdf28f08de65e798");
            when 2489291 => data <= (x"70969cc206cc2259", x"c3676e22c7bfa1f5", x"ef7df1e309177742", x"138758db3c4fdfff", x"80bb0aab63587aca", x"320bbb15fb95db97", x"4dc5100e80e77d95", x"be679324e0dee673");
            when 4043043 => data <= (x"7f8673c8485b79e1", x"49a17f714088bb9e", x"e9a7427efe017e9a", x"278947b193318849", x"e76bdecde294768b", x"1b6834bfc7d7ed0c", x"af9f789bf4a809a3", x"4b67260a3f31df6c");
            when 16239709 => data <= (x"f1c86a062abc7f42", x"b8539ae58e869081", x"9af97c20f9502d05", x"9b60498a22881571", x"59cadbc7a8b5fa15", x"263c35415ce52ee6", x"07612110674d81f9", x"237f098407a774f5");
            when 19730729 => data <= (x"00d4f6326c771d80", x"1ad51c338358864f", x"d94c394db8bcc09f", x"da9bb912278f0b34", x"30e3d2baf6124688", x"86edb42c267d7c15", x"7a0d4dfcd0f3d0c8", x"bf318c6c17c657da");
            when 33355560 => data <= (x"f92468ff2d2bbbdf", x"ee3df06bcc8d5bb5", x"f5fe2ceed84b613e", x"51c677067d1ebd8d", x"893d8f6fa30a3a4d", x"e634d9b7a3d0ba2d", x"246dfa43a176062f", x"2dfed9c01859606a");
            when 2903171 => data <= (x"3ec4e7e014ec1065", x"7580d37061ab2b18", x"301bb14c8fde60f4", x"3a456842f5cc94c9", x"092f375e5301cd7e", x"33701cf90554cbb3", x"771845a4f4cdb823", x"44b1e932b14b66df");
            when 15265319 => data <= (x"f83eb366540a96a7", x"fab3a4d5233fb540", x"5835913651cfec83", x"3ae045854ceee80d", x"1906bff3df7326fc", x"61bcb1a231cafa53", x"13096111570e5b75", x"f798da4b3476e086");
            when 22297274 => data <= (x"877984ed5740ff20", x"0060a75a3c710674", x"21023e62879cdc5c", x"8a26002d0dd87b52", x"08f9dea7268b3eef", x"520c8dd6b577e74a", x"aff1ee0dc34e609d", x"23e2d7d1e44309e3");
            when 28553339 => data <= (x"0223c0f351020ab1", x"f01871fb180575ae", x"48368192c7ba3b6b", x"123f7020e930d752", x"b6657cf3e6f0abcc", x"4b09678bd65695a5", x"b1122ce6cb416e7c", x"84e30f083a81b5ea");
            when 5039219 => data <= (x"2ed828537c02febf", x"30c5b349621e6c60", x"c6e1e054d2634248", x"ddd8ec28a5f6aacc", x"61d389256bea78ef", x"b380de9f97755d06", x"2ea69b72ea254ff2", x"9c08b090bc4b02da");
            when 6735844 => data <= (x"86887e27caa23f65", x"1dc432efe438316c", x"d8e644eb6b706b15", x"72f97879ece1cfb7", x"51ac54653e096d9d", x"c7131ee37e4a9aa0", x"1e305155320b47bc", x"c00b53f49442e6a0");
            when 9834155 => data <= (x"7969dd643e919271", x"e5dfd58e18a24f85", x"4d8e6b4dd34b428d", x"fc6875c3691b4705", x"3327cc4e19747e90", x"c638f1ad341c9dc4", x"5bed1a0affbdb0b4", x"2e86c3cb0130cdc8");
            when 23832064 => data <= (x"64b5c656ac77bb53", x"6524ea19b0ade60b", x"143e3e82935a584b", x"51eb6428994ce76d", x"2f2c2fe7ac02ce50", x"326edfd7d90acd2e", x"d88993e403682178", x"09985112b7e0907f");
            when 32776316 => data <= (x"d7459fe340ab8b3a", x"8459ebae5fbd6916", x"b8904146ba08ff71", x"185337f66000bc9e", x"4d5ffd4aa4199999", x"b22342056cab3862", x"a5400a969180ea49", x"9e152797424a3c0c");
            when 23473597 => data <= (x"8e45ede9abb9f758", x"224fb24ea75c5ff4", x"834e6c7f5f20c300", x"aa5dd1231d928544", x"47fd40dad6e0033f", x"81ca33e9742f1b13", x"b97ebafe268ae270", x"48508a8274ee525a");
            when 17453207 => data <= (x"13fc0fdf8f7963dc", x"fff43252535e8565", x"58d5403b678c24de", x"0ddeccc080ad6817", x"7639fc9a0789e625", x"ff856dabb392ba73", x"452e349aa18c5a55", x"8f219bb42a71af80");
            when 27021489 => data <= (x"35bee206d577d54f", x"dc2b9bc36021e7cf", x"37d1614d5590b165", x"2128e333541fcb61", x"18d3cd6d32416b2c", x"7308f97b34539438", x"bb1d1ebf4e520a97", x"848056dbb76980dc");
            when 27950583 => data <= (x"0cd9e457df99a0a2", x"3defebb07ac8ff9b", x"7421b23b32965df8", x"37304d3bbcdee41b", x"43d07222e0fefe0f", x"0ae9668364b3a895", x"85513e8f2cb2dcff", x"edffd68bb8d3373c");
            when 8175282 => data <= (x"984b296bf9371c61", x"85ffcccad2bb3933", x"5a254605813f789a", x"9ee596d87b9d9db8", x"7a943c7310a4d9dd", x"fa9104bf49ab144d", x"19b716d84af2d41d", x"7096590a80498a05");
            when 14170808 => data <= (x"1fa6bb33d40251a6", x"602b5e99a6b3e0c5", x"3df58764e2f7c1f9", x"debb81cd617cf569", x"f742c7c62137d99d", x"acc9deafdf51c2ea", x"7b53f7899298c8b6", x"24bde1b98488ffcd");
            when 16735655 => data <= (x"593fe89ba6ef3252", x"971e74bdf208897e", x"896144903516d43c", x"8633a45c45147ae7", x"26026ee20ea83348", x"d7f90a86efdbb25e", x"ffb3c96619aee4c5", x"de3851ac5c4e4934");
            when 10834102 => data <= (x"a338d59682d8a01a", x"45672f9325fc2109", x"9d9c70f97f9b7255", x"d28ae63898007fd4", x"e3f6f2f30db9575d", x"41e04ecd36a46fd7", x"fb0bdcce1f399f43", x"b3bf73ab799c148a");
            when 11215508 => data <= (x"0de0ff944f56b34e", x"22eccd2cc711e41a", x"d73966445dfc61e7", x"663602e310e2849d", x"b0b63211958340e7", x"5634d8806080cd29", x"52a521c7779dfeb0", x"63526d41a7ba97b7");
            when 12862149 => data <= (x"9f9fb9118360461f", x"6c6306ddac538491", x"2661f51d0738238f", x"bcb54c1cf2c2da21", x"e3ec5a9f26302910", x"259abf504b1d42d6", x"7d1e473e174dc619", x"ebdb342600419507");
            when 7677885 => data <= (x"e997104ba4483755", x"b74b5917d75d8aa1", x"b52ebc18e579d96b", x"0dbce12799eab3fc", x"10667ae1a0546337", x"ae28d58f82dc9746", x"4c709e9d83829e4e", x"f1368c3337d00e53");
            when 17763338 => data <= (x"dfa2437130c92923", x"0268f83836f8d870", x"ebdebefb2ef16c6e", x"1625507d2ebddff4", x"51c1032e5161c169", x"c90006e29ac77bfd", x"57bdf7fa729464e5", x"4d7eee9b0d4aa4df");
            when 18106455 => data <= (x"8bd1eb941aee0120", x"352428480ab64ce6", x"c1d09d79aec54876", x"6dd8b90af765c41e", x"42e56c3a1db2e6c1", x"1281ea3e899a023a", x"7f3dfbff5c4f55db", x"5520e3a0eeb2dd96");
            when 27076337 => data <= (x"4828a3b5cfb0919b", x"48465c8b8445acca", x"f6fdf9144547f1e7", x"6bb329ce47ddb908", x"a1d3b8d13708860c", x"0327a2b23eed0c36", x"10df70e251dacc7a", x"63717435e8ac21db");
            when 4898498 => data <= (x"abdfdf7a4b47f618", x"a16a1b94da978a71", x"97a286eb34854fe1", x"b76e2082f1565870", x"4081432b43308c2d", x"df12acb95a448f26", x"4e51391a5d030e3c", x"1a7ac36bc5ac24ac");
            when 2394184 => data <= (x"717c26c05112dcac", x"cefd264fad8ff239", x"e601aa54f3eb9d17", x"e72c82758d0ea992", x"eba83acd3f6430ab", x"04f11b174e571be9", x"49c6a16ad22c515d", x"a3cf745161584ffe");
            when 18544917 => data <= (x"00b079be70da2a4a", x"3379e7ccaba3b4a1", x"aa811cc6d5faca3a", x"d16a3ca830a80b64", x"d0d286c69187075b", x"2f3516d280ebb22a", x"49bd45e91d325637", x"8c254f50d0340a8b");
            when 15139391 => data <= (x"2d9f8b16c87d92af", x"56006b85534e9319", x"1c883600fdc7e014", x"b7c2d483aba8f40d", x"9718a739b6c7c474", x"b56bb2f6d2d4e5fd", x"7b71731747d46843", x"8b8bae6ff6102694");
            when 6516709 => data <= (x"44e80c62964842ec", x"2a20bd67584252c2", x"43bcca0680195821", x"756720a67da14d7b", x"620ccb5dd061ee60", x"246b41360215f650", x"467bc7cedd142229", x"a91ca377313d0149");
            when 30174631 => data <= (x"9f22b7c3b3e109df", x"5825acfacee9da11", x"f1374107dba74ee7", x"aa801a1983368577", x"2749585084d82dc3", x"ad17d6e340dd8070", x"71fe7dd21a1fa00b", x"75e57e0ee6563ef6");
            when 12422138 => data <= (x"63a24afc37ce7e92", x"d8685cb80dfd1bee", x"5db15599d5c6eea8", x"4b0d3553089c0080", x"13b4c8b98535f61a", x"2e969c5c60a42090", x"802941c22526af40", x"2dd56fe0cd90244f");
            when 20659888 => data <= (x"1f3c8a8b5e483b04", x"3ccf213665330dc9", x"35ce9ed60d0f8514", x"9061373cde8cb5a2", x"a1fd885f35016412", x"81c1e22aeed9fab7", x"78a11db7db5bbcfa", x"969f91e9419f08ee");
            when 4242331 => data <= (x"6bdd7440f0da4acd", x"d28f752ce3917274", x"1b3fb2fd05b6ae84", x"b865d652f7dbf699", x"8adc283d3999f0f1", x"6641db74e55e80da", x"5b0730427b95a341", x"d52ffed66a076985");
            when 26605841 => data <= (x"b11e45f4110bea3b", x"cc29a9ffe8513a5d", x"8d752fbcd41ca495", x"eb33b94218d0559d", x"d66838130e7c18de", x"ebdbb748c62390e3", x"45151ec60b95453d", x"d0145fd02dfb3845");
            when 10767039 => data <= (x"07dc08d211cfcc5f", x"ee99c5372a720b0c", x"e1fed70066dc1e3b", x"aa8275e98346c27b", x"9e47b3098453eab2", x"30700599250f319f", x"8cd1f6800ae12332", x"06f0856689da4408");
            when 12951867 => data <= (x"0dda165fc8a2e8d4", x"3970cc777275140b", x"05a482d36dff739c", x"5cc04110868ddf74", x"50f7206b11b3aa3f", x"96b8df7a15e7b64a", x"e3d064003aba1dd9", x"0fd7017375384d14");
            when 26986283 => data <= (x"8cfc692c32a30430", x"e4aa0c901befb77b", x"8b2faf36d113b0c3", x"3ae2be0476d82947", x"922eee20363c8c0d", x"b45ac14f60a0ac59", x"35526d1d91e902f2", x"4057ddf852b8fdda");
            when 8520155 => data <= (x"fe8ee59b63319c65", x"d8123fff0abc83fb", x"33b59f7ea8a7528b", x"d52589330d52b58f", x"e5936788a6e3edb6", x"8e98c7b1e5fbbd84", x"b7e56c5c16d972d8", x"8072a549306e246f");
            when 11781424 => data <= (x"c0b1d7cf865ded9e", x"63b7ef1689fadb77", x"77ebc1ca4cb4ec5f", x"c1e461e6d7a421c1", x"8dfdb2721274ba9e", x"265b2526b2d051c2", x"533bf8bd19368e39", x"a9126041b913c980");
            when 31255122 => data <= (x"f1248431f8a6112b", x"d84d53854e8eda3c", x"3f1a61686b4d2e44", x"7d9c3191f311c835", x"fde495a9a436d304", x"0ea04c37bab1233f", x"ec391241ded4a760", x"c73decba0a43573a");
            when 2245637 => data <= (x"6b35b5b7e5cf54b9", x"2ce8aebcd501c1e8", x"dc50085cb73b32cd", x"cff287ca73b1874e", x"87fed9e50bc40c3c", x"bc2f2f5c0c4e4a7d", x"bdc73a6c35eb7513", x"af5ca10682618ed7");
            when 10148004 => data <= (x"5acdea1ecd4d7d0e", x"ed7641254d541fc7", x"b87d1e70cefab384", x"5b0dc4a3afa9841b", x"780a384d2aa2e5ee", x"4c2f06d36a4a2d02", x"be5aa02e4644e946", x"5f5ad3bfe0b89a5c");
            when 32247111 => data <= (x"edc0b59655dd0f16", x"18b5ca6c7225feb6", x"409c9d893bc9c8ae", x"e38aa4275b2a18cc", x"d7d836517994a6c9", x"aadccf95bfdf3d2b", x"4f4adafb1bfee2b6", x"de6f2f85d5b9e643");
            when 2126705 => data <= (x"dfdffca3a05421c1", x"8e1f0ead4e8432b3", x"9b9db99fb7ea9b5f", x"96be228d4ddfe39b", x"706eed6266f868b6", x"f0e75d2d76fbca5e", x"075fbe54a61025bb", x"53386715f253723e");
            when 16422561 => data <= (x"7819ca0f5bd0f592", x"7dc8f361e0c6901f", x"cf7a071cc0c06bf4", x"9cae2c6f17b05f19", x"d746201d1830cb38", x"8419fbff98c6d6e6", x"03ce60ad0af9e69e", x"def41cc102c5f0d8");
            when 28861539 => data <= (x"0c0f0e42a3245946", x"a53a22fee70c5936", x"594472874655570d", x"6509a0774c252473", x"560d60ebde309d30", x"bf7428563eb2cafe", x"ab2c72ff4e28fe7e", x"eb0e92ab1ce1da07");
            when 21613509 => data <= (x"7088bea0be495884", x"430fbd4ca30ee015", x"005881feee9084d5", x"697e6ce02fc58e9e", x"2ca30c7005bad5de", x"6ce61d3fd42c47d1", x"26928629bfd0aa5c", x"a0657fec4dd8f7b4");
            when 30809947 => data <= (x"de55b0bea3626c87", x"172cc04e9c43ceb7", x"7bd864f7ffa49d87", x"32844ebd0f21f2bf", x"24d199db2441bb85", x"90d3ebfcaa80657a", x"b2112054d8a538b4", x"74cdd6481815d029");
            when 33183112 => data <= (x"cf1f32120e06983b", x"45b55279e88ef64a", x"a80ee22fd6b72d83", x"5b5b5036500616d3", x"97ad153a88b2983f", x"f69f5d195ea64cf2", x"4abe6d94b106060c", x"6d5a8e75e4d5192e");
            when 6285525 => data <= (x"f27c97303a3eedb1", x"30ca8a37d6cab5fd", x"21dc96ac6720e2b4", x"0b3e78519fb25941", x"d803abb85ebf3150", x"9aca02006ad688b7", x"498636acf769af6c", x"6f4482ae890c5115");
            when 21666110 => data <= (x"cc0927d5b7494a58", x"dff54078102b51bf", x"645f0d4e9214c51f", x"8895340b7753d2b3", x"abad82bb47ca441e", x"27f6b71db8180699", x"42ca1e0b69f016b2", x"2235c1aec9c23799");
            when 18594107 => data <= (x"b9fa90bf909b08b8", x"73a6411c1d33faed", x"7fe4b58cdaf2c21f", x"dfc2317bc48f4f60", x"dc6e4195cb0a35e2", x"c47e9f8b6e5bec60", x"7811d729c3bd5a20", x"36169d6f21a37c74");
            when 4674844 => data <= (x"95edc8d9c49e43b3", x"2d4e33b993e78435", x"15f5a9e49f9e0454", x"aa04338ff88d2db0", x"0931ec616397f7e2", x"7570d7f813cfefc9", x"bae8bbc8db825198", x"63485e8ede9a3eb3");
            when 7136991 => data <= (x"a3669d6d83297aa6", x"054211d1e2e06809", x"d3a00cf5b30d53db", x"0a3bb27fca74d601", x"e38cba9bc82ad58a", x"ab3088d91c232873", x"763f03bbeea9813d", x"6076a7342e94c0f9");
            when 17168314 => data <= (x"dfd89c2c34e36116", x"ad232b20fea7f240", x"e104bdeaf1513470", x"de7c222e4566c394", x"c239cf827ba890ab", x"28ae5ba8b85d13e4", x"240d78e6d896cf6c", x"a9ab4e075e2bddc7");
            when 24662795 => data <= (x"ad97dfd56b4d708b", x"1732bd92ca178dac", x"9d2b739c25104478", x"2df8b70e0d4e1b9c", x"adf8e0897089e70b", x"7cff9f784ff56afe", x"ed7b568376f433e8", x"7a46c0d9c6bd7ede");
            when 16928730 => data <= (x"66fabbf60a7ba371", x"950daa166d5360ae", x"7cd1bf8e2f210e04", x"2b6719284037ab68", x"f320354b481e02c2", x"9056167062a61d80", x"689010bd7b86117e", x"8b6a60a3e4f599f6");
            when 16851352 => data <= (x"a51e260fee5204ad", x"f7de0b1db76331bd", x"0af66e0a974da8d2", x"6a5e5a4cea8671e7", x"2aa9fe822e80aea3", x"c16236726d1d0aa4", x"f6f682c1ca9df49f", x"efceb8027fd7f050");
            when 11251499 => data <= (x"4468525fec294a9d", x"ecd53d11a3b8b49d", x"e3131177ae6472b8", x"2e6d63a7a374246d", x"9b4121c7596ff413", x"90d896fa946e96c2", x"481772dd0d1dbd22", x"5bf4a61601c0d765");
            when 21667 => data <= (x"c19b6c0b2bc1f596", x"d016018058a7df41", x"1df57f1bec8a55b7", x"09b5a600570697d6", x"51891ab12693bb8f", x"e74f893bc4bd3fda", x"63901ec46d998fcb", x"f64381798c721b26");
            when 11265602 => data <= (x"5c9ff8b94bdc635a", x"7b000759fe1e7d0c", x"15caeed356d48d4c", x"08647d04660307fc", x"d813daeccb8c976c", x"5868d79e1e5f1f73", x"297161473e5b50ff", x"25f6358df771d95e");
            when 16389855 => data <= (x"f351f43d531356c8", x"6b3474133f796b57", x"0a1a29e245fb78c7", x"5f50bf145feebcf5", x"bfb0230bc409ff6c", x"58db812d0d4dff39", x"2dabc1f5dddf2dfd", x"4a9e612234ea74e7");
            when 27902516 => data <= (x"b6ecedb8a058ba0f", x"42b2d746886b96bb", x"1b733d623a5af479", x"665bc964bb574c95", x"439e3e80ed10d9ef", x"245c93f4101aff8b", x"f4e385dd90e496df", x"17e92f634e2e7e29");
            when 20519375 => data <= (x"ebda8885e53be21b", x"235cc0659fa98e8c", x"0a158c2e0b98bc89", x"137a1ba7f5fba1a3", x"fbd9dd8f51a34289", x"2c157b655b63e8a7", x"779d0a778934c75b", x"7e0d6437f210ecba");
            when 12104053 => data <= (x"f2aa4f06c759491b", x"d308f7d8de8026b9", x"bf32d0444defa70f", x"0208fa0cef15823a", x"33d47db65043a1fb", x"98da0c3be1db2e69", x"7c9b0d08f1fa5a7c", x"77e296158078f837");
            when 1344327 => data <= (x"1d1f8e0e5c9e9132", x"4b9ddcda6c22e407", x"4f82fba61ad47b98", x"2e2be3421006f0ec", x"22c598e67a3c93cf", x"10a2918e7c70af9a", x"a8fb110bb9dc4e08", x"a1ece5f720ad82c2");
            when 31663326 => data <= (x"1264517fd1deaae7", x"e9d97e6c8fcd771b", x"0ee314c00ced5e18", x"b37a8090e7db611a", x"ae07a29147790e93", x"5fa36cb271a14352", x"85c88510e8db896d", x"8559fa5d2ff32aae");
            when 20346336 => data <= (x"52ea4d3d3a23d912", x"557fe3c4b1feed81", x"27e0569bd07275bd", x"b38769f3673e5a31", x"d8f83f02b2b2f592", x"ac6e6e6fa199aef2", x"07ee1f113b16c8b3", x"1fb02e13c32b74f4");
            when 27596173 => data <= (x"43411e69998c2517", x"4f3ff7c36436d8ae", x"e9d84c0f5365fa1d", x"38ccc280cb79f65e", x"2a36cdaad113b62b", x"2afec39a104c4c3f", x"aeff1b978df29ff9", x"25f5b60947dee7f2");
            when 26216041 => data <= (x"6eb0083596d1be4f", x"ccfead5d3c14499f", x"d1eb0138249fd375", x"419b5ee5d0648a14", x"8849caab8344aea1", x"2305f3c1ffedc248", x"ea566302f7fce99b", x"2ce5ef299fea15fa");
            when 19042714 => data <= (x"b47b6882868c4bfd", x"95dbb9ba0e433e21", x"2b99a84943953d5c", x"ce7413523ac96385", x"07a6234e2f95f661", x"581c634b0113fb19", x"5af0aece7e5f8219", x"ff59d0b18efeaa85");
            when 26608840 => data <= (x"810e6bbb76845f3e", x"7eb334ba8ed73eb6", x"69417b395b8607ce", x"e3a0932ae7487ab7", x"0d49965cd5426fc7", x"149171dcdb9cb402", x"16d556807d6fe901", x"967401ad894b27a6");
            when 8423331 => data <= (x"c2b78b5cc8620ed1", x"7c9bccdd81e1bfe2", x"ff368c6ae35f543c", x"ff97e542f20105a6", x"7260053a9729cf98", x"c75766d8c78ac872", x"67495d2b8a1aaf7a", x"1bb4d1c87d9ec8ff");
            when 3340081 => data <= (x"60f57790a15f68eb", x"e609f6f5d4763ff0", x"1ae4664a8a360e68", x"9317df969e001c73", x"34d2616a98ba661e", x"5dc08689a96c687d", x"7a15b294693c11ff", x"fc97c9c35445b83b");
            when 24177009 => data <= (x"5c071379a893e3c3", x"d380341d7b87246b", x"568d7c778fb014a3", x"b7911c3d5eb30d58", x"6e6639ceb1947221", x"86d3d1628bc79ace", x"68c2f2708bef527d", x"50eac71ecb3319d4");
            when 10684982 => data <= (x"f422d5f3f2bc46ea", x"021952ee17c9d477", x"1f853507dc3783ca", x"09833ba75c1f5c8f", x"f41543438a85dbff", x"8d8da4b15f3a9022", x"b7cdc1746d8da7e5", x"867c628abcaa2b88");
            when 12241327 => data <= (x"2f5e8fcabb44df55", x"e476814355814995", x"15e4a29f038b50e1", x"4538d81980209bcf", x"2d179854a43b2f7f", x"8c47eadccfd40f10", x"4b2d46349f934d70", x"c5919a9e0c30b10f");
            when 6872284 => data <= (x"a6dcf38a5bf19044", x"c5c3d9406f52bd4e", x"83ed46dc9b0031b6", x"b9e34f3dab560e0f", x"941cb10d73582c60", x"7e4a01ab6f1cc48c", x"f2b4f0633373f8d6", x"b88e961fd1fa95a3");
            when 23189824 => data <= (x"af0d256a01fde33c", x"7eed01521133687d", x"ed1c45927dfc5840", x"93c3e0f6a5859a87", x"4007f7feaa625be2", x"1cc35712f6fef85f", x"1ac26e0f2195c1ad", x"f10da52b2e26d957");
            when 10421024 => data <= (x"a4898a8a9706df43", x"672305324af942e0", x"b0ce31291cd9f0cc", x"f31051c7ed706f56", x"9533589dedb1520f", x"cf3f030a5b934a7a", x"ff7c6367b011007f", x"064127246611087f");
            when 27363842 => data <= (x"73d2e0a56e53b831", x"6d77e352cea8d0e9", x"c0c3c710c5ac99e9", x"e09922b35201653d", x"05b97c9253d63af7", x"b02007f5356535d4", x"11bcad6e61589b22", x"3520b2a47ea4fbd5");
            when 26480663 => data <= (x"2579ff57589732d1", x"8ed17dd584586187", x"68235475c028ebcd", x"ec3ec20a21b14bb4", x"0370ee1bcd4ca91b", x"3ace50ff4ed26f7d", x"92473239391641c2", x"02289250b0596ff6");
            when 7558019 => data <= (x"e5c66d3e2db884b9", x"949e357d34986a6d", x"a0609311abd2d0c3", x"b39672b601766cd8", x"b4c950587ab200f5", x"7ca989bb80eddc78", x"af9bd1abd6b793a8", x"3583c6ded930a102");
            when 9922015 => data <= (x"0726208dcaf3434c", x"2b460f0cfa774eac", x"549abd6834981a52", x"7245690b4e89c007", x"2ede67b4b8da5a2b", x"e859f2b4230e09ab", x"89a7c3b9c3efc824", x"fb166ddfb9ab743d");
            when 15701833 => data <= (x"ad27147e3764efaf", x"165cb76f20ff14fc", x"6e842fa4806b0853", x"5e3b0d199998806d", x"36cee22a71c99b53", x"a31bde6cedf2ed8f", x"138bfc82a3bc3153", x"236bbd20da9d28b0");
            when 8999968 => data <= (x"ec016d004dcc10bd", x"749a5481f7744d72", x"761546bfcc5f4a79", x"de2efc985f9cb3aa", x"339b02839295ae19", x"bb268632cda4c0f9", x"4130bb0c71ba6794", x"7d1e930e96976f36");
            when 13142211 => data <= (x"94739e7a72e97d64", x"f15b61ae69c90b36", x"b7152e6f90319106", x"5aafa28a583b9559", x"1f888f32d812c66f", x"840da8908eb9f177", x"519ee10a32f1fe25", x"d44f68a065120fd0");
            when 13154583 => data <= (x"ddde231325263e72", x"e3088a5edbd0feef", x"642024d52c3ab04d", x"fe75dadf210df431", x"c3e1f5905d1e5438", x"9c5856d4fd9c14c8", x"a372d2227c2cc0a3", x"71092bd96788681e");
            when 12053599 => data <= (x"5a33e7412fcbd36c", x"2378b2e0df6d25d1", x"748bbcad0a7955fb", x"61faf4ccf2576ece", x"931925610d3e1786", x"3d7753355a13e8db", x"de1b6d5d84ea2964", x"7bf02cabb07ac42d");
            when 17449064 => data <= (x"767bcf6e30ac419b", x"3a00c1aab8845680", x"093d42c0b481d4e1", x"1b6e3fdb56fc1d54", x"7ec71db05dc67856", x"142f5d9e31dbb93f", x"21be756cf682e6c1", x"4f592f7c2f142643");
            when 17020545 => data <= (x"ca0dee371a3b91d5", x"a844877622278741", x"6353e9401d281767", x"e076724b846f2510", x"ced4d26daeb527cc", x"93bc7dcef86629ba", x"9607b00c7d27d0f1", x"5a64424078bf272e");
            when 3433310 => data <= (x"2232d3a5b9141b31", x"cd86611112aaeb8c", x"5a505d52b81dd0e0", x"05792002dbdb433c", x"aa41243ee0b2406f", x"81ddbd850ee6cdea", x"b6e557738fdfcc29", x"e6d266dc5039b81e");
            when 14849329 => data <= (x"793891ffdf9d77e1", x"ecf2d386c968a2aa", x"064bf06443c0b56b", x"cc8a85520083ecd3", x"136636e7f2162dc7", x"9420d1a7897ab797", x"40472da5e3856325", x"52bd53eb02d29d9b");
            when 24936720 => data <= (x"9140c429e660dc39", x"1256d8235466e924", x"c035c966f380755e", x"d2407c0c46786754", x"b969e662979f9388", x"f7fafe7efd4e5fef", x"73cb0bf56d389774", x"06f4417a49da5356");
            when 2304864 => data <= (x"80a1aef4e7cc3283", x"bec6177c75839ca2", x"ec99cc95dfd79e49", x"72117752e0f1a2c8", x"c83914ab7df7f086", x"b841606018203e9f", x"aa99dd4a61bfc0fb", x"e14d2a3ab8941b21");
            when 2658668 => data <= (x"195624e19f7125a7", x"e1a1d6a68d200a9a", x"ec64961649fc2562", x"faba4b57afca6469", x"96b51510dd116e0e", x"9fd7c04da92ed1f6", x"f6b1ce3347829d50", x"1ed96cbd03a9dd55");
            when 9343351 => data <= (x"1d23a902a506ea2b", x"98969dbfb471b7c7", x"21bb310452cba3f0", x"e170ddfc59081934", x"5f19c2ef8df2b20b", x"2f18f985b6313f79", x"25ab7d0c03e18fe9", x"6ab4917a0e9b0932");
            when 19803997 => data <= (x"cbc6c4491463c14a", x"fc4a0f97618d3391", x"e8f16c27e5c0e7d5", x"a6c8c3c1e40db155", x"d575df6dd8cd3545", x"bfec0915b1be7272", x"fb99c93811c8e334", x"4c7ac04ecebf0cc5");
            when 11474411 => data <= (x"95a616c7974d2f10", x"b102192cccc8f9ef", x"d57bf36df2292bbf", x"3ebf67b6545e4e60", x"368a9c812a1816bc", x"0bab54503bf2e8ad", x"db4e7ad03c2aeeb8", x"44cfb54f6bac15ee");
            when 28610908 => data <= (x"89df50f8b2d4daf1", x"b3c76769a4502a2e", x"2181c77e0af17f3d", x"4be188f4da3420fc", x"1ecb6603b135c92e", x"42a22dcfd42cc8b8", x"e97ce4accb4696b1", x"13465ab33d65e03f");
            when 1281315 => data <= (x"b80efbd8728ea826", x"8d5279256041d4e2", x"17e5637596d3d596", x"de94fdb9d0b8d868", x"663e8daa768c9275", x"c785c26c54851295", x"4b6252468fc7d049", x"1f354a6e30b0459d");
            when 30707130 => data <= (x"7e992311ee768663", x"9f5c45db2ce84a6a", x"7d020b4140a63d28", x"7156a0bdf30a91a5", x"a66eb5bd3b77469b", x"d04ba405716ca484", x"1a42d57f39e74d8a", x"1aa1f0aa09cb7853");
            when 15642543 => data <= (x"3170066aab1649a2", x"6a252200204ce90a", x"7c84090578427c71", x"8fda6e9ffb41bbb9", x"92339524374f6ba1", x"4419f342a9218949", x"d3cdfb20c09c60c6", x"9c8af40cb134fb35");
            when 3107479 => data <= (x"943ae1871c19eb5f", x"b8518f59ea5485e4", x"953e4d31ab8be289", x"a593f5ce0a76c62a", x"781cd7e2979c223f", x"77eda7b9dc48ea28", x"aba178445641eaa5", x"2786cd91be57c91f");
            when 10737158 => data <= (x"9e7fa5aa16f149be", x"43962f6191c1a477", x"304059f0d34b920b", x"1e4e40b40f2e3ff9", x"69597f575b18d84c", x"1a2c629f77672887", x"06403e50f89c8a8a", x"981d3cfd025e85b2");
            when 13083251 => data <= (x"6097201b72454922", x"9818744dbc15780f", x"c9804195bfec4bfa", x"735187194381e473", x"e551ad8644efa461", x"a674c48d696814c8", x"0a9749af54510d52", x"d03921b87a695697");
            when 5260545 => data <= (x"5fdb12afd8c3a1dc", x"c4c1dcaa1f504f77", x"18e69492be486195", x"4d8c97d74d9ce5c5", x"9602f73bfc1a53e4", x"95ff195979772709", x"fa28243601504bef", x"127c4ad550b53265");
            when 32639763 => data <= (x"1accfa9afb911746", x"1c75f168600c15f6", x"0fb624477fb9d51f", x"359ab7593495cbff", x"6d4c9ef716956ebb", x"90bac667239fb29e", x"89e1f25c76a96c33", x"767b16259f09a98c");
            when 23052926 => data <= (x"cbfa38882e8c0a45", x"abd23cafb9f07701", x"59c5eaca27721bb5", x"75b3b3903631aa08", x"906ce118c5ab6704", x"1de7128893a5f0ce", x"9c482d93d5535137", x"191183cbc8ef44bd");
            when 11315145 => data <= (x"2d9aba4806556dd7", x"b5741a7bf4af8c4c", x"a311fad103e098ad", x"05f7dbcaa01958d1", x"256dc33b18efdd06", x"4552963c083ebf27", x"7ecac037ccb39b30", x"08c15f6de838398d");
            when 19113181 => data <= (x"b3d2c2f3da7e7fb3", x"b7dd2ef38b0cddc9", x"68cb10d51c5717a9", x"08e7f0b6dea54dab", x"2e442a8e010c365e", x"5df8ea83d00b94f7", x"8bf0afa8fb32b516", x"8ecc1cc452df95b2");
            when 30641807 => data <= (x"7a1cf756c1524594", x"fd495d85a3a6dfc9", x"4ebde62ce8f00148", x"994465102f09fe81", x"851e2c0f95313158", x"9019d02022b34a60", x"9df5f8710736d584", x"63915e43504a856a");
            when 4917652 => data <= (x"0321f5dc1c7215c3", x"a1e18a996a821df2", x"a318e59db7570aa8", x"868bf1958610230c", x"85d36e41415480c3", x"64982b70ea354793", x"2b32b7ebb85ad792", x"06493cbbdc7b7985");
            when 10245686 => data <= (x"daae2a36ac99b3b9", x"1112f2312c348e03", x"51e8baeb1376765e", x"f47036a7f0a3197b", x"f5480d74488a9695", x"c7eedd6d269285fe", x"bff453eaf5e01cdf", x"ec63f0e3616a81e5");
            when 5075801 => data <= (x"773e3aef9a0a4dfb", x"4ae0ffab5c266e93", x"417698833e3ab642", x"88caba91d47348da", x"d1e268387567210d", x"e21f887f8cbb48ef", x"9c8cc3a5a2270375", x"b888aca134d573ba");
            when 20502709 => data <= (x"4d6ece535b419bc5", x"043ed5fb90e1cef8", x"74fbcbfc600515e9", x"5379de81e8d89dac", x"c0dd772a074d09c7", x"07bf922b0534c498", x"606ba426e75fb0d2", x"6d86cc63915fb7d1");
            when 20274382 => data <= (x"59299e06987ffbe8", x"70a5fa96f3d0638c", x"2c5a19e53f9ea47d", x"775660e9c3a1f86c", x"a5c86c0e5442c6eb", x"2ca30c21ff102c05", x"7d736f5a61d8ec73", x"0f5bfd47a5e7725a");
            when 19318154 => data <= (x"5b10cc364c750e40", x"90ecfda02da39fb7", x"a014a0a3e34dc6e5", x"04759935b3ee77d3", x"f5cdbe914f7d1682", x"aa0fa11ae0941537", x"77babd8bbd8d5916", x"a21ff1ff924384e3");
            when 32474485 => data <= (x"a243ed205a72267f", x"fe65acd515acc234", x"df57ffbfe414ef22", x"afc9b871e61d1fe4", x"95f734f463ef0f4c", x"fea585e6da2e42c2", x"399c7186a0926aa1", x"ba42bd5f5debcbd0");
            when 33008009 => data <= (x"a5c3041c9e16b574", x"5ddab11a5d039398", x"e8fcae68f90fae3e", x"95fe88b7ba9172fc", x"16dc3a1b3f3ef1a3", x"2459c9d740196992", x"c70d483845b86f37", x"299511815c7df2be");
            when 10138174 => data <= (x"5d6d375c8b837713", x"78bf6d47be9302f7", x"3169cdb969d66dfb", x"77a117321e0930de", x"6f86b8259b41695e", x"7644797345c7d2a4", x"664a99cc9af438f4", x"fb656ec78324038f");
            when 14959336 => data <= (x"9f494ba778079528", x"c0c83334cb3310b2", x"d327abc751063605", x"00eeeb1ef0a61d9f", x"99111594d42ca599", x"348b951a05cf9733", x"c9ec0ae97e77bc6d", x"d88b6dad042a4cca");
            when 29130000 => data <= (x"da8184fd7399bf5d", x"0d4fac978f6a2c4d", x"32f8ca356bf49f85", x"05bcdeee32ed64a3", x"153faedfdede4166", x"4e1616298652d2ed", x"3a45a510696b29dd", x"44287d4b55043023");
            when 17842898 => data <= (x"f8aec68dc6703673", x"a607386b0fc6be98", x"5a2a55232f68e718", x"ccb9e6bacc80b043", x"59931e6d354f2b86", x"0a197411dd3bdacb", x"d7ef08af84d16c32", x"0e9442f7d9afaf1f");
            when 224589 => data <= (x"1ec9dc0225e5fb5f", x"43989cbde3a8ab87", x"7b9ea668c9b7dbbf", x"e04643edf38240fa", x"280b19ff5e6dc4db", x"f433f0f46c5e9bfa", x"36d7812e40b084e0", x"fb6975e05b0a447a");
            when 10208083 => data <= (x"a0b3a0b5e05eee5c", x"0d33df52900bcad0", x"ea31d20d0bc12993", x"93df26f2661c253a", x"95413de8d2255430", x"af2ce6d0f2c91e66", x"48f3192a6ed0fdea", x"49e23e9ea4071049");
            when 10720382 => data <= (x"c6eee68820edeb00", x"570a14ab5ee53116", x"5bf6ffb5abf5d98b", x"cf2c30453cda6098", x"4736e662ae4eb089", x"c9274b8240ec429f", x"c22263154bb2f1a3", x"c3bf3d67502ffbda");
            when 5534413 => data <= (x"7923e267f5918430", x"5b224e93428e96e2", x"0ce23f5732680c93", x"cc444e6d97070271", x"26e70502c18d73c0", x"869f84480a8b9a5d", x"e9e9d4c877cdd5f7", x"356acc9798257a4f");
            when 31331218 => data <= (x"ceaecc13a6304f04", x"62582b511bb5e437", x"e48acb13e2a64d36", x"ce7791e6c1a5a859", x"4a65a9a8ceb97849", x"430d3153af5f58dc", x"1381b59dfa4eeb09", x"0903ad95a2822532");
            when 12724675 => data <= (x"f1892ee97d1b670d", x"43a70321eb40c909", x"88f5b19477402439", x"f598b0330ed038fe", x"4b591afb1b0bd834", x"c61d2f086c4df7f0", x"5e44a4c6192a29f7", x"618ca54cb48ebc5a");
            when 16997334 => data <= (x"a4dde333ba6d8204", x"8ea352a51c72ef39", x"aaa16bbf375a5ca5", x"b6298182dcc55ac3", x"f9a6c3c739de933b", x"74ab3e39b0c726bd", x"850011af0c7472b7", x"f988cb88d4a8b8f2");
            when 26649161 => data <= (x"6666a2eb824de247", x"057e9f84f08404dd", x"bc6113b359f8d69f", x"2d194d4202bca6f9", x"6e61ba04557518a8", x"3ed60ab5688fefbe", x"69659050836c76ac", x"d8c3fa055acfdebc");
            when 5961498 => data <= (x"09f8389cbb22898c", x"2e345d6bb9663eee", x"0819e5c6b1af9ea5", x"491e2ae75cc80143", x"acd08cf97f1eaf0d", x"781fff06b8950249", x"85a58d70c9b7f0ee", x"e2f9025bd1b3455f");
            when 17084321 => data <= (x"2977eb76f7480d38", x"6464dae4055abf1e", x"d0fd21fdf6048ece", x"6e56f7384df0d393", x"5511bfafbb1e29fc", x"0958f50e99fa5ce1", x"0b2b7822d68bac97", x"4bdd4c8c8116355e");
            when 2836701 => data <= (x"90655f9383dec884", x"129ef516e81cec28", x"6fe12b95325cc95d", x"be8381cb4384d6b8", x"3375262923f0d9f8", x"32cb8ae28af4fd43", x"d91d9bfd181b9a7b", x"33bbd377891d5259");
            when 11185352 => data <= (x"db1b0e023f797cdd", x"0a741fbca849a745", x"688aef6791b118c4", x"323e26d2dec2ec71", x"869c55edcd3dce60", x"cd4b20a2c52afbb8", x"8b6080d3e28add46", x"4b3d48c8e212bda3");
            when 4736970 => data <= (x"6628eb5b112efd10", x"1f731c5858d7d33d", x"6f6ec48cfd4f82f7", x"3b9801202585b6e7", x"cdf8ee366a79d462", x"3386ef00a31a2954", x"eee932c116a6dec2", x"a5ca5c4c0f02b005");
            when 31888135 => data <= (x"65b5f293db9c67ac", x"1fdae3edf5562044", x"cc6fa0f5e6d3b2bb", x"56daa70383d2a0ba", x"d1c186aad4be50f8", x"cd86c796bb55cf77", x"a01384ee256df609", x"f4fffb9536d2aba7");
            when 27759473 => data <= (x"ecde0824a92e82db", x"a2b651173fbb6ed8", x"316c0aadf6b99abd", x"4e0898ef3764fe70", x"b4b2f7d0dbee4360", x"7803ad007533f8aa", x"18ee319ecf6fbc74", x"2803fd9d6215fdf6");
            when 30353828 => data <= (x"e36c11819ec4aec6", x"a4e7574e3ec8063f", x"248635b3bb993ecc", x"a510d0210b89cbc8", x"3ab8735929570c04", x"ef6907d4170ccd53", x"2d8f3c0c472bb97d", x"9970b7988d35c978");
            when 7851448 => data <= (x"3534f6e7f7c8832a", x"14bdb29384c47e6f", x"869ef2501700917c", x"f5864eeeac4a2cd5", x"d3d9a801c0200d07", x"d999b1827dfa679d", x"5569447356b4bed2", x"71a101c12da50fcb");
            when 8561852 => data <= (x"2ee6f57fb344b4e2", x"1cd6ef4aa18f2a9e", x"94964765ccf35f2a", x"fce2959e2500fcc3", x"ffec92eddf3dfb3c", x"451bbe2c76402007", x"8636adfbfd51981d", x"326fd31b89eb3c70");
            when 22926901 => data <= (x"e54788115502d7ac", x"f23ed8e5a388dad0", x"fda685d0db6191a0", x"ecd1470122ff057a", x"2464c1287a6278d2", x"1b9cfb6c44361835", x"e478f46b464816ec", x"ed09c513e3e4ae75");
            when 15844941 => data <= (x"bcc1f5888051d0eb", x"cf242ddb49703f7c", x"9068f61c093c20da", x"fd53589e8dd0bba5", x"53e03d79e04571c1", x"b17868a3ca1e85ae", x"af484f63c707fa39", x"9f932f991271a7eb");
            when 3502339 => data <= (x"ef8afcbb1e012549", x"bb87e776bc7ec130", x"f5901bbb31b2570a", x"51c8919f1c464f6f", x"caeac00d20d29894", x"e654602159fb3b78", x"b35c5396afa08fc9", x"3a30a208d3da9249");
            when 1294964 => data <= (x"4ac8df85349101b3", x"45af97cc30463ada", x"6ffb3616cd6eaf22", x"34ea23e0b60f998b", x"5cbb035865fa81ed", x"180f1ef0e5ec9877", x"9b6308e5583db879", x"26ef6bd734882051");
            when 32983370 => data <= (x"bf18cb001350093b", x"4117d7e291133de8", x"290bf82bea9764df", x"10b58a5eebbd4094", x"8ea4c708defb318d", x"18fb2ff64e51ff54", x"7284085a3133abe2", x"a4eb2adbadf94f12");
            when 22750006 => data <= (x"ed8b1e4fd166e55b", x"344e5df9f918af95", x"2c4af2e890df10b3", x"87970665456dec3d", x"3a9de905d9a2c816", x"4b6db1fdb05042e5", x"71776dd4a43e6be0", x"d432f1e8b28182bb");
            when 20916831 => data <= (x"a3677a622dc8e7fe", x"e27359b6b1722d57", x"4838bd6f3d34d3a0", x"4847955ea36ef9ae", x"1113907fd02caf1a", x"40e21ba6ed7c88bd", x"2d505d0648ec24f7", x"0ccfde104db252f5");
            when 16071469 => data <= (x"9f188c5261b990ab", x"3376792a5fbdb644", x"28c26da785465c76", x"dc9da3ff24b7e34e", x"7df040777a4a0e72", x"9f93b4ab609e00f0", x"aaa4d94e1129d6b9", x"8b7db40961771a61");
            when 244630 => data <= (x"839bcba3c77e736a", x"74da40269f958542", x"c8d6b1c663f193e5", x"473c01c282d6c7d7", x"2079b72a9322e16f", x"1360d64eb81ede22", x"56b9640dfb21d2f1", x"db08b0767e44cea1");
            when 12955676 => data <= (x"6999b2b4a966ed9a", x"ad99767bf52503fb", x"dca55885af11b0af", x"ea13b64f1c338d85", x"12d7b0040fbe7a90", x"95fac8b04c6b4fa4", x"e85d6427a1203c90", x"c484c9fbe8b7f655");
            when 28495129 => data <= (x"e90964851d85bb94", x"92581361effa54e3", x"ea7982b528be6399", x"125e8ad2a47437a9", x"432a56c4f8993be5", x"714dc98fc82bb0dd", x"d9d761508d2e95d2", x"b8ca6ee23f483451");
            when 30678127 => data <= (x"febc84002f51dede", x"89ce1fea70129157", x"c3ec3eb60037d739", x"01089a9ff086820e", x"4f6d696630b3d7b2", x"cd368f438993d6c1", x"f7a2f2f8665ce961", x"03b3d0fda81d6152");
            when 30640540 => data <= (x"07d2f5bf56ed52e8", x"ac260143d176f9d1", x"bb3e50cb758b0380", x"b744468ee7dfa678", x"5e3f98dbadc545a9", x"24319416eb4db8d1", x"a7eb9d36b657a6c1", x"246ee1f07dd336ae");
            when 13313678 => data <= (x"a78b553be9b20dcf", x"95e128772bff6304", x"948022669efa2c1a", x"156d674cb9f0953d", x"4ccb1b5cd563bd0c", x"678007bb1d45b3fa", x"49026ffd457aa0b3", x"e3b4711597888f7a");
            when 187490 => data <= (x"1915c64f735a5ede", x"95f69ca15989b190", x"7df3f743a549a6f1", x"ca69da31c2d8b1c3", x"fa04d96cca899499", x"7bdf6132bc8e68f2", x"332f55f9a70035b0", x"20fc0577d9f472e7");
            when 28840701 => data <= (x"6e15ad2aeb9027a7", x"27edb0d86f2da00f", x"9d4cda3419a694b2", x"662a166e37fc536a", x"d5a16fcaa4752750", x"633cf80183ac1a06", x"3cffdf97f63338ae", x"ca38a416e151a544");
            when 20552744 => data <= (x"09f0549cff3d62d9", x"21102979332706d2", x"c2fdaacd69f926f6", x"5d2d880ede0c2cdf", x"0888ca11cb523000", x"4bf9df7e68151eea", x"a96fd157d718220a", x"16db3f7719570b1b");
            when 1386384 => data <= (x"ab40f424177e88b6", x"e6fd4232db528bb5", x"d7be916cd1ee4637", x"ac162bbd4879da27", x"b65b07ab59fb1c74", x"f588126d6961c39d", x"0cd5848642ad7477", x"5b60c8849a4c8ac6");
            when 5567242 => data <= (x"e29c9ec4bd583d1e", x"4285a2607ec33d31", x"1348038c30334531", x"14ac8dc9369be5f7", x"8a667f5f2c49464d", x"f1e081082254a139", x"8202b78c145c5c6c", x"32e944461425459e");
            when 5703971 => data <= (x"6721229041218583", x"866a217f012b0cf9", x"0bcc1f366f93eac8", x"fec2711a2632848e", x"af6c9d624730283f", x"e850d34a7ece4c4e", x"53d023927f2eece1", x"4a50d24fd514614a");
            when 3806973 => data <= (x"371973568d26063a", x"1291799849f1f729", x"70e3b8ac9b1c86ee", x"a53dedf2ffe679a8", x"3bb75073a8cb91da", x"0c456ff04ec2957d", x"8708ba28a9da0a3b", x"f9a4d49ec7534292");
            when 4510707 => data <= (x"770c559e4e2542ee", x"6966916960f89387", x"d8790b14db27fb19", x"78839038addb5a1c", x"b65a08b0525a5938", x"21deef9a3de84d66", x"0c8825bea1147cfb", x"7c0ea6e41c9d8aad");
            when 16299042 => data <= (x"6fbfadc4b988bfbd", x"8b50a5198a4846ae", x"240ed6a5a1324b26", x"6927868f42f2587d", x"29f941e854dcd342", x"1319a76b2e6e3259", x"b03098e3293ef736", x"c469865d74ee8c42");
            when 3526318 => data <= (x"a88457aec6ed48d1", x"254e6ed6d2c17918", x"aea9ea334a94717e", x"820fe55fed8798fc", x"2c2b6030895152a5", x"a4041a5dad823614", x"aa6dd8280488145f", x"5716a4366b882b8a");
            when 1381145 => data <= (x"109fad5e9463ab49", x"14b6e07ed2b81124", x"740cc7b809082a3f", x"68899fa49db6438b", x"543b0c9d81425a41", x"a20bbfd5010007f6", x"5c4ac20eb93dccc1", x"eb9aeaa201905ca4");
            when 1584185 => data <= (x"dd933be6c0dd881f", x"a1b39a7306fa3fa3", x"ad17aa06b97d3d1a", x"808e736b5eb520bb", x"5b938314270f98e7", x"b520fb3415cb58d1", x"9b757528d77b17ea", x"50c06a902fef9302");
            when 27294872 => data <= (x"b6d8ba8d901d219c", x"928a48f18c9f74d5", x"a769fafac1f72dc2", x"160378becf4e6c34", x"faf753976e70ef48", x"6e46fb3fef4007ce", x"20c8af493b9a1b20", x"2361aacb4889aedf");
            when 27662133 => data <= (x"af8af194a5c6bf27", x"2768ecd9f4295f17", x"5934844c288a2267", x"749d4bad136cb7f7", x"9549a2ac06ff7e89", x"16af18009ebdc651", x"247b0df64cb26e08", x"c35f81298c803d61");
            when 16592257 => data <= (x"f63329ddc16169c1", x"dd4ea8649db783f4", x"07c43137467b6544", x"a4b1dc1b021d6c1b", x"77a12995c676122a", x"d54177484493728e", x"21a2d7d893754d4f", x"a9c0ac00e7d26e70");
            when 4037399 => data <= (x"c65392bb81b6b4ff", x"5f0f24f101be4828", x"aa690edecd58f9ae", x"2bbb9dfd41f677ee", x"9150cf1d4d987ef3", x"ccafc77747098f11", x"03487aa6a72b3031", x"ab6d2e2133e88c6b");
            when 5265819 => data <= (x"601e8bea9be54cbc", x"783d7023896b3919", x"69cee6f31c4bb553", x"473ab3de4e4431ee", x"84566ef97e5da08a", x"3d2e9e1616d5e903", x"42ceb3abddb1d55c", x"79c2fa51941ab3f4");
            when 28089735 => data <= (x"a7d320ff3368f99d", x"c1d97120a4b5ce06", x"745ea1f31a833757", x"9731780250b6633c", x"34b779289306861d", x"180e1f71b146f5e4", x"ea9639165f7f183c", x"c8861cdd271f36d1");
            when 31299616 => data <= (x"6a52a815442e9163", x"2870fbc3580c078a", x"2c650389ccfa7839", x"0e70904f0b3ed780", x"21e3ef1bc7af6b40", x"442fcd2d084cabfb", x"6dae9274a198b9d6", x"9bd5f2180ab3036b");
            when 2262241 => data <= (x"7204e2d6f07b9976", x"bc8bedbb8eb013f3", x"1050a213a890f6db", x"e1fcb25c8bbee953", x"c8ca495e475b8258", x"cbf6028081afbb9d", x"3800b946dba37c88", x"dde420deb8f1eb2b");
            when 7662388 => data <= (x"1369ad37c2cc03d5", x"3d4d97f55942e294", x"42cd0805b69e042c", x"a6b599adc172747c", x"7b082629a3519771", x"d23c93f36a606658", x"7ad992212bbd0e7f", x"8806e131b3275f51");
            when 7242004 => data <= (x"8379d7959b2ade65", x"37d32e92d0929e4d", x"0af443e7e711d38d", x"a4b07a30eede299d", x"8f22a2d394f7dc4c", x"f33f224df08679ec", x"07e6e3d84c72f95b", x"65d3e5ca5f42f9a2");
            when 13284908 => data <= (x"9eae89e157543630", x"3dc3fce8c4764e81", x"20468ffafed7bf54", x"6f39158bdf6f50c3", x"aedb4019a768cc34", x"ddd191a70c921d90", x"146bdb946b3504ea", x"859ccaa5f689984a");
            when 18902700 => data <= (x"7ece597565deb6de", x"03e5524b39a491a4", x"4aad48ddf58dc11f", x"d36e7365ac9d695c", x"694d32537af8d052", x"740a90e9ea3a315c", x"34e251e1344cc59f", x"efd168d0fd2f0c4b");
            when 30591133 => data <= (x"d379ccdb0f3f57d2", x"246bddbd53dd0cb1", x"55653c66f5865ad8", x"2ba86fa24a48a931", x"e1c2f4be20bc5625", x"338cb91bac8103cb", x"110407f762561269", x"263922aaa3c33abd");
            when 8594177 => data <= (x"4f36aa02dad3a00c", x"42f35f0c4cf43ca5", x"31fe324a683dbf8d", x"3b3fd541adc9189d", x"4ed70feb76e11655", x"820c2e803453590c", x"b85e47673002fa5a", x"f777af9431292bd5");
            when 16856707 => data <= (x"d3356867a16182b0", x"b358bf2ba3079b61", x"e63278e41a22e681", x"d27c26a0075a4c7e", x"48645d5b72bd951f", x"a3092f430bcbd648", x"413fa1a84b205cdd", x"0041e32111b86385");
            when 4432394 => data <= (x"03801de388257040", x"843d5019a66665f2", x"4776492b8c96ea52", x"46f1f5d944480ae0", x"fc79782eb2194184", x"a28d12f893c578e7", x"ad692a88db592fb0", x"357441b3cf4d4035");
            when 11071043 => data <= (x"e6aa69d7f5520d49", x"c79b1389b60a62ea", x"c5c39302936ca5c1", x"b619532a7bc03403", x"97296c354393edff", x"161cfba12fe4e60a", x"5a226355d1b701dd", x"5d34fc27802d6776");
            when 24335000 => data <= (x"de31d396f92cb7ef", x"55da07132aa0b0c0", x"287fbb7a8f571113", x"201dd80694b277f1", x"9023ae80394dc2cb", x"ac10acfba461ff34", x"50a373e6eedcf345", x"b474ce094c3185e9");
            when 30047338 => data <= (x"0dc87bafd4763fde", x"3c586a9a8a6ff5d5", x"a8a1a80daa244573", x"7c91722cc2be2e07", x"1acc034efd0c370d", x"1ab94ecdc6010ca6", x"d6f150e575767c25", x"f6cedcbde1c4bd65");
            when 28669297 => data <= (x"d4866c9361eb12d0", x"e1ca41b156f6c449", x"bd1d657c154ac7eb", x"dbe3fda5d280b320", x"c297218dfae2e0bf", x"ac34d290d3e55e77", x"52a0ade15dd204df", x"7cab4e9e6c9f85bc");
            when 7883258 => data <= (x"d92f08adaf8c3946", x"41c54f39354db952", x"79e5f7765f491bd4", x"5175b2086de3927f", x"1a2cc098cc979075", x"573d003bc5aab62d", x"5d1c8a3ea6c3fdf1", x"14dcfb3fe53f78bb");
            when 21016419 => data <= (x"ee5abbbcfbc265fd", x"e39257d25016163c", x"8eb2785f0f26bc15", x"fcbe48af9d29964d", x"7d1216e97aecbd3f", x"6f83d54f730d856c", x"08d12b67d02baa47", x"bf4ba6bda8855e67");
            when 26888771 => data <= (x"8bf1782aa97163bd", x"c32892544ee3a050", x"d765114a75d805f7", x"4960f50cf5c498bf", x"796a2b37adc19818", x"ba6f3394139b4e9e", x"6b27eb6e2d97fd77", x"107b83795af65440");
            when 27937666 => data <= (x"e521fa7f494f2170", x"ba4df03193438b4b", x"7a5fe60f6aa04789", x"0c3c6a5708ad1e84", x"55b6e3bfb2963df6", x"5f2c4e9c2363fd1c", x"c11652ced891994a", x"99983966f3fe869f");
            when 30395571 => data <= (x"be57a1c4571fd07e", x"8df173fce94137bb", x"8216b192e3b46727", x"0f5f98a2ddd39844", x"71409ab2f3c8677b", x"f0c26d3c93d743ed", x"93bcb96126743e09", x"59117ce3a557ed06");
            when 15356448 => data <= (x"483ed590cf82363c", x"80ed100eed330e67", x"46fba40cf9a0617a", x"4f0557900955cfb5", x"7e418451507d9791", x"0a54e834a1705189", x"e14dd3de2e6aec34", x"7f631ae70dc7d37f");
            when 236334 => data <= (x"b2823d79d83fb37d", x"31e1455702bec29a", x"864349b8954e2a60", x"a101563671f6124b", x"cc800b873fee927a", x"054ba1a4e75828ab", x"19b76f5fd2596295", x"2b9a8b8359686a3c");
            when 31921858 => data <= (x"33c604a8c3191b35", x"4bdb474031cb7503", x"54c93be26aa2148a", x"4223dc23d8801276", x"e00d5e14dbe8e632", x"c21451250a8e2763", x"9117a3aee93b5cf9", x"ed9a4fdd53b45337");
            when 20242764 => data <= (x"21083394e5b98af1", x"4b59da0bfb90052a", x"3bfde8648fdaeccc", x"9850ad1820ab85ac", x"d93efc93d9564ae6", x"b38520013e522dd8", x"3e28adb86928b14c", x"40d489341d71d95c");
            when 26037710 => data <= (x"76a9c85a3f1c3cdc", x"50112b2b02901b82", x"ad4a4558ad99e30e", x"559ed0cf11af65cc", x"9d7abd8b19f4275a", x"f3b7974b19ad1a23", x"509f4b719b47a942", x"3a12d5d6fdc06507");
            when 22835870 => data <= (x"ad1b6600f1c4ee6b", x"ccff4f161e483fa5", x"21a8adb6f95b4913", x"95e4d843092d44b1", x"18bdb371067addfe", x"c91445588c65cc74", x"e9d653035eb770df", x"1d02473dce0a1a70");
            when 3630892 => data <= (x"ef06c7adbaba4fa9", x"855a6730e27a43c4", x"d5686e7089c2b3b5", x"0d56e90be85d7344", x"99364efdba5611ba", x"be2fe49e8882dd54", x"0c2cea0aa528ca59", x"8c660ea62d7062fa");
            when 29269601 => data <= (x"7ce8df4b5d9c53d8", x"d609779d7f801f2b", x"97d8295c0399e318", x"da3f821e36203234", x"d90c335324796d65", x"dd6be77a04def6b0", x"9cef5ae64cd47824", x"e200d7932e8987ce");
            when 14815463 => data <= (x"7a94eb24947a57ed", x"ecdc384a32ae1190", x"6e05d34b88b7de01", x"33d0fcd43e2700f1", x"692d7c908d1fc607", x"2cc108f850ef13fd", x"f40aecfce14cdf4d", x"509b651e42e0e196");
            when 2039893 => data <= (x"0931d281df14d367", x"5c6ca9daf9bf4a3a", x"e2634f5e94996fdd", x"18b93a4e469f3021", x"3dac9a9aa355e517", x"2ff3c8dcd9bf2154", x"cbc565b80d2d372d", x"e620edd4615a75ed");
            when 19331267 => data <= (x"2c9fdc46c532565e", x"6cbd4cddaa0342ca", x"550d3cca430b40a5", x"afb7972685cf3752", x"4cf9606b8ddce1d0", x"e26ae2e91690f9df", x"ab5f443cf1c1e8dd", x"cb89f5da5f17bc54");
            when 23186200 => data <= (x"76074da9835ee5bd", x"95b3973ef5c38f17", x"a873e593bfca01ef", x"8f59279e9ea9ffeb", x"5f9c27eb6f07d116", x"c758d4d366b0f769", x"05493a1dfa0261c8", x"06095f5f8cb0c3f1");
            when 6446882 => data <= (x"e14f3f73a41b8b23", x"7dc5abffdddcf9c9", x"4bd80dbddbf7a069", x"3f13a6c8765399f5", x"a693277831a40831", x"85770cb4bf4ac307", x"553940329bf48e68", x"aac98556779737d3");
            when 16716495 => data <= (x"10ab57ba3980ed35", x"bb5fac6a95020fdf", x"4afb19b834a78ed0", x"e9705195a24b8a01", x"b0c6ef1aae80dde5", x"e5890361530f40ee", x"77b2b2ed04627a3d", x"f9a156efdb69ceee");
            when 18688392 => data <= (x"35d00a21a17e9865", x"41b6afba0bb68b98", x"dc4b2b9b4221db23", x"a009434f19bcfc3f", x"c35210414ce3bc44", x"981c6262916b2fc7", x"a0a8abea0ed88972", x"c161ec0b0ea8e2c1");
            when 20474894 => data <= (x"6d881eb134299d76", x"db0f73112a6ec03e", x"481a6e3006f7d28e", x"2ef4d4fcb77c1f54", x"f19549f02ddab408", x"6872f975aeced1fa", x"53e8fb9aa103cdb6", x"df9b5597a61d9d8c");
            when 27449714 => data <= (x"73305cc1e521e66c", x"d254cd13de5dfaa2", x"fcaee9da0292fb33", x"4625586d5b4f702e", x"b6f1c1b06e3ed121", x"ad3f01f26f29569c", x"566912da04d38523", x"9cfbc4a4e81c121a");
            when 31344090 => data <= (x"545ef3b0c8f48a68", x"a8a3eff121f0e9a9", x"c18f753936fecf21", x"1306e8c598637810", x"3132061ccf4a52b1", x"da5001f30431ac99", x"e5a28512deb6b548", x"5196a1fcd0c5c2ec");
            when 33140842 => data <= (x"8bcfe9685fd2b37c", x"ecc10a61696579c5", x"965ce9d33420005f", x"85dc8faf422ca3d1", x"18ebf3e5a1a71291", x"0a072b443e23caea", x"c77957a4f95be0bc", x"26746194d089ff9b");
            when 25108124 => data <= (x"41ec2f95b34feccf", x"6e4645e3c8702853", x"cead5cfc36241de4", x"c614236ab7a32f26", x"500cba9c4e2af6a8", x"1586c0e4fdad877b", x"139b809e2078265c", x"ae3ed5b7ba916ae3");
            when 7364704 => data <= (x"842bbaa76c579104", x"993f77c679ec2cf8", x"97fdbf414ffd3ce3", x"3480737cc80a58b4", x"01c9ae643eb04024", x"7589db71fa373323", x"7297f42064b0a448", x"e409ae58652f0ac9");
            when 17441636 => data <= (x"536f2359893b39f5", x"b151374fe4ed5f02", x"86eb74022e2e34b7", x"3f7393a026dcfe6e", x"011147569f7c9b46", x"b2bab78d2b9e4430", x"6456566b714e23f3", x"375d3348686333a8");
            when 14222822 => data <= (x"f3cfa019c51bb5bc", x"4d71b0612d2fc757", x"658d709d795fa76f", x"840f397a37dbbf35", x"0b5aeb29fb42f1e6", x"d7f8581efd52a20c", x"af10bbf96d25a2f7", x"8373829e8ccc4e12");
            when 25734202 => data <= (x"6f5e9555377b9459", x"e05c5bb29a0bd93b", x"d354c260f542dfef", x"02695be8ef35e702", x"ed60e365fb220152", x"92eda78e9c27ad61", x"df31e379588227b4", x"f97242024567dd13");
            when 32598092 => data <= (x"f17fb911d150d010", x"414abf511af843e8", x"b911e7dd393e3b45", x"af2974c335acd9f8", x"72d9c224b3c39e4a", x"7f56d53421cec90e", x"038a560ac8425aac", x"2653b726f328a5ed");
            when 2689242 => data <= (x"97c44ac5d4e7fe1c", x"095e6b90c4c4870d", x"9b21490a79c5a1e9", x"bc13eb7c55f2c266", x"7dc60f0ed98cb9f9", x"c0232859185bde0e", x"63842adb4d48f1f1", x"307205c64f62a170");
            when 8472232 => data <= (x"789358f782ec051c", x"dc6c62b58e96f270", x"e4fd2c1f91f449e1", x"cb03b391b9c513ac", x"3e991e140b5aa25b", x"8ba390e0bf495738", x"b99658e2302360e0", x"9f1249fedeeea743");
            when 26873683 => data <= (x"a73ad0bd2882b2d7", x"523290608d9b527d", x"8365be1fabe39646", x"2f6e53088d95490b", x"eafa3aed1e163510", x"a573f9bb137a7e91", x"a6065ac84a74ab17", x"4c9606dd4db1f250");
            when 1447174 => data <= (x"3f976e53271b8ea6", x"d45e4c2bcdc057ac", x"d1f21b48db4c1a22", x"a4cdfa623741520c", x"6f92819dc68d611f", x"9257349a618dd9c0", x"07ed6fe1b1514379", x"0c37aa4d88603fca");
            when 17692099 => data <= (x"884369bf7a1f31a7", x"6048499c213d456a", x"5ca64ae896f17518", x"0265806df8df3463", x"6915055bedf7e7c1", x"96969909c163fa0e", x"70f8c17e0df301f9", x"9fe57671b46d5f2d");
            when 5118509 => data <= (x"487cd7dbc320d05c", x"674fbc72dd1c97b8", x"5f9e3c55cd9c7fff", x"cf8411803116fae5", x"63b92ece3ed936e1", x"ad15140bd5246cbc", x"89b68241a4d83374", x"ae368066e234de96");
            when 30786974 => data <= (x"cda01125f641f145", x"0c073aadb00497fa", x"0c318ee7703130d6", x"32b5f92917275133", x"6df6f825309ac04e", x"d00e1652afa64e53", x"2c6a331b3fbb949e", x"4465f890dcf6b6ca");
            when 2676465 => data <= (x"e2bcac9f78ef43d9", x"1e96d9e91ff3de80", x"7626598db476d7f0", x"aaa31a497d95a155", x"6d7071de102e6347", x"70f892ef0ebf91ba", x"bde25f58723d43c1", x"f8f6bf2733f83f02");
            when 13750826 => data <= (x"5be1e79fc6ed401f", x"6256ecefb03b819b", x"4d7cea8a4525a89a", x"0088fd93b111f342", x"f9e78a0b8e11c3ee", x"8d221596b2a4594b", x"c703354db916b6fc", x"f258b07bb7ffb9de");
            when 25527732 => data <= (x"b8de1d2814c89258", x"8cf692e3283765c8", x"7bea10e1ffc37902", x"90240011cc81575a", x"3655a2b3e94a442c", x"13d628ad3d4c1bae", x"5148c9abce612459", x"5826d8479273d091");
            when 9113935 => data <= (x"a9519bd932d2e320", x"31ab972cb7c9e393", x"aded5d4bdb47a36e", x"bb89859487dfbfb5", x"dec8733d61cb4eca", x"963fe5d710977b6e", x"90376083a524f022", x"611a05996a8a6a5c");
            when 15051537 => data <= (x"aef7a9bb8d5246a8", x"8591d7d8057066e2", x"e20e5cb5863cdac8", x"7123bd67f0055816", x"d921ab4623987353", x"ff325be4e26eec47", x"0a79dab26d11d037", x"dbc128d8d35a1f2b");
            when 16975712 => data <= (x"9f65a5ea2118b918", x"2a6dadc2e9f2f86f", x"ca0a65e9ec874333", x"8f70492fd6c536cc", x"85d1c45aa5348f07", x"c407b450e46a36f6", x"93d459f69bc1c54c", x"fc0350dc1395c093");
            when 16675157 => data <= (x"8d00613b04bc7ed0", x"d2f4316c98749715", x"577bfa47dff60653", x"3581d27581426c4d", x"42085e4ef65abc8d", x"548bf7d0f7bce6f6", x"9c8ba809e15799c7", x"538c10513d1fc211");
            when 656531 => data <= (x"7e977487ecfdab96", x"574811bef6677997", x"4a51ce17586479a9", x"26608b696c17072c", x"bd12dd0fa330436b", x"8fabb44af78e3678", x"dccc7ca2d7abc7ea", x"88eadd07993e7fb1");
            when 7544889 => data <= (x"df92f8cc508d867c", x"e6a3416fb7583373", x"12fe6b1730ab78dd", x"651be0317770e560", x"8880c90e59234d5a", x"1f36c3f5e8ea337a", x"d2c86207b9ff4600", x"f879f5181006e0e7");
            when 32663445 => data <= (x"b4726ea72e266a5d", x"d822657dd683b789", x"bb0608fb8dcb7588", x"3c1c14e5ba003b0a", x"a4aee9ffe618b585", x"198e0b795c13c320", x"d98c89892085260a", x"7477a0244f9cdd3e");
            when 33494530 => data <= (x"fe0165ec54ab4f77", x"a892e3efbc3be619", x"e17c787581b3c607", x"0f38ea3142665b4f", x"7618f0a0c41552bd", x"11e948fe2b08e2fd", x"b990c06e64690a19", x"e5f8396fa649d4d7");
            when 30521047 => data <= (x"75142595b2c6481c", x"44ada93f2af31746", x"af0a91d7d1f12fa4", x"c8b350e48393f34f", x"806644f8b47d7eaf", x"edcb9ac7a6a1d4a1", x"466eaf855cbaa482", x"12b12113fbcf08f8");
            when 979247 => data <= (x"b80f40e1e1cd65fc", x"6f9ea2662f6207e4", x"675583a899d1ae6b", x"8681bb8712526ac4", x"f3f2c3a06f847701", x"eeb55892f78031ec", x"be41d14406514aca", x"3c8a7174e41d9115");
            when 29218469 => data <= (x"d8c6c1dedae18422", x"1b562710443a2dc1", x"09fa843c40870fa3", x"78e5fdd9822c5f31", x"ff37c61f56a63156", x"30381053614e1c03", x"46ca13a30d70e164", x"e578659cd51e6a4d");
            when 8499834 => data <= (x"1b98fd4827ce329b", x"7d6d72069e74572e", x"34079609d8bf54ab", x"aaffc63cd1aa5cc1", x"16edac325b2eebe1", x"60ca84b0b23ed87d", x"5b71133fe3a8bbf4", x"25ef6f3598479eec");
            when 10727277 => data <= (x"f074e9da5a12face", x"c6dced5e0666d42c", x"962779b75b297e56", x"7648b7a120d1cf61", x"becae6d6121cc3da", x"ab87705b97d51b17", x"562b53a78d5a0c9c", x"da2f2d96b89bfa08");
            when 10656410 => data <= (x"dbc189b1afbad65b", x"a62e1167a44aa144", x"d30d2ee8a3786e03", x"46ba09e99b8ca873", x"37cad2241a029da1", x"d1bc0e0a8c072dc6", x"fbd15427eaa9c307", x"ecc0ee0347ed0bb6");
            when 11116001 => data <= (x"677ecde573ada427", x"828d15ac4b2adbde", x"8625c95fb3ed1082", x"51d43e0b0a1bbcc5", x"e3992008d010ee3d", x"5ec0bd2e1ea4040c", x"d2c303b1ce44997a", x"30a2020594c5cc96");
            when 18650683 => data <= (x"ef0773a5cc0e3f4c", x"93e114b84edbe71e", x"b336538f47882b66", x"acfb63e4dc162edb", x"f78346373ff0f2f0", x"5755b426d13eb8f8", x"3df4d788f98ca840", x"2346557e6eda0d08");
            when 21068584 => data <= (x"39015c009fdcaf5f", x"7913180ef390fcb9", x"b3f6eafb839ddcc3", x"a2dbd89ed49d6879", x"9d04601a6c789927", x"c5901b815f52100e", x"96bf74c2ca2d3ee5", x"1c4cbe59ab817f99");
            when 25901003 => data <= (x"9219ce4eaadf1c47", x"d68ea769b1f68b9a", x"51b8649ee24fe868", x"9adca84e41f551c0", x"98016c60cfba0e42", x"0a1400e2f894aa7b", x"b0bcf51d3fbf5995", x"2907aebab5dbe20c");
            when 12448022 => data <= (x"3217b561fab53f0c", x"ccd6bab3c791b9f9", x"ef7291e7675a0408", x"3fcb08249e530906", x"fd3f9701b2f943b8", x"70668668b627a57a", x"0511f8d7b84d5d9b", x"f54a2f144f6f6496");
            when 33325143 => data <= (x"4152a90145a1edfc", x"95deec2802462002", x"e72f661cbbe8bf59", x"6586e301ca0699cb", x"173bbeeccbee76a5", x"d3b5fade52e4899f", x"418810f69662899e", x"7f02790dbce018c8");
            when 28082368 => data <= (x"35afe9af19f59163", x"89ee355bf52b9c75", x"4eb21956765b6f21", x"086472091208b6d3", x"70a84fb9c6c93883", x"2c7c7d1be83bcf00", x"8bf0023f16f942de", x"c53f0dcf4eb91e0f");
            when 9929288 => data <= (x"4c7e7a079b368406", x"4db7a4ea0de0153c", x"733f8d4888d3e100", x"2d5e74199c5b6672", x"16d5f05dfd4691db", x"7475f95a064d82ce", x"3dd1141eace991aa", x"3b2b69e3362037b2");
            when 1447191 => data <= (x"ea513ced6abf2584", x"03043291104fdddb", x"6578f1f1a9b8c544", x"16400c0dcfd3bc4b", x"052382b2a3b30388", x"016cd76c4a464555", x"6854305e028735b7", x"09dcc0126e7d9627");
            when 22544131 => data <= (x"a242f2ceb37c44a0", x"80c54004681033d6", x"b3894def591398c8", x"c97cae0c28b644ac", x"96147b8658bc97a1", x"05346719678c2475", x"ca7cb87611eab483", x"b38a2b3413d49dc8");
            when 27082473 => data <= (x"297b7789e116493c", x"0e305022b91f3f7f", x"ad8d6f92a983809a", x"34c62cab316940e6", x"a1074a024cd16e3c", x"09d7f7048b97e74f", x"0d21ee0db10a6fdb", x"f16202d6c0aeea99");
            when 24310713 => data <= (x"1831f792677643de", x"b016917490d13939", x"19296f92623550fd", x"31ba3c95e8a36a69", x"cc3d911e0439cbd6", x"0fb826b15e2d3672", x"dbfc1ee8904fb386", x"e1eae32244ff7167");
            when 18776653 => data <= (x"65652b625790cd60", x"6fbb87d75cc130e2", x"1a8805da2bae6d63", x"3b3446e94e57b522", x"a9c859588b0e8b8b", x"0493e82a3dcdaaf8", x"26a14905305c8fb1", x"272e1d04449bde19");
            when 20334459 => data <= (x"0d3ce4e052c96d85", x"cfc73799df704ff8", x"aee2f407195d5c46", x"4e15d89a60c7f930", x"c387ca9554a46bfd", x"fc28a2e6f63fb415", x"8c4a67f239dee9ac", x"7bdb1aa776e5c092");
            when 1298638 => data <= (x"2d2b4a081bf09d13", x"ea46ea6c4b92648d", x"e128a1dbbb992cd4", x"4cd9134bc933b0c0", x"969ab000a033b95b", x"00b409a3b55672c7", x"71af5929fd15164d", x"1e6d6b0b1b268dbf");
            when 15691114 => data <= (x"534027944aa7523e", x"02bc6cb81702445c", x"b0da4172a2571353", x"5c50fc793ff1d964", x"61856badb99a780f", x"3d4a68f2e252a4a4", x"aac7108dc445e2da", x"28fcc1079d813acc");
            when 28175206 => data <= (x"50efafeaa2480a82", x"e8b3945e64b87e8b", x"cccb4302a0e96806", x"8657e9b630deafe3", x"98806a1da08dcde2", x"7b4a7b058a63f921", x"8a15a685db6e0178", x"34350b1a906b6152");
            when 16719170 => data <= (x"51d052d0fadf37b9", x"e10ae383b5727f64", x"eb57c7a3552d7cea", x"49015574a1afd2d8", x"332cb947705b0ef2", x"e0067fd46d7934de", x"0abffe87538f28b5", x"b42f49ba74d53380");
            when 5603710 => data <= (x"3ce4c1be56172ac1", x"ca8b19811c412640", x"f4fc9c08c0d31160", x"b43ff7b0be79ef41", x"371d314a05ed6f16", x"415b635df88cf4db", x"b7669dcd2e4a5383", x"44d41c11e5c403bf");
            when 29842962 => data <= (x"4d3710f49ae64d64", x"68741cd92856bf54", x"e8dfd49b863474f8", x"331a5509ed4f58eb", x"d89c70e1df302dbe", x"0199fb6dc48a3df8", x"4bca5713b0a03c31", x"2bb234c75ac381e3");
            when 26075856 => data <= (x"691ac5537b952a1c", x"37a74a330c422309", x"d4a068012ff55588", x"58ae117aeed0e837", x"fa64117f36ee8869", x"78c1609538f24dbd", x"c49a8b96d554547c", x"7a6000bde2f319a5");
            when 26621712 => data <= (x"fa69bab742fca547", x"a2f1e065970a76a7", x"221e596fb6ba8f97", x"ceca57c705bdddf0", x"27236a229ff60769", x"275c09f8b8821859", x"6c48136f28058acb", x"4610fe3f42178e62");
            when 28650073 => data <= (x"6c0cc99bbd7c2cb6", x"6d48eabce717b72f", x"622fb7646c2ae3a0", x"9f13c336a8423479", x"84aa4a907b6147cf", x"678283756943cf00", x"30dc07f3fcea30b3", x"229afa714daf5ad3");
            when 32426322 => data <= (x"8392bac404784456", x"fd9bc4181b4e127e", x"b14eea276070d8a9", x"70a62e8bb4c9c623", x"e9313c57199569ff", x"6e9595c8cf14a427", x"4c3cb62db29ccd67", x"a9b648e0c901d674");
            when 20133687 => data <= (x"90c8f589afc9fd52", x"fad925f6e5e95cb1", x"5905c95261506323", x"0f33550b7bd25871", x"b435c3ea357744a3", x"c4e03e85a11351fb", x"01d97ccd16ce1049", x"4cf61522d8bf3cf9");
            when 11520496 => data <= (x"791339c5a293cea9", x"29461645caa926b2", x"d62a98024bd19a40", x"dc1e4e858da2c308", x"402a2737e465cdc8", x"7e48d3a6c2b7405d", x"8be843edfb06c0bf", x"abc83918f599cb39");
            when 691364 => data <= (x"af0e022cda7bd9a6", x"9b9c2db93243d879", x"43f9fe87704cac94", x"bfdce812632d34c8", x"d284dc94f4a5c923", x"c2acea1cfaa1cf88", x"a5d8084367eea90e", x"5c251ce3ef3f19c3");
            when 2702690 => data <= (x"2de5d84b84f252e3", x"c54641f3e2a2c45f", x"2bbd242c9d3766fc", x"b605b6a1ba89d65d", x"f01014a7c06b8f93", x"ac03218adb85aa2e", x"86ccef2d17ded656", x"5becfb6954b0fd3e");
            when 22843563 => data <= (x"d641e914e2c011c1", x"427d7940e41f2c6c", x"9e3771a9540bc070", x"7875e00e378febf6", x"6f9eac03d3771d54", x"eaa0a0af8fb9c48c", x"51fbd4f01bad08f1", x"d969d3a1fc0667f3");
            when 23839359 => data <= (x"ee53b048c4f3e740", x"7db38d09842ad8ef", x"50ef6ae888d67163", x"d0a777aafd96d7a3", x"88cfc175b3e0e8a6", x"7bb373a1831c1c05", x"9ac6e09b85a6027c", x"19ef3853c05f0fc5");
            when 32582201 => data <= (x"d1ed4ea4678e7999", x"5aee78525b075e62", x"437e89120e8b3d89", x"3f67e39642583d60", x"f901e817e1ac0d91", x"c2031b1aecfe015c", x"79c2b2888342ee69", x"86ddc5c69768c2a1");
            when 22568279 => data <= (x"854385df880eecaa", x"e7f28a1a5d936da2", x"d0a379030dc8ab19", x"3d0afc68cea02073", x"7a1db11aae1ffc36", x"53a2f7b1da17fdc4", x"f3ca88487ef2667d", x"1b7d5b2650b7811b");
            when 2370836 => data <= (x"4df24c098e1eccf8", x"412c0004ced81fe1", x"40cf6a46fe7bd3bb", x"a3507e5b54d9fee6", x"1795d506263c980b", x"a58937060c7edc2f", x"7a1c80bf530b7e92", x"982220fe4e2b267f");
            when 30017883 => data <= (x"9c99fa36d60c4aaa", x"f33c306ead8e5d92", x"33d5a41f24cf48f6", x"cc0e2ebaed5b17a1", x"475451e9ff54b1f1", x"f77cfd38761ddb69", x"7aa7d4984e0d50a2", x"bdb5fad78bd92672");
            when 19410520 => data <= (x"78d8b43bd5e39785", x"c7ba30ffc861b83d", x"374a5fd5a1ecd631", x"734a1e483085e16a", x"7299ed5d080d6b32", x"b799fe7756dc90a6", x"d6256748f73e68e8", x"8f3f37121b85b587");
            when 29141918 => data <= (x"73761a4892aa1389", x"786354cf76063fc3", x"5fa98d38b4dd93be", x"4c5768147639e8c4", x"4ee9c804a7eb32ee", x"3e2b9dbc7cdfdc61", x"229337450937bcf0", x"f2d7db4840441d49");
            when 13481396 => data <= (x"b20a8cf338c39ddc", x"ab760740de36cb9c", x"8f795a0fd8f12341", x"c4c81c62cfcb86c6", x"a88b6b1003a6ed1e", x"24fcd004b6ee9f1a", x"cd1b124a32b5c536", x"a3ca9e231c935991");
            when 10457121 => data <= (x"ff2d484cabb648cb", x"b57769d0a32f0858", x"6bb755c6b470f920", x"2a3c7ba0c60fc27c", x"37bf9290e4a9e156", x"3c5990238fe14007", x"32dd74f7fb87cd8f", x"66fd8e6624b129e8");
            when 11057585 => data <= (x"90b5d083b0b535c1", x"202ee731a96710bf", x"d15ec14603081c70", x"6582d8480dfb03f3", x"0f137463dc235955", x"298f32ea486d3ea2", x"236d75857dd6498c", x"53fd6fc324a43d45");
            when 31567656 => data <= (x"453b1d9879208182", x"0c3567f0ce34b90d", x"af45e06916b6cf11", x"2efa90d7345b4e33", x"e65baedd5cd97bd8", x"0c7812ba05d388fd", x"8dcf98d3bc7625a3", x"e9b80fd23d0a24e8");
            when 21154525 => data <= (x"09eb4f8262bd5e27", x"7f5af99983a89a44", x"128494982391219f", x"c0d595cd24b69362", x"799757fa14984619", x"d8338a252107b298", x"bbcb7738c02a7425", x"466e8ee67688d0d1");
            when 33153759 => data <= (x"603b835cafda3826", x"5bfcc1e9e575f78a", x"b90c3ad1348c1d21", x"32b9db6b37928e7b", x"5581702a78be7d96", x"fcda9f27e83015d6", x"246ff6f283d2531c", x"bf8a164da1f9a9c2");
            when 5992978 => data <= (x"a2b8c958f8800fd0", x"a662053a5b41ee1e", x"62bb2bf01c6ec9e5", x"bbcf677bea2d4a3e", x"afd2d9901f10f5af", x"27af85f92bc3eb68", x"fd737caf02822665", x"257f739981cfd47c");
            when 17861744 => data <= (x"e69b7bc886fe8777", x"69bc44564ed6fc1c", x"d3a65c5c2bbcf7da", x"6aa9847313aa7041", x"734a2fec6233aba6", x"6a7a1a6fd255dc7f", x"8f1aef6bb8f90239", x"d47e010dfff46674");
            when 29580997 => data <= (x"e68621c0a3781b2b", x"f57f66a8bae1844d", x"eb8783c5ff4d7304", x"81f09b9e1e72e13a", x"9fd488ea3225fe45", x"1bfdc21e1e41553f", x"8a8fad98df9afd55", x"a4281377a89874ce");
            when 20310103 => data <= (x"ad516fb14d4a0e64", x"608080413aebb9c8", x"4687a63c10ead9e0", x"c18b0b2a9faffe4c", x"bd97542f1346f890", x"14eceeba56f8a0f1", x"311a81b49b5efb37", x"2645ab084b466330");
            when 19784090 => data <= (x"27077d3c3fc8ea19", x"25f852e5c6dcafba", x"72d9cc9527c732bf", x"f4f0ef4fad512367", x"a0fa47afe10972d2", x"fb934ae2dc71da33", x"ee743558869105c8", x"418dc31146de1854");
            when 6678819 => data <= (x"52f1642dac2feb6f", x"0a3d0fd952eee67b", x"b546d4eba1e7a0d9", x"c1540ecf35175ac4", x"cbf15af08bff4943", x"f634173ee3b3fac2", x"96811b5576a3b89f", x"d2e9252956c1fde6");
            when 6564300 => data <= (x"1c939c6bf90b3ee4", x"93ae6bfd47968cc8", x"55fb87df6129681b", x"635f13fcfcb151aa", x"68901853e9e6797c", x"4ee16a160a9bfd65", x"7e30c54129ebe72a", x"433136160f940615");
            when 23558199 => data <= (x"1073f6089dd25cb6", x"76a30b35a184a735", x"f3cbb97d0ed5bdf0", x"6c4500ebe1d2481f", x"6607a718925008c2", x"f88f121d1810d25d", x"9ba6000d484e0537", x"b766ba56b49a07ce");
            when 29081933 => data <= (x"bc0d4eb7e7585a64", x"27792fbea8332250", x"92cbdf7bd904c097", x"c068a83e1ff84902", x"c89212c072e6c980", x"6384c6639615fa6c", x"b79f999da2a3fe99", x"fa8e5273f0e33835");
            when 26612778 => data <= (x"deb6ab04bdf7b197", x"9d604532f6087777", x"0d530e0040655495", x"3885802fedc52465", x"90e1ae6bb5c0347d", x"815a827716679170", x"3c3eec180bd771da", x"9c1b7447b30f01f2");
            when 28531987 => data <= (x"429b678007cf786a", x"7a0788a8d1179361", x"f5da4fd4f36409e3", x"9173add0f51ccbe3", x"eca3b924a3b18061", x"1bfe295e4c43a522", x"db3b8283c1041456", x"beef8f25e03ecc61");
            when 28077503 => data <= (x"b8ddf475fe0a9612", x"aa32608a63b73b38", x"c5f0d4fc8160f405", x"cd460fd7a33a54c2", x"e3818b4d9c8528c1", x"bc683d8db1348f25", x"a9c9ce84ed8d490c", x"b21ff7c1f0bc0883");
            when 14736026 => data <= (x"a7ac1f88a4951624", x"9639f4bf343224fa", x"fe994089b3f2bd51", x"7777b0129120e9ed", x"1f1acb3c13f65d01", x"17567afe73457c89", x"49fbefaa9b1f75f5", x"a28362ea35b00766");
            when 6148975 => data <= (x"987076571563d71a", x"7d66d957c6762897", x"460979e0f9da0dfa", x"b16933793c890f61", x"a6da26a03bd22b4f", x"733d7224c0178e8f", x"36b5de3607ee5a89", x"cd7118d5f3aa5b94");
            when 8041334 => data <= (x"1f1e39221eed7ec3", x"6af27e6db8ddae04", x"2798939973cf9b84", x"18475b8e482efbcd", x"0efbeb1ded456ff3", x"d3cde4c847794685", x"6c0b80f287aa8fef", x"935b47f296ac6075");
            when 12995769 => data <= (x"524df96833477222", x"1ba47f7052d39f53", x"c9b65694054d4462", x"468787face35556e", x"7f3688a6372310c2", x"7a23000c32d48de2", x"6715009add5997ed", x"b3b79ab32d0ff139");
            when 7014331 => data <= (x"f6e1cc3ff54e65f4", x"cddbea6f28a21ba4", x"dd25585ad50664c7", x"6f9c44f1c30b41c9", x"969807c98d8671dd", x"4c6ca957d735ac16", x"2e93addfacbc1d44", x"9f075cf1951dc7d3");
            when 16641096 => data <= (x"7e87b018a44e5512", x"b24f0b16f3a8f7be", x"45dcac79d55c8a7a", x"158b37210bac93c0", x"5016757790de9734", x"532c1497a624f578", x"1fe98a8492a4ecdc", x"aacaed280259396c");
            when 876295 => data <= (x"5a5f5d35f827cf00", x"f6abd4d15a957cda", x"af2292b5de32a685", x"05b87e2f36183d1e", x"6c7ed7d66c0ea12e", x"2e2a9c2496069470", x"706aa0d3cab8349b", x"5c02f4b2f0dba7d6");
            when 20493753 => data <= (x"87a9f0fe3f0292e3", x"ee131f3358b6a08d", x"c49b9fe351fccb46", x"f6d8f79f08e68758", x"d69d33c6c4cf8cc3", x"5ce7e8c3d3a8cea3", x"4ec641ec248ab045", x"8c041d373571471c");
            when 26879430 => data <= (x"d7793ecdc37ea200", x"896f745bde249bde", x"81f0fba4ec55777e", x"83618360819cc559", x"e125b5a6455389bf", x"c80ffb40d2f90648", x"e727f7e8a671ad40", x"5b97d7ae6510bc5b");
            when 16244874 => data <= (x"f685597a04f5c938", x"51344d35dec2c5da", x"070d10b03fc1dca1", x"2bdfdde47477d754", x"dc7809678c9378b6", x"f195a91257b8c81b", x"88f1dd9e92097eff", x"6ef96860d231355f");
            when 5833802 => data <= (x"16424dde6b133fc6", x"3b9f0b69de155218", x"fea02c0b98765d30", x"3d67f9070b584a6c", x"6fce2956f67b51ae", x"af5286cb4889f729", x"db5f21d72cc54045", x"a55b091caef054f7");
            when 24604816 => data <= (x"3fd68f80435de500", x"ef23fa809b2d7576", x"120a8446f70f0f2b", x"a6cf0fc348a1a6a0", x"afd09cdc2e5dac10", x"7613132f23574043", x"85d00efda20376d9", x"d3112257059bb884");
            when 720243 => data <= (x"111b1061686bbb07", x"57a36d064eb3528a", x"397e3e30789a9ca8", x"89f4b732572c989f", x"801c2ddcd623346f", x"46903b0c6df3c424", x"ac261639ec4a0b35", x"8d28ecc53d86f968");
            when 29605525 => data <= (x"0e9cf37ca20cd00b", x"8f1f43a572d6e9a9", x"0545c1b408694484", x"9fca0840946cced9", x"fb692c07b6f455dd", x"bfb33128ec5fee8e", x"2e67a3a3f42e9ea5", x"80a6aa466c278ece");
            when 13891063 => data <= (x"b29d148e96153795", x"46ee90e00c0487aa", x"cdf4711c2d19ebbf", x"c1aa8d60660ec3d4", x"486c6b46c5b4e8e6", x"3fdf5a7c4d3e8d90", x"7e9de2f157c37a29", x"9d33697afb28bd9d");
            when 25221922 => data <= (x"a3800e7b97e3bca9", x"6b74287ca761ad3a", x"d7dfd43b7c2eebd3", x"52ca95a13e69e1bb", x"9c19b6a909938857", x"518a0c555725765e", x"35df5ac4616cbc5e", x"e5df0d1b5ef02e7c");
            when 12747314 => data <= (x"b0621fe6c9882b2e", x"96cb5015a618c24f", x"5dfaf10be0e305ae", x"1f2e5d210a14fc73", x"3ba1e0fd1ae6b8df", x"aec28153119b7f9e", x"7e8d40811467fa7b", x"158b598488e58ad2");
            when 15864211 => data <= (x"8d7ed118be65da42", x"c16727b3c5662735", x"5481536b3a12eeaa", x"7fe3e21c96737ece", x"caaad0502091f7d9", x"b501457bca4008af", x"587ebf7c78c598dd", x"b555ea568994485b");
            when 3295024 => data <= (x"b72b7436ca565ee0", x"06f8bedde94048a7", x"52691dd51298f8db", x"4f7731351a808ec8", x"d297bbbf9ef12902", x"cb22bccb042c5fc5", x"0e82fc9f90833922", x"5cf5ce988bad3737");
            when 14631554 => data <= (x"6e18e09765300a1c", x"fad5ddce26f95721", x"47a7d0f440070f96", x"ad9f0524b1ffe8da", x"92a8dcd61986878c", x"381401419e2a38e8", x"65b5ec778663f4bf", x"88477733dad79f87");
            when 15722851 => data <= (x"ccc57460f16a8054", x"8a3fc95b27773e0c", x"ccb5482f586bc9f6", x"d0291228bbd0223e", x"265795c660e31764", x"38e8fba20cb37ae5", x"eee850b66d302484", x"514a435d2cc3ed01");
            when 14980366 => data <= (x"9d1690babf79d6eb", x"7e7c6da61c7fe80f", x"4e1ade1460cca4c2", x"a0f82eec12d450f7", x"2f9c26be9ae75adf", x"5e7c36ceb1c3893c", x"95e4b38b585e5c38", x"7e97b99c7ed80cb7");
            when 30963758 => data <= (x"47b01a0afc2fe4f9", x"6af3f72fce241cbe", x"3fe2bd51f3f80735", x"8038a5a807efb830", x"112217f9ce7c66d3", x"e2345333ffb24f8d", x"ef360c91cded2f1b", x"c7267eea46d70dee");
            when 9954314 => data <= (x"64579de89ef4de11", x"1d581424c563fa2c", x"ec37223e0d25247f", x"ce9d0a8dde9eb7bd", x"8f0a53a75c4eb0f2", x"4f0f0ae47b41b966", x"2ea795e590b9d6da", x"4474386565fe2bea");
            when 11310311 => data <= (x"e2e19e7452f66ffa", x"201f256981d336d0", x"e2093e31d5426e95", x"7e000d911367294c", x"35943d103ed2104f", x"6b975ff45c6a237a", x"0230c41be6583ae8", x"99cf5527ac721d99");
            when 29385563 => data <= (x"80191e695c2c078d", x"419f3606b620da30", x"86d0731a3772a5f4", x"038469965ae23577", x"75a4451b56c859d4", x"3209d3038482a341", x"4f19b5ef7d58cdfa", x"14baa02a731b0bb6");
            when 23477495 => data <= (x"7fe0631e8faaa7fb", x"613664f109d9afc9", x"70892f076d455c9f", x"4c077ee0dd8506fc", x"71a9f2c8c9100a60", x"a760a8e28c171a0a", x"f86879a3e91aca18", x"dea91d75594d9c36");
            when 20406858 => data <= (x"c96d259115b785fc", x"393bbaa41cef861b", x"ab934b8a4c6adc89", x"bbebd67b57bfd1de", x"bdb4cb3a729ca390", x"df1e5c99d603a965", x"9ec48017042c238c", x"d6ec09a68371bf94");
            when 28165774 => data <= (x"eb34397a8077ab18", x"8b5e931fc474cb6f", x"671282a8b1e1848a", x"9023317fdc5ed5cd", x"cfe3064138dfce99", x"b83276ad23e95968", x"676cd5ae0a5b4b1a", x"78480945abaa4fe4");
            when 19966912 => data <= (x"a516472ff06bb6e9", x"8555ffa792409261", x"8db94693e9329def", x"cd72fc2e3547f078", x"3881af2c159a59f8", x"114fc859b41f37ae", x"a6ea12651592dbfe", x"7ae6e481c90dc311");
            when 39464 => data <= (x"e6696cb8b3e15bec", x"3301a6e25f477930", x"2ef02a61a82bd01e", x"e49c196d38e37f35", x"6b0c19a8c22c5699", x"360b317afdf8e687", x"5a27e42630923ae3", x"c67f7e9cfd361a57");
            when 10734022 => data <= (x"63a463e16f5c557b", x"d5afa177613d3190", x"d4d80ce1d37512e9", x"3c758c3a0872bfc0", x"01f81ffa60dd5d49", x"76c1932018bf8f5b", x"a595ffe98ec35b8c", x"e6ebf1aec46fa7ed");
            when 7275483 => data <= (x"2dabc4aee48db07d", x"19d67b7aae9dc8ce", x"54deb1e615161dfd", x"da52812f6ee0b02d", x"b147157a28e9d9ad", x"f2965808792f87f5", x"0c12197a228c8a16", x"6373820815f89757");
            when 29475997 => data <= (x"b2bb210e7bd70a02", x"80bf17fdb82fac0f", x"2db4cdbbb9e1f23d", x"a6e82c556823f4e3", x"8ebb330c11d58a90", x"6ab21e719a74dd9d", x"3522568a7db94aa1", x"dda943d00bb78720");
            when 13191975 => data <= (x"663230bbd14ab0e9", x"53a5e39a88c0c843", x"e2f535a89759ba76", x"ed86c4d3f10f46be", x"2a577b50943adc4d", x"9ce308a05267dd08", x"2f6db7b4c8ed5336", x"a7cb389ba7c9de2a");
            when 12459128 => data <= (x"7e34767b363a5af1", x"c8dc181e0d80f199", x"fd0e75388b4c658e", x"8851456099964b79", x"0551d3e99968861e", x"376a32bbfaf06a09", x"f5f3b32bac4cc794", x"3fa7156e9c393659");
            when 12520963 => data <= (x"29573cc964f6299f", x"42992219902622bb", x"7ff04b17dc696f23", x"d531a04285a57bfe", x"e9b6831b65b3ea4e", x"e2e33565917474b7", x"d9adc7ba6ede48c8", x"0c109c84d241e5ec");
            when 21532341 => data <= (x"e5868a7e02f891e7", x"6437f8295cdb9d1f", x"0139c48769aa9ad7", x"5d71331f74fd5c07", x"17b451e038879218", x"6b874307ef88ddd2", x"4dedaed065e52bdd", x"92b90c274bab9208");
            when 18715266 => data <= (x"12ac7df57450ac8d", x"515418e2b7f3ba6b", x"b24caf207db575aa", x"bbab3118ccf8ac1d", x"cf7cb3a6da0ee6fe", x"384f6f3dcb15f946", x"3ea4d2cccd99134f", x"3b574eec76662199");
            when 26363076 => data <= (x"4226b637521c36e9", x"3b0074ae6cb18788", x"c3fd80eb7666fd65", x"548bd475d864964b", x"ec1cdd750f147711", x"165bbfed1a9a79d7", x"a73a9b642b00d806", x"a1b0fea22462f086");
            when 5866659 => data <= (x"4946e10de9d7810a", x"33acd3e0992d4518", x"7c32b5ea35c5fd9b", x"896a1402fc4b9fc4", x"b2313a269c094589", x"a0ec9973c6ad2b9a", x"b6c4196ab7fe7f3b", x"fe85ca1b898d6be0");
            when 4329204 => data <= (x"f36cc29d433c8d2d", x"8a709485b2d64d59", x"748d6a5326d52399", x"41737b9fbe460294", x"8c8384c0e24188fe", x"78d32fe919fa091f", x"15c6fdecd814eb35", x"5dd9bde7868aa741");
            when 14509871 => data <= (x"534b96b8ff6e9c0c", x"49f31260a32f2cb7", x"79d690e832a21c21", x"620bf6f142f7deef", x"a5e8a45fc7f52256", x"46f8feeb11c3d6a8", x"63cdef69d566909f", x"a114ffe040ed5dd0");
            when 13613714 => data <= (x"8c85353d943599c4", x"ce0a91dbf8a894a3", x"aaa0789b563c97b6", x"4bf3018d7b93cd64", x"9ca3a81e90695bde", x"d1a87aaf50d6e31c", x"bed93b78cf4e54c6", x"260e373d3c83c4c1");
            when 9779725 => data <= (x"ec3aebee48925f7e", x"fdb48adf8f32fe2f", x"77ae5f54a88964fc", x"89aac857282c5e7a", x"080e448e698fcb9a", x"5303e8110dd1aab4", x"df7cab982a3b343d", x"1a2033ef9bcd9709");
            when 22268491 => data <= (x"5d93b5b8d82c99ce", x"01cb02b2c034cf93", x"cf5a114f54e7542f", x"bb510f22906e12c6", x"b613ecf9ce2a8877", x"6e1fca55714a3361", x"3b7e5d80806ac5d0", x"18b3022dde3b51d3");
            when 20794900 => data <= (x"1048fa3015afae6d", x"90ce3dd81ff6d421", x"712f6bcdca4be840", x"e87e7a22230ad8e1", x"94cf351da1267c1c", x"8d39e502b17c7619", x"d3b2ada4d49e9031", x"c5699ca82fcd01f3");
            when 17789592 => data <= (x"81f73e4bc3c8b652", x"01cce5342759bade", x"95ee2a67e4fbc161", x"ae79286c2f95be4c", x"7c5973b31767f1b3", x"fb088f0a2a395b5e", x"fc14f615a94edc1f", x"35488fb6821a7a2c");
            when 20838262 => data <= (x"cfba7bffd6912b29", x"854dd318f5f22600", x"ab51a5b09a1c9618", x"6b7466a071f25188", x"16156077c575771a", x"f44309e3abbe3441", x"4a0e975ab0d35296", x"c28e700b7b9a722b");
            when 295602 => data <= (x"72e4de236d79996d", x"92675960c6086523", x"ea6c9c44be528356", x"d74cbe84053a1e38", x"d2f643fb6e286620", x"808049d460c83230", x"432313cb70fb1410", x"e5a84dc882587f2c");
            when 3941924 => data <= (x"031ebce9bc3045e6", x"3b91a539e563621e", x"8e7455f91bb562d4", x"0f17e21a8bcd71a5", x"fb842ebbdc77538b", x"449c8f40b8c54499", x"256e2e70d85a4fbf", x"ea5b12199e1a7c6c");
            when 26584594 => data <= (x"4cfc52de1d94c5d8", x"f6b39f91a47f6ac0", x"69642b4fc69f762c", x"486689f606f9e36a", x"1b8532250b7f6123", x"58dd1aec4ce18efa", x"3834296e9b5c1ad3", x"27019ba58c0b6898");
            when 3951874 => data <= (x"42bb1eedb8f38267", x"7db8db4ca5ed9193", x"e24f4969fca932dd", x"0f0d2459f217f9e8", x"0460bec666f9c0bf", x"85c47f5759608dd9", x"3bc5ea7b083ebf13", x"846d0d994428dd2f");
            when 32332391 => data <= (x"6b7520f33bf1619b", x"3ed9b6b35cae88cf", x"3acd2928eb0dc019", x"e2672132e0eb54b1", x"3abe8b6ba35f79c6", x"20e28d0da786b282", x"4f5de484504a75ba", x"c111518c58c26e9b");
            when 33536132 => data <= (x"91cd14a226e948ab", x"ca4bec92c7c4104d", x"4e50d5b92a9d8d3b", x"d2625dfc0140b845", x"fa0facc47a69be0c", x"5170b0128987b560", x"988b39538772d80f", x"870251781a46ee19");
            when 33075413 => data <= (x"2e5f50f636225790", x"12743fd694b06f7b", x"406c18d5020e81e2", x"bef8b2fc229b8b94", x"db9ed302761b2033", x"12ba50d8bd106d40", x"7686969583e82b41", x"85694d89dcc16ee6");
            when 26048763 => data <= (x"6d23cf8d30a4e6f7", x"6c3289e5c4829923", x"3f23ba328a3ad0ad", x"01c5733be954964a", x"828e61966b5f675b", x"c04e9852bae79555", x"661e5265929b3519", x"717f814120a87ab7");
            when 24727117 => data <= (x"5f4f170ac981c340", x"8385eaf70aec3a4a", x"6ab5e5fdf6fb51cc", x"8ecee806309e92a1", x"add0f5eb4b37561c", x"d2e4c122ed1959e5", x"e6a06d1f189805f4", x"ec4659e9a08dd1f6");
            when 16337485 => data <= (x"b9189dc089445287", x"bf692d9499f56452", x"666a279dadf7d6e7", x"b36367541338b715", x"08a0462e4b77701b", x"2b69efc72283f82b", x"27e2c9d4199d6c6a", x"bc861a461f13a21c");
            when 17924927 => data <= (x"21b8659cb24bfc38", x"5b7896e5caad7b04", x"d22082cddd5d4d13", x"8ee68a2ca6344516", x"e5bdb1ec7a191baf", x"414ba68391821dbb", x"19a7d965c2b56487", x"5405c11c16dae025");
            when 10793433 => data <= (x"01b3bf94663c5f7b", x"0262bfac25a64969", x"30e3c640b01f4184", x"f5d6cf8cdeb9fcdc", x"a060cc0085a78b16", x"94a0a36c3c72ddb6", x"104898494bb82178", x"a1405dd92ac52494");
            when 834026 => data <= (x"05c84da8075069da", x"fa44f24a4f3951fb", x"9a9154a4a8f3dc6a", x"2bed78465fa81e94", x"52395bcfab2338f0", x"48ef109355ab3141", x"1e39a3dd9ea4c62c", x"c7f21cdae4795a5e");
            when 16708057 => data <= (x"a36a8c2d5def8265", x"2a4abf8dae939ad0", x"f06a7b110cd6fce1", x"fc411464e0096626", x"2f1291de630871c3", x"6c5ec2abac4f108d", x"cd5634919468e844", x"8d6e5ade42346191");
            when 16044332 => data <= (x"90d4755e0f7fbae1", x"c323c62368193091", x"7056205599049ca9", x"d3cb9674bd55b83c", x"88eda8019b914d6b", x"3e4e5bf73ed42184", x"af549b2ef6859209", x"1a9a925cd16e2c4a");
            when 13014656 => data <= (x"780ea212fbe87e32", x"00d38d922875043d", x"efd6017262d18be5", x"e44f59f14efb9899", x"00ea9b17011596c6", x"cd9e7e57818f15ef", x"89593991dc33ec2c", x"5a861e92ee086700");
            when 30967642 => data <= (x"89eeb6e4ecc2cdfb", x"cbc5aec01e54cef0", x"eec854f5a9089a79", x"6c2dc1b58e5c5160", x"c5d3aebbc7570b63", x"d6cb956da215166a", x"4d8abb96a6b6870f", x"694d6ed5739491a9");
            when 21106701 => data <= (x"f71925ff0e296bc4", x"c9050930febc9597", x"75e4203d2b35c205", x"35c476898c352b0d", x"48a02ae854e3ba1a", x"188519bd152cf423", x"b6043981482c2804", x"29b9e4bbec75bdc4");
            when 84203 => data <= (x"1519e6ef88824d19", x"c113e8226c41fd45", x"f6766226865de9fe", x"057cbd05d1dcf3a8", x"76d15c2dbdb32f02", x"4de15a3bde3f9aee", x"289ae1da82ad2794", x"3bc9d10aabd2b816");
            when 21700364 => data <= (x"e3c55e96b14d90bc", x"7bec0f282951e515", x"e8fd7f729448416b", x"0c996753723255bb", x"85e7fb685af79b7b", x"c34afb974603cf20", x"03b4d2dc79f747fc", x"87a8c82ded7fabf0");
            when 20105655 => data <= (x"f041371c1e59c008", x"f853dc61c570cd62", x"9f4a92e211bef7a5", x"05ffa5c9ebd8f361", x"a48f0eddffc22418", x"f377178db483d5e1", x"8e7bb3d79798a7a8", x"d1fc0a512d7af2c3");
            when 28879207 => data <= (x"b5658fe298b38472", x"b0d1afd6537941ca", x"001baa715d461d70", x"3b873c92ba4dd0ba", x"3e665a8778426f3f", x"f88d45b98477af95", x"23c8aa933df0e1bf", x"0b669ca6e834d869");
            when 17405208 => data <= (x"484853aebcb56289", x"a03be61d9dedf512", x"564f03ae75c6052c", x"e6729879a583f05b", x"284f8ae90923b05e", x"5e7262bf3de43810", x"77a4f77b62133f23", x"ce825f4b9ae98492");
            when 21406220 => data <= (x"77e2813352725480", x"d294cc4477b7bba0", x"a36177b980398c9c", x"d106db7a949a5287", x"7aa0050532175cd4", x"2ecff472bea89acb", x"a07ff7e8339f8b2e", x"91683c2c2beba6d1");
            when 6426024 => data <= (x"c1aa4fae4ad1abfb", x"9d44d1860cd1e39a", x"6ff460ae463a8d98", x"d70e49513c5aac11", x"998b5136a7a6f36c", x"9821840dbabc33cd", x"9ca2fa2ed6372f41", x"cb4679321e748da6");
            when 8553742 => data <= (x"be585ff81f086455", x"8a54985019d9233f", x"96f618bc037359cb", x"b0e2a8407253c381", x"cfc443c1c6411122", x"d3de92145b1a52da", x"7e3c99e9e26d75a2", x"65136502051a2a88");
            when 15708056 => data <= (x"1c40557a2d665da1", x"b6acb78fc68a8697", x"5ac51de53a02c8a0", x"e94470ce81dced9b", x"a87a085bb134a87b", x"df36cb83c9b98618", x"9f5dc05d7ad68526", x"aabbb169d0360fa7");
            when 1770515 => data <= (x"288bd6422699937c", x"83db48784a221049", x"f36154907b3d18e2", x"3945d9d64a84d5c1", x"47c028c33ebefb2f", x"fd233c9d4d82520f", x"4b04e7cf1da42ed5", x"f583f2f93747dc4e");
            when 6449616 => data <= (x"7c79247244f7ce2a", x"bdf4f94308d0bfd9", x"5a4c7e922d45b3a9", x"a4287bb8fb81f65b", x"fb49a8fed04e3c11", x"bb6a2785482f474a", x"2da8fae589880ab2", x"0df85c15b2933ed2");
            when 14204003 => data <= (x"c7e46047c88ea1b8", x"d7ed79c1b1f81835", x"abb848dc0e188b77", x"5a7b99cbc53b308d", x"65d7e2cc08185179", x"fcd1f5bd3e81ca2c", x"4a9a5a4f47b83194", x"81f31c8c4006b09a");
            when 8761535 => data <= (x"7c4e4c22f8b8b061", x"5aeca82c74566af1", x"5daf453eb74c7d91", x"480217ee566850ca", x"bbe5eb6f49ad50c1", x"3ca61239dccb988f", x"9fe43b3a0585bc43", x"97fe6f3f0c53153a");
            when 16967003 => data <= (x"42fc7cc6771a5c8d", x"6e59794f2d98c964", x"8d4d2dc99857cea5", x"2eb247ae0f77da85", x"b51c01bd0c1ae282", x"83ab5a4bf75a09d6", x"98a736dc86bd69d9", x"66eafb18ea2377f7");
            when 21496501 => data <= (x"4795da03938e0aa5", x"12c8d78abb63acff", x"cd52b48b5682f809", x"e1b85653a4ec0054", x"25f2455d73fa31e2", x"0bd8d1706b7e1791", x"41c9e35159264263", x"f220e829ebbd08d9");
            when 6645327 => data <= (x"2998cf397d355050", x"6f37092de6705b2b", x"b79b725d8111e9a5", x"3fd4d0459309da69", x"56705acc1c1dcb69", x"b04d57d2aee3f479", x"e9dafda40df337db", x"10b9273f5b85a135");
            when 25396702 => data <= (x"4d3feac4d8d9adab", x"ddd050447028706a", x"e6661281087e90ce", x"6fc2cb363ac4d6cd", x"3b4aa70637d8dc34", x"d339afb7c74548bb", x"bee4ff5d450490d9", x"1411c46d07b986d9");
            when 21097543 => data <= (x"1e09359a6548ba70", x"76c462cacc0fc981", x"dc0605abc13746a2", x"352f361c852d2116", x"2e46110c2c8818e6", x"1cfc05c309f41826", x"4b04a211c070dd9b", x"e36c000ea5562d46");
            when 11062789 => data <= (x"aa744ed4450ac7b9", x"ec9e044c26f48894", x"8b07d0a0c755d559", x"a5d7702be9f02d03", x"d16008260560ae6c", x"1d52f5d8eafa0ed3", x"f9abfb70402bea34", x"db1f94aeee2279bb");
            when 27468291 => data <= (x"f0e53a3414ee0353", x"d352fde53470ae51", x"c2154ee1f1ee1f11", x"d3390fae10e1b582", x"b4e347aa81119caa", x"96f5ebe540bfb9d8", x"ca60ed85594c91b9", x"e75ab32b1fa753fb");
            when 6993093 => data <= (x"32a591cd623d4b16", x"cf040a67475d9d51", x"0c2e9d843a072c20", x"154165893598f459", x"f92cfc5af085bcfc", x"be7568a3f004343c", x"cc8b56b0f643012d", x"07fbea734d352582");
            when 28141638 => data <= (x"e2562f813d9a1b8f", x"cb155e30a78bf5cb", x"6126279dfcb76e5d", x"afe4545e5ccff4e2", x"4dd4715c6473a89d", x"10d15014183dec9f", x"501cd23ef9f35909", x"ca81e19c35dcc168");
            when 8978713 => data <= (x"c08657789ae28345", x"22173e5fae327c2f", x"d93d020381dbe3fc", x"be5e79701601ba17", x"eb94401488678895", x"671b08cb24381255", x"594c8a04e42683b5", x"b78b3d51cb36e55b");
            when 2208875 => data <= (x"40362cc424eb8ea1", x"e6c99bb71481f45c", x"85d8433a7f1c7dd8", x"bb443f2ab6cd233d", x"8fb0e8c75f34ca4f", x"729a5c185e769991", x"79cc7f1ccdd7dc6c", x"5a30e12f3d70e2fb");
            when 25911541 => data <= (x"2418316e99eb7999", x"ffc89e71256af4b7", x"d7b70dbd4942a138", x"00794df04ba39be1", x"3fcb81d59951578b", x"90a5679e468b13fa", x"1a7acf1df797a0fa", x"d1b15253e3c84a8a");
            when 1731565 => data <= (x"70a1edf84f70c136", x"71f10d4fdc7eced6", x"d8f9e831f9816249", x"e7ee7c19f66609a1", x"7e8f672a6521f59b", x"077aca65a1294400", x"1cef422bf36532b4", x"98a57b121547dff2");
            when 27115504 => data <= (x"30a6f43a51209efc", x"ef3a15623649e2fd", x"43b879a7bd86178e", x"0e230cffee5fe228", x"fceffbd693bc251c", x"3e2efa259f600a9f", x"4b94263f4bb677fa", x"4c3d134aba44ce96");
            when 20271879 => data <= (x"7dcd74a263918478", x"3551b19f80620242", x"b43bc091877dcb44", x"c069bb3f6f9a6677", x"d9a643f4510d730f", x"afb84b952969f266", x"050f62db668ea321", x"97f4423e73731da4");
            when 22258631 => data <= (x"2679666b9d6d16f9", x"b6e7bee051d31f0c", x"53a721f1a0e0fd01", x"dd46ff8f2bc9c94a", x"9207a1420401bd0a", x"4f33f919d246dbbe", x"f67fde90017bf1c6", x"57120ca614b4b4c0");
            when 26641473 => data <= (x"83b04fcf20c76322", x"e34ec2f7d49de9f1", x"e5101b19526c8a28", x"a149fa0e18592cd6", x"bc6f9c74bb5a333c", x"82b7f14e4afb1a8a", x"b6ec50052428e403", x"58cabb19693f6e99");
            when 11224365 => data <= (x"e87b781859c7f7d1", x"586175b5fc6fb192", x"4610ba354d2258d9", x"f62a111bf5051107", x"76406a96484bb817", x"bdc008e1ca25c6ca", x"f50fb53d4bd2c364", x"cc73284828b484ad");
            when 13278213 => data <= (x"06106e0866a962c8", x"962f3556747139dd", x"118757414eba75e7", x"490159a1557e2471", x"f395e8eb0b0be7a6", x"c5e4b4373b6a954e", x"e6cd9d9f0a3bb31e", x"420f29b9efe4e7d3");
            when 24616831 => data <= (x"f9fa3ae5ef4ec091", x"8ec52ee7b07d2ab4", x"5fa607a192e9047e", x"47a2977712b56d23", x"9b7faa735378d0c4", x"a32d040e2c6c7490", x"aadb6d8b1a88bac1", x"d1b3ad3e97450217");
            when 30185619 => data <= (x"977f5be9e55b38a4", x"253e009430897f97", x"6a94bfce25199629", x"307c6d31b2a3a3b9", x"2b3f792a27f701eb", x"68d77cac7e83bbaf", x"93b9fe16365f1149", x"d810fa5f8f987108");
            when 20709317 => data <= (x"2a2289d995d54f7d", x"092a769cb4995901", x"3ad5f98e60aa4170", x"cd07629424980541", x"27c8b4a9da8f12e7", x"f3c51baa5747d57b", x"0c101ace9bc7a435", x"712996112a28184b");
            when 21185376 => data <= (x"fd03ad4df947c711", x"ed99567d55ffdd63", x"4d069bcdd0377dd0", x"ab82ffca193f01ca", x"3c9151a954fbfd4e", x"c080a3d54a9a6a1c", x"2cff7e84ab6018f8", x"b13dc778a98f04bf");
            when 18841401 => data <= (x"53472d86d5a37301", x"76c1847c3ada2917", x"8779cf3b38d8590f", x"cdb9cb50e25765ac", x"add7e21f666334ce", x"c046c700e3e8674f", x"6ee4c48f7e03fd6c", x"65da9c23df5c6782");
            when 21631969 => data <= (x"19805a76e57ef0c2", x"5dcbc37538115e90", x"97ee41e05ff013a9", x"73b73b274c13e0ed", x"62ed0f455e4c2ee8", x"b63ed0c2c92d3a17", x"70933f6b882e2cf8", x"31b23f618bffb33b");
            when 18195310 => data <= (x"4c5505cd5aae2bda", x"d28890f37a7e657a", x"f1a32f35f57c2b02", x"4d125e8c8827463f", x"64b626364339dcc6", x"527c693f726d96aa", x"3ecdb3d56e235903", x"30f00f3c2da2447b");
            when 31393040 => data <= (x"f7b540fd2018bc26", x"a3037a74b8fb5b02", x"b9ac46e6edd5aa9c", x"6dbf20904e5fdf7a", x"e6f9064898246484", x"a7fed3240ba3d4cd", x"5834445e62780eb1", x"39f8372700abb13f");
            when 13535597 => data <= (x"774a907156eca242", x"384734e0385ccf21", x"f9c430791f41f7d1", x"de80919e3e66a0b4", x"ef07cec9d1a163e8", x"f3b4c245bd473818", x"c1ce55f66dc44974", x"fa9be3e933e72c33");
            when 3999151 => data <= (x"a5a40e078251858f", x"992ec9b0f5258950", x"53d189366c4577fc", x"9e15808c230aad60", x"8db9551bee67331e", x"b78a144c8a20e2ca", x"211c0c484d683914", x"2d756a8e737a71de");
            when 18004888 => data <= (x"3dad7c8aae256c5e", x"8dc8499cb87d8451", x"038c152a48e70da3", x"3c8239b45422f696", x"6f804777a12cebf2", x"9d99cb474006fb65", x"0771ed4fa49f6da5", x"c49b46408f7bcac0");
            when 1517452 => data <= (x"f51eb387f246b426", x"67de514fa4f80058", x"405914a648cb3e28", x"d4eb364a215c608b", x"f35750dbb4df71b2", x"1a82c9e1ef9341b2", x"801b428ed35ba298", x"124900aada539ba6");
            when 26599318 => data <= (x"477351ee551d4ba9", x"e9aafa78cefb0afc", x"f9e2a5823b768776", x"cbf55a05e6a24db9", x"1ffec2edce0c0ff5", x"44237e50aa9ad87e", x"88a834583f84c859", x"bbd7c49059f91705");
            when 6267800 => data <= (x"e7993c2a4f71cf11", x"498668dd4093bd6c", x"656c517341f37dac", x"74da01f5b1991088", x"7e16ed1a0bbb1fef", x"6da5c449ea32bd68", x"53298f3366496b9d", x"ebdfeaab00af822e");
            when 19636291 => data <= (x"fbdb65f113424639", x"263cdcd856a797ab", x"acfc5da79f36b3c7", x"c7a9c1f295f9cd9c", x"74c31c4078738745", x"abce88d89e731cb2", x"df86cefab46f34be", x"c5a75f5f5e4d32d4");
            when 12274110 => data <= (x"26b2988a2b692c2c", x"f6e4a42a54d46349", x"555ba858229d2160", x"bc0e6eed300f456e", x"157fc3af8b570236", x"84d40b14fb7b6704", x"c7e44ecc9b5f418d", x"9283adc21fb862f2");
            when 22146999 => data <= (x"b1422eb89f0e1bb7", x"4e9a8a1322fd7251", x"a1bca6daaeb1a368", x"0e71a480d0402ef8", x"0d1db6f85a8a4871", x"84404ad372a12fb4", x"7c7bd8ca943eaad9", x"e8509e111fe7d3f3");
            when 28014837 => data <= (x"2eb80b615e22717f", x"7791da78fb2b40ce", x"1c6f2fede030ac58", x"8377a2c138276f68", x"3de2dfb454278e78", x"03e4e9e62a253469", x"deedd6e4d34683b0", x"fb1e60bedca9fccb");
            when 30489449 => data <= (x"081ace0228bc6a35", x"dd02f19f27e49ddd", x"d6d54c1b14ff7b79", x"dca5414b68ae15f0", x"9442a2c2b2288551", x"72c173dc58ac34d4", x"d5dfdd299d0360b7", x"814dc14dc0a405ca");
            when 3320752 => data <= (x"b4141c1e0669fea2", x"0ee5d1be75750ceb", x"ec444561b3d3d4c8", x"8448dfeaecd5711d", x"398c53a462378b20", x"0d68e5fd8be97d48", x"e4489aa84cea850c", x"bad061e89141ae3b");
            when 22891482 => data <= (x"7ac1a8a299992326", x"2c109c1923bf72dd", x"16868786b1157bb6", x"8891ebdcf2e70b53", x"ba040ea9c9580688", x"c5baa38d585f9d78", x"5f08834a601ac23c", x"24860156e0985882");
            when 3439025 => data <= (x"52c81fab7909d45f", x"6cc896981ae12f7d", x"55bc77e0f232a55d", x"000b596f7f85311b", x"0d91eb11955d7903", x"976727bf809baa1f", x"d87bcd415ba5977b", x"5ae640408aa2bd97");
            when 6422408 => data <= (x"1074a32e5868257e", x"72926c5c263fe9be", x"af16b4179adb6d30", x"fb92b8ff0b750134", x"523c56b127877eab", x"c56d3b223377b439", x"fec3672dddb7ac4a", x"85cbfa4a25b5120b");
            when 29234685 => data <= (x"394c786b96b239de", x"77ef2f5e61020857", x"d29196f86519af89", x"3c03a3d4da84454a", x"f029cc5cc15d4411", x"35b715946ddf8ae3", x"d9c274cd5a0daa0b", x"0f2786faaf63d9e3");
            when 18139245 => data <= (x"1181bf148d5b7c4b", x"433c3d61a531a45b", x"8c536c5e812dde73", x"315d5d1b4c4b6375", x"a9cba78528bc17d4", x"f85a51cfa7264a3d", x"88b9aa69da9e5f18", x"07c66df85008ed7a");
            when 10169951 => data <= (x"6d7ddcabdbf17a64", x"f093ff29de52514b", x"5367c7ccb520efcc", x"cbd10941f3bebcd0", x"8410251658c76ef1", x"46057bc13b27b16c", x"df911761ad9d58cc", x"552e77509135ec16");
            when 10954308 => data <= (x"5b2783b927e25315", x"56ffa885fdda2144", x"4defd164a492c939", x"73d485d964d1abc6", x"5cddccf541843f0f", x"0fd38bc3ef4380ac", x"ba6acb3ac96481b6", x"196a7b620535b0d1");
            when 19065900 => data <= (x"8e764ef7d2b3c9ce", x"1b70e730369d4c7c", x"4dfc9d85bdd8b910", x"9766c33126ec9996", x"6faf3ddf8525f323", x"b66cd4b4f50e9002", x"74e0e90cd0dcfb24", x"1ee2c70841bbc916");
            when 13276385 => data <= (x"a31fc3149aa7189f", x"ca8e5474dd222680", x"02b8dfe51ee975f4", x"212eb866bb3f1b11", x"100739046506dff3", x"fb789168231cc607", x"297a8306c9d3e8dd", x"da09bc78eb61013a");
            when 31108461 => data <= (x"b9c980f22c1a371c", x"9ceb08f7868b4757", x"0d0e280fad43f588", x"0cef810d7529aa1a", x"b040901bd6d8492c", x"55b790fc368ce4c6", x"fbaad5a0cec2731a", x"905d8e8b39d554ec");
            when 16621123 => data <= (x"265e8828656d83a3", x"74871229ba1acc89", x"ab057ea1a6914ccb", x"7c71334f593860ec", x"af898499b77437e7", x"2ad5ea1634c234d5", x"edd53f3a59a036f5", x"c9880214e894a82b");
            when 9018052 => data <= (x"99984eb8188a9c2d", x"7032fa9b0bd3c2ea", x"3630bf8a3dd9e8c4", x"b41288e6b0a6c237", x"49adae9e714d4855", x"d6318405c3ff53ed", x"a35af66b3c6340e0", x"4b45b8aafa2b729c");
            when 25507705 => data <= (x"226e6d6d61387e56", x"e3c637700ef4fbfb", x"78b2a4e872d56f6e", x"626bfc161a8af9a3", x"47037057965466ad", x"9826a0e2e4a8325f", x"53c744286509d906", x"5092b96f6f7f0c2b");
            when 13591160 => data <= (x"e7f7111a623a56cd", x"22ffad482e5667b4", x"357637219a5538db", x"a19cde77457673cc", x"7f19a68bfff52f9d", x"683e25b8b2303186", x"44fa13e2a9569202", x"7633be5d73c6d5fb");
            when 8775617 => data <= (x"4bac49413de51cbf", x"096f62d02f38231f", x"b85ebaecaf8a4fa6", x"7e4fd81026b9428f", x"3d4db248dd662d90", x"cdc6428c8bc6926a", x"5b0b2b368aa378d2", x"952790d76159a0d4");
            when 11850771 => data <= (x"b9236d4ab294b70e", x"24b217a4272e6e95", x"5957fd0b03564785", x"2bf4bf0f477fb039", x"2e0bb2c3d2b609c7", x"a087392e4b5d5ca0", x"6373f9a59257b6e9", x"ddd03182f80199cc");
            when 4389361 => data <= (x"71232caf5e3d5c29", x"56669c52d62ee898", x"b2755d35a81acc22", x"d0e8f9d4b64080f6", x"477ba9b99d87f3ef", x"f90228f9bae97b42", x"8af43752a49aba50", x"aeb3cc236c615abc");
            when 8408581 => data <= (x"b91085b0ec783f82", x"39fe63f6b27cbdc6", x"578f9a08b8a76c8c", x"149bcf537a651c4b", x"5f00d75d02a13ee2", x"88d8d7c63d09a65e", x"21d063a295d008ad", x"3273fb43c4d7bf72");
            when 14603796 => data <= (x"c8ba8057719039c4", x"7350c2a6bf94d9ff", x"b38451f7c7dd3c2b", x"5f7d7159ad13c901", x"a4f84f4fd704134c", x"bf54a557b632fd38", x"6b3cddcb57dc3e16", x"e15063f758ec9598");
            when 27820172 => data <= (x"e96991294918d365", x"4cf684077dc3740e", x"ecde66a377b51018", x"2fdc721e38f4e454", x"89785f58a632d2b6", x"2579656361fc9fa5", x"2185ddc20eb4c1d7", x"6b8e3d560bb2e5d2");
            when 17215359 => data <= (x"bcdd40ddd1c1ec1d", x"568e56c692c60d6c", x"7ecb89e351eac215", x"e414b2d58433dbed", x"390d7feadcccec29", x"19075507bd4a3b6d", x"3590d17d5a11617a", x"87e33acc8624a15a");
            when 12236812 => data <= (x"a59fcca6889be667", x"57c49e7ea86458fd", x"b70312ba0a55f3d8", x"d0bb7dea4c4011d6", x"da76a879be8b7caa", x"4838704b6550fa48", x"f3755925ddfefb25", x"70a078b7ccc46581");
            when 7074029 => data <= (x"9041d860c2c6452c", x"1dee996c09ee1fc0", x"f92a9a5fc5108fb9", x"a31d2fe523020d2e", x"9b19a0ef871584d7", x"d156f4767d1c7886", x"c225e0620a68969f", x"701a48296756df92");
            when 15324145 => data <= (x"4d72211f1ef32591", x"8ae37d60293b6855", x"3049d293aabafc28", x"cc498eb119dea147", x"5dd43845391645c0", x"464ce2dc02167c2c", x"b5ad4818b97139fb", x"6c9782885aa5b097");
            when 12580536 => data <= (x"8d9356b61c03e3b1", x"49c29ae968f6de20", x"d25d7b7b88817384", x"ae7b382221c80120", x"0ab24e3299937b18", x"91b6e299678717b6", x"3f9026426af0e89c", x"319ac5dd79e17b5b");
            when 7494450 => data <= (x"b290a4ccdb56a02e", x"b47adf7a5b7888be", x"69aad49b944654a3", x"4e5b083feca9b1c6", x"e8ab396279b75fb5", x"dfdb590eb45722fc", x"3b00a5ef089dd6d6", x"391a4d7ff19f7bc4");
            when 26562708 => data <= (x"e9c97258f6b008b7", x"9dc088b2f6228067", x"7c91fff02b95e3c9", x"c0cd4a09361808cb", x"1ce91ddccbd157c8", x"e9f26cdc95ac3d99", x"ebe244d8179f8abe", x"0d9ca30e737781f3");
            when 21773389 => data <= (x"ff169ac4ef1f57c5", x"cfda398a0f8865eb", x"43f34db580384d18", x"d455db8efd8330a0", x"49900aec9e9ee074", x"9064e98a2d5e13e9", x"8f5b4fb100397a7d", x"c4fdf4a6cf5e21e9");
            when 4994700 => data <= (x"2012f5cc6431aa71", x"a25bf0b5cd9fcebc", x"066e6990eb2f3eb5", x"cf005f8c3d9a3d10", x"ac7a0662052a5d72", x"01ed89349c9d6f27", x"96de4d65003ca207", x"ac575454d5d923e3");
            when 8959869 => data <= (x"d4ad81560e9b3813", x"d8d647521c74833e", x"79ebf3531b71ab24", x"8112fed431bdc018", x"bc7b0cfdfca30560", x"3307e149ccacb14f", x"7a40f74adbcabb1f", x"06f6ac79f0f4d06b");
            when 18275881 => data <= (x"edf79e12267b733d", x"f5d97a2226ed3c2c", x"99193d0b1c552d70", x"10f38f8db4c6720d", x"a9bd2a960585c909", x"b653f9f7e62ae536", x"23dc557585f1f9bf", x"bb5de2b3fbbd2f97");
            when 13071983 => data <= (x"0b6091ea4d7b3c5e", x"d4438143fe640555", x"3d12e86d80f0610b", x"3a94b367c8e08f7f", x"2a150a85c9635fd9", x"b3a13145afd17440", x"b2312f9619edb364", x"aa0d1128ba23ce79");
            when 24247312 => data <= (x"5c3a484b5444eb7e", x"5a47d62b9641d67b", x"c76045e7495c93c3", x"097ab555d7960b34", x"11431aeea1b2bd77", x"54c127c0309e1d2e", x"00f68691523d1f6d", x"77645f73c92ca797");
            when 16199386 => data <= (x"e9677f7fae1adb70", x"e98918d908a34f62", x"24188ff4164881e4", x"f302ebb11453d22c", x"e48b4f4291e5ca0b", x"a75bc52c580012a6", x"a34622ee0e9108ab", x"c497cda6e35ace9d");
            when 17918577 => data <= (x"d4a2850f6d2cbf7e", x"52d1762d41fab0aa", x"e02ad4d338b512f1", x"68352f5b1a71c1ca", x"0f157ae76ca07ffc", x"cc97172060ae6821", x"e327102a1d6ee785", x"222f848802e493b2");
            when 8827854 => data <= (x"6e40458423cbe0c6", x"0030fcb13c116269", x"c503c2390966bb22", x"dd0486b0360d9c37", x"1f41ecb31b28866b", x"6e5ac351d044b220", x"d82ce6d69a723458", x"aa99996ef9ae0043");
            when 24130734 => data <= (x"17937d21faee52f9", x"6551225b38197a28", x"cd8b96c097c2c473", x"5a3a91f6fdfd3840", x"a2f6d669e4a66500", x"75a85abb475d7dbb", x"99f69a9aa23947c6", x"4579fbc46036370c");
            when 33172890 => data <= (x"f24b35aaa69f7c45", x"8371dbb9e8f2a495", x"f34819b3da616af5", x"f41063871336c449", x"c377ce3b6446c9d3", x"8b2d6bb3fa18f83a", x"3017c2f1bfba39b4", x"a1fa6521133e0c0d");
            when 4445102 => data <= (x"404a7577b171366c", x"c0f6d3a6582e3495", x"7cbee541c2ca4ddf", x"563cfc849c7ab84e", x"38dee7278131d7c7", x"9ec21ccbe2100c96", x"6587735aa4542b03", x"6a918c5d0d870430");
            when 6347118 => data <= (x"b8a78699c0750a48", x"bd61ee605f21710b", x"8930b615ee7708cc", x"ade1b1238a5ee75d", x"be41baf901c1a0b2", x"3978ddffcee3a1b0", x"568d6b23b49fcf81", x"3e8417abe88b449c");
            when 7840357 => data <= (x"bdb5d833636e7852", x"222c55e198e4ba8f", x"a3fc9052262158fe", x"6549c8ac9e8bd167", x"cd2afb760f699865", x"3888ff93e17687ba", x"bfaf0fac63a4a111", x"92d94b19ac1afdd6");
            when 17553876 => data <= (x"a39179212d6d3175", x"57f24aff649ef24b", x"91385385607f0a5c", x"9ab5304f3870bccb", x"80a82e0d8cdfa32f", x"6edd803097b23a1a", x"259b5ff83f00c55c", x"a0a5783c40fb5f55");
            when 13515462 => data <= (x"36b4ab5804647e14", x"b79f5dc5ed6af748", x"19b12b9f2569de88", x"74c7bc7b8784f592", x"82e6ccb910754688", x"ef28692bc5b54526", x"080eed68bb8d829b", x"889f4f961768e21c");
            when 18006024 => data <= (x"afd62da5bf190233", x"0d3846c2614b042f", x"10a0cb7fcfb3afb0", x"72da2cd995d3c545", x"1a4a220baf0ba174", x"31a175a24a36c173", x"bcd11fead718e08e", x"c5b1df0f5529b66f");
            when 28845422 => data <= (x"2a272dc322d278d3", x"1b2dd534b7d8d29f", x"4ef36c2e9a73894b", x"3ab3d4830fbf2e5b", x"f684f17481263475", x"8aac8a89917fcfe7", x"c408fc297cbde477", x"4e7cb9018ddae9dc");
            when 29086534 => data <= (x"80b3e62e73d96672", x"2ab532758254b0b7", x"d7f6956118cc5521", x"00720acbd8cc354b", x"c8ffa967265b6ef2", x"83d256fd5795cde1", x"48480ff40859e4eb", x"be2f23063a68ae9d");
            when 22052987 => data <= (x"3b69c5417561f74b", x"a10c834e5f54fbde", x"1aae40b9be1a2fb7", x"a214637081324c5f", x"48bb0c39ba04a26d", x"6163da8e30417d50", x"5854df6447b604f8", x"bf688385e8117580");
            when 26650040 => data <= (x"dd127176b282fa6b", x"c0c548fd55e9bd5e", x"1e2f21984008a79d", x"91f8203989383189", x"7698e7bafacfbc34", x"25287cacce3de178", x"eaa728d2757ff6a1", x"ba36e009fc7fdbd4");
            when 6499182 => data <= (x"e050e00011433182", x"b7b1ae15f42b5d5b", x"b2585f302cee1b2e", x"889a2cac825992e7", x"d303a1144aaaa5e8", x"d69d049badc0e767", x"74e0fa4c53d30cbe", x"13a4be432f1c1c85");
            when 6861741 => data <= (x"cbd0c88077e9992f", x"33d207247cfd277d", x"0f48be0a97ab3268", x"7b44209105e2502a", x"ad1f45b2c2e85be4", x"e5ed2ebc093436cb", x"1711542433b9c02b", x"f53a91b27ce03f38");
            when 742990 => data <= (x"7c73d5b8195643ec", x"c6c9041b4a15b8f2", x"756a96c82e77e0e9", x"bc7b99f2dd410623", x"94b4efa85d66cd59", x"f9314f00df100cf8", x"7b2dadcbfa517c75", x"9a24c5cb4d796cec");
            when 11271712 => data <= (x"13464ee758b3e2da", x"ad31317cc0ecd107", x"24a88ea97a15338c", x"a194c3a091433054", x"ffc4e70afc368fa0", x"37fd08d5c524189d", x"06bb5c9559f2b781", x"506726878c97ce89");
            when 8549326 => data <= (x"205dbe5dd35633d0", x"739758ad1587e654", x"59e495ae952ea280", x"ed9c9aea41f68db0", x"eea24ba2adf1a014", x"0ddde6bc551bb5ac", x"e0cdc790b04f8e95", x"b7bb01629b4cdeb7");
            when 7480274 => data <= (x"a9899d45977b3e72", x"38853a667cab36a2", x"1bef853e8a8f1490", x"94d7c04ab77b5951", x"0fe56fc51f65e6b7", x"53eecdfdad05d8c8", x"6b83dadd8c9fc0a8", x"41c4594d0c4806f1");
            when 18128380 => data <= (x"044cb2ac20cbbf0e", x"3cab5349426d1b94", x"599c4d5441e31509", x"6ed1aad224b10e26", x"17f1d976ea7b0a8e", x"ee46cf27737835d3", x"981afaeb61169388", x"62df5da7c39ec065");
            when 25946408 => data <= (x"b4c02117aa8672a8", x"a02773fc03aa5269", x"c5d3b07b24bfd688", x"072514a4faf07504", x"5dd1b09fe5247155", x"02b1ca455e9a9c4f", x"c9dc8831ab2e5543", x"f565dc94acba48fb");
            when 21058257 => data <= (x"1c9447e39ae5a2ed", x"5636ef95be4c9f92", x"3e27304918171d0b", x"1ffee991b689885c", x"a85468c17875b0b2", x"24216baa3dbfcdb3", x"8bc35444f2fad5e3", x"90e4f7982376ff8a");
            when 12948414 => data <= (x"bf3d79db376f2e38", x"3de276f9a6219a40", x"9ce813de4eaaa55c", x"d3eed8954af56f59", x"79f6e894056e1518", x"c15eaf99f582888f", x"ce8c68db6cb1e8c1", x"b0c707eb38b0210a");
            when 18263214 => data <= (x"bbf1f475c353316f", x"ccac827ad34d790f", x"28a60cae83013d4b", x"6f898086801aa2f9", x"5ebb8ca089bab75d", x"90d845fdc3bc46a1", x"bcff0ab7ad8212e3", x"b6b0b4e0c34dda00");
            when 20757331 => data <= (x"af260798637e17bd", x"6640d6d2050ff94c", x"1c17d5a44c6df879", x"fc09e12d127c4be9", x"7cf22b05c0c8c01d", x"7ff6cf2bfa08182a", x"e5d17dce50e00377", x"3b31e9a338f2b107");
            when 25216174 => data <= (x"2aebe797785f4248", x"efccf083600834ce", x"105bbfb5c7748e7e", x"dc45f6b6843b4aef", x"0663e322e8eea5d3", x"2e0b27b16dd0b0b8", x"a04be61e8553acb0", x"a1c2fc1e3ed7936c");
            when 14212452 => data <= (x"0e71068f5490df10", x"6599dd1507f9e6ac", x"e1a193ea02567df3", x"2ca0d97e22d462d6", x"7b49d016a7a99862", x"c14b833eacac0f4c", x"8d4b9d481f3ae18d", x"ec5263724348576a");
            when 2102954 => data <= (x"e6bb0aebfc6c58bd", x"f073c5ed80317011", x"8d7e7cdc085387bc", x"3c6064a12981fd5d", x"b4bd6d2c5b1b4509", x"2a6c44497c6a30a9", x"a9034ac60e1986b9", x"4b3c7c804a37aa88");
            when 30420572 => data <= (x"aa908c40ace93903", x"18efb5439c2b8c86", x"76332fbc214a22ec", x"0e7faff73c253653", x"7a6e1ae74d3a2b8d", x"aaf52432dee96cbe", x"a5634f18815cbaf5", x"0b23e947eefc86e0");
            when 12306448 => data <= (x"6bf9506d6c7aa0ec", x"0b18ac2f70269a8a", x"3d3108000c9e8fce", x"02320701c0939ef4", x"5db9708f276aac7e", x"a8d3b83280423957", x"98f5c24e8be4b033", x"864f92e9ee3e42c5");
            when 24286232 => data <= (x"621601754648c0cb", x"e2bfe4f1f9dc426a", x"f9e66d32d987f0f4", x"f5251c3a3344f303", x"3b9dda1bd77b4156", x"f13a86f2aff4e6a9", x"ba9749c8027280fb", x"5cd52b4082a6cb83");
            when 10103039 => data <= (x"cc983e5e831ed6a0", x"778f8251b83e1d29", x"3269635845bad0e3", x"83a1b4552075c2b0", x"36ca83e27bd8253f", x"492b3ad4cb08133f", x"bcdc784d8d76b028", x"8b6a0be54f42d00e");
            when 12890466 => data <= (x"ae4507fdeb2fab75", x"78a20a4f0adf20f7", x"1cfd43d8f9c56f78", x"2ac256e22b309dec", x"099a449cbbeb5eb6", x"8823867ac3619804", x"e624c163aaff6884", x"d36ecced112c670f");
            when 17385201 => data <= (x"7ce5221dd0f6edb6", x"a0e1fa48315b3697", x"20575a0613bb2979", x"8e471989f60dafe8", x"cc5f1edeee6037bb", x"ac0c75c2dd1d9204", x"7f0f38d5bfedf882", x"40e2c25c34365f68");
            when 12331849 => data <= (x"354de295a817e942", x"377ac167f38e6572", x"1ba658a76cee064a", x"05362c3a1a1f2097", x"4694b9c9526015b2", x"818f9a6a8f8488ef", x"a8242089b4742577", x"c8f38b83b7846629");
            when 7183253 => data <= (x"fd82b4ff1232acb9", x"c4fac1de09ea93aa", x"5d95554a4cdc3d62", x"e810191f6ec7faa2", x"3e4402d9b7fd3e58", x"d653bbf48c0b25d9", x"39bd97a8f38307b5", x"eb73d257a44aabc3");
            when 5202464 => data <= (x"8c952bff15ead44d", x"d632603f0cfcf632", x"e3b288570e73a42b", x"bd1e168a5f2ae188", x"8ccd0a6992b3f7bb", x"180491b863fdb9b5", x"0f1726eb74eb0837", x"f64876b658a472d3");
            when 3660823 => data <= (x"30708166452477ac", x"312ecc44fd43af28", x"e4e8d17099c02884", x"b41a8e42f1092d97", x"99c23a0ab6130851", x"2e8c9305f96f8485", x"976c61fd1c78f655", x"2556ac3ce3907b5d");
            when 5255830 => data <= (x"fdf8c60d28065900", x"785550b9eb40c192", x"d653621b8dfd3bd5", x"509af86436f58f2e", x"eec6134aad6c4452", x"ef49fd1294605183", x"80067d78e77fcc9b", x"7b23cb54f3b243bf");
            when 10901134 => data <= (x"a4ebfda882cdf290", x"ac57a81333c65e4a", x"20230bb489ad2b2e", x"531616b5ee49dde4", x"340f87b157a5e291", x"8bf73942bce909e6", x"25c3a22856912266", x"681c8c21956f622e");
            when 23475768 => data <= (x"05085867554dbb18", x"6d5402b951bc2d68", x"868307d0ca3fbb4c", x"ee3229a5c0ab6d04", x"b4023ddfeb250290", x"de817fa18ff7d739", x"b589f21c8b70d626", x"8fe28de8301cca3d");
            when 14766155 => data <= (x"a6e90a2dc2e994f9", x"bedecd3649d0a987", x"7749cb84b765d474", x"6aff477d6bcbd711", x"60ff1b4b574a4323", x"30ecc20c7ce47751", x"d68302326eb4edc4", x"7b2bae352950f73e");
            when 8900114 => data <= (x"d018b34833b8ce92", x"9de7271a7fb4b3f9", x"615239fa736b2fa4", x"ffa39a94b8128e78", x"0553908f1c08678e", x"0236851f8fc176b7", x"3f8f5383af973fa1", x"c5777e43e5df3245");
            when 18859134 => data <= (x"dd7ecccf326edc60", x"740248b4d1417bc8", x"25ff5e706df1f039", x"cf31c82f8471f858", x"c281f14a3cbf5685", x"eeee9f6840baca42", x"c3b411ad6f5098b1", x"e041907bc670f252");
            when 31289483 => data <= (x"5099f498d76a4059", x"de8ec9b2b62c942e", x"1980364e608b439f", x"db277d3064a52121", x"a89094a53bfd62bb", x"0d730e295f54ef95", x"5662433ee4efb07f", x"1cbbcfca62c45932");
            when 28035317 => data <= (x"0408e8d3053dd99d", x"a4ca0129527d5b34", x"acbda273a4b8b04c", x"bb55187e9c4a7ca9", x"4f99e622bca8dddd", x"a76a75fcc03fc625", x"c41571ca99760395", x"9216bf3f2fe07a6d");
            when 29655006 => data <= (x"fed30ea4452793e9", x"e1b93d7e82a10cd5", x"82383be744ae5c1d", x"a5e5ebd3bbf9a16d", x"0bee2d476896fc20", x"8f564d580f378827", x"3e3e4d6dd00ce7ad", x"59025f158a0089a3");
            when 2875868 => data <= (x"57bce9acf793c28f", x"af04b6e00b6d87ef", x"33d4d4510c3e7ad1", x"f84d41b5c8e3be63", x"48d38e8c6d6b9ceb", x"cd20a4a1c66233e9", x"31634f2b1ebc6eb3", x"0f82f911b9294190");
            when 22347309 => data <= (x"920833ef4ff59010", x"aac2ba3ef5774b77", x"e244f72965b26610", x"8cd1e3c1313252ff", x"099f4a079716c03d", x"8bccfa5c6a1aea02", x"0c1a8ebbc4dc7b19", x"a966257c53017ef9");
            when 11548651 => data <= (x"f2f67fb3f8ad6eb3", x"2fa8a37c90506e5c", x"6ced1c6b3b9049ab", x"edf37e79ee943516", x"8e82b63e23bcc83e", x"732e47fc822f9ae1", x"ac64d5fdae4451e8", x"6537457460795e31");
            when 31448017 => data <= (x"a5e8176b65f69955", x"9b2af4c28fdaa81e", x"297a5dc4e463f829", x"08c2be10b7d62573", x"e2dfb7c5b07960a5", x"43539596dab9eff1", x"a47c697f83101b3a", x"cdb354514d6cec48");
            when 31775538 => data <= (x"96b2f9895ff6daf3", x"ee80d6fe910bf0fc", x"d62ddb34ea9c8d9f", x"1d3085f7edda9e24", x"7c1b769e7c308fed", x"4882cd99b007bbb0", x"2ec51e6b8eca1007", x"4a3b71b6f8106aba");
            when 21176797 => data <= (x"55b7033c659f350a", x"825e2ceb9b4034ce", x"d6e2244b772af50f", x"0e032fa2ebdc3501", x"c7c742903a087db8", x"7e884437ddaed0ac", x"0a854877783fc6d8", x"0a81b656755a64e4");
            when 22276029 => data <= (x"9cb71f0d4dcd0b09", x"5183a2380933ade5", x"9f7c71d8e4531c30", x"cc0a25ce4a771e5e", x"eb89242667f43cf4", x"87f587d4f0a28ff0", x"9ad2956c90dfc86e", x"a7c8abb724fe7965");
            when 32347235 => data <= (x"4f7e433c4eb4d5ee", x"8bcf9b4f22fbfba3", x"6a340ebd06a4cb4e", x"bc0456dee7535464", x"ea1a5ca859984845", x"399f0b1617f0f4ad", x"5495214e8414f63a", x"bdb5e25ac80df9d4");
            when 25038963 => data <= (x"df445bd950b64c1e", x"bf1205e8fcc333c3", x"b4cb3f5130024836", x"96491d68e99a2db0", x"1204e2d56eca2faa", x"f34f557938cfcb35", x"907ef2eb3d2ae042", x"f82fedff93052461");
            when 22933188 => data <= (x"efe456f26d841b95", x"785dec85804db2d7", x"836a02b8cf3d6708", x"c83896d5e4694337", x"8d9504b3209ecc52", x"54b5bc9507d38a1b", x"874e16e92daaef1c", x"a0db95f44c46a94c");
            when 133047 => data <= (x"10e1ac652bafaf19", x"f83fbd3cfa073976", x"822296e199417e95", x"b94e7ddaa81b0fa5", x"bc164a39e9709460", x"d737b0ceeb9f5278", x"3f9d3936a711a3d0", x"194a34c6217f11d9");
            when 15100591 => data <= (x"11ad9157d54b0f33", x"c4a7f95a74e8b70e", x"aee3843453f89bfb", x"cde74c729d8e9d7b", x"c36d679d69395111", x"56fae74d8c63e659", x"9cd7075047620d09", x"064fe2681b30c770");
            when 23056729 => data <= (x"489bfca51f11fb78", x"720ce572d52c55cb", x"95a38064cf32ac5d", x"1a7fe9f4e2b4a1af", x"eb089d451ab40ccf", x"e20ee73021cd679c", x"f25173b4a639c1b9", x"59e0406570b705c0");
            when 19469287 => data <= (x"ab9c396b24567b2d", x"a443171c6db49208", x"001c47c74a181203", x"0c5257828d55e38d", x"c88ecfb03d9b18ed", x"c7d2e115f6132655", x"b3d1e25951bf5466", x"391450d8bd91a495");
            when 1899002 => data <= (x"4c722291f31fb432", x"f82ad3a5a72b37eb", x"8f43b7f60b82137c", x"8ee0a4389869af2d", x"5b076f958048aece", x"2b339e5c1098cbd1", x"b2f598375c9d980b", x"df783d7c0f5a3410");
            when 14972622 => data <= (x"cea588b4b3c146ed", x"c775a79dee925f89", x"b8399c4af2831f2d", x"2c6b56e72a06b6c6", x"88ed03dcee08c4a3", x"2dde3fe2b2419a4e", x"2f60f63ce485a8bb", x"bdb3186497a52a1d");
            when 27593464 => data <= (x"3ee30da5ed6e8958", x"94346fcc904b114d", x"ba91835d72d1d30e", x"d3cb1814cdb6347a", x"efcea9e09955a181", x"247f741bd482221f", x"b7851f3587a617ca", x"481582723a8eaed8");
            when 3783014 => data <= (x"920fcc464cab700e", x"33654888eccf3ab6", x"b1ab83885559a75e", x"83b71b58910ad445", x"4e95db7f92ba2e6c", x"3e6d4c3061410b1d", x"819e775da7304721", x"283d9c9e0335c4b5");
            when 23388505 => data <= (x"8b5b61529d4dc2ff", x"0cbaca46fc0d2164", x"461e36cd38643cfb", x"0ac95ee8ddec31c7", x"d17edc9078c1c6d3", x"f7181699a94e0a2b", x"e1b9deaef55794da", x"179263c03512d55a");
            when 5809379 => data <= (x"88c54481f62678df", x"1f5d504715580ba6", x"9c89fd2d12a1f567", x"9faa382860827203", x"5c1b99957ec93811", x"a16a5280705935d4", x"89eabb268b62f72c", x"d1c7f2d01bf5a0e7");
            when 4332126 => data <= (x"a4fdf8aa5b84991f", x"516c7976ae41d9f1", x"000b8f6a90104705", x"27d66a8a0eb36bf5", x"9d36440ddc90d1b6", x"17a956c964de3abc", x"c97af0490bcb4ea7", x"f6d002109b3cddfc");
            when 2532148 => data <= (x"f763c26d709a513f", x"264c551f9eb6df35", x"a30ee6340438a016", x"73c74f52683563db", x"d6a40c2858846001", x"85745f3c50f23940", x"f8510e2d1959df72", x"5bfde4d07667cbee");
            when 29677218 => data <= (x"81bedc64f36e32bc", x"8b034396fe76ca2f", x"599d907b2565dc65", x"97b40ae174d4660e", x"48b8e0b9bdddab8f", x"5e13437e89a3750c", x"d158114c0a3a714b", x"4815578cd2fc3d96");
            when 5781298 => data <= (x"78a0a8b98a543125", x"0b0934213e73f7d2", x"8420f8c8bf80bb9f", x"ec7a5c78031d0204", x"126747ec53350715", x"33cc33cda99325a9", x"6efc5cb80234fe4d", x"cd00f62d0aa01989");
            when 21031457 => data <= (x"c83ac25860b92ac4", x"ce409a1036dbf3e2", x"6f7977cb01181604", x"4a1a7b0b816146c7", x"bcddcdf70cada48a", x"0abdeffcc3c2959e", x"bcf7794cb8d09fe9", x"4d144c799d2fc007");
            when 25578879 => data <= (x"cad6eb3ca676a7c6", x"671b1d166622dcf6", x"871c57e9e7bdc571", x"8ea9fa29bfbd3f7d", x"09ffc55867ce14da", x"595b1ba94c1199fa", x"5f9d7f8302fa0426", x"50d277e9bca17e35");
            when 9957199 => data <= (x"afbb297edcf76b1d", x"18095165a5204d34", x"8dfaa977e65ef9bd", x"a803452e908c8bec", x"18ee04e17295499e", x"22bcb3a0581231aa", x"219e50eba5a2d997", x"17d4a2325a6cb51a");
            when 9976269 => data <= (x"dd4e05632bdd59e3", x"bc4ce3d9847dd791", x"2c5afac7fbbffdb0", x"f46ede48ea39b619", x"85cf3860936d9b7a", x"bb109b1a0159d715", x"549bb392f174a9f3", x"cc20f005f5934862");
            when 26020812 => data <= (x"76fdc4773f60276c", x"d11ac0cdc53bd7d1", x"ec66469cf89cfa0c", x"ae19559c57847285", x"fe53d3a5cba4e504", x"6692498ca72a5e0b", x"38e611abf9b0abea", x"e5c39d9a015ffabf");
            when 31284873 => data <= (x"84de91b2f8254db5", x"113d371ae8655449", x"8a4aeb479aaf066b", x"6873d9414ce6aa03", x"afd9c24b3d0e749e", x"04f7a56b86a51f15", x"e8d5e03b7259ee8c", x"f1301c4fecc09afc");
            when 24686367 => data <= (x"791334f74d412f8a", x"fd703a3210630b88", x"842b88c232278335", x"f4f84a8583d6b50d", x"791056c768c109af", x"ab7c3d2580fddb4d", x"eb5b3e7a24db65e8", x"055d4c5610424b3c");
            when 18647708 => data <= (x"fb484916b3b9ba8b", x"6966181c1b4be43a", x"7b37a4b653d83be6", x"a50668b65bd17a64", x"2c4ff019017d927c", x"584bb1adfeeee5d4", x"bf8d8c0fdc8e8c88", x"2cdf3b13bc922432");
            when 23227744 => data <= (x"5b9c8e3501cdaeb1", x"f63b87d83c752a9c", x"ca48421cc9a64f11", x"4100da870618eb9e", x"53c4fb20abe0e7ea", x"1ae7567ebb354b9a", x"2c21c36f316c61f8", x"2d370eb0e4d3ec8b");
            when 14283635 => data <= (x"be000d25a650c93f", x"bcb3a7079e992d38", x"54e7f60222e0064a", x"a724d2115b112986", x"b8c754c94f590f1f", x"07f100d2ae2b2519", x"bfa3145e482772f8", x"fd0ea10a6a949e69");
            when 458038 => data <= (x"11668f63b2f89a8f", x"625ffaf9ec3f825f", x"f58f2796c0a1210e", x"01702d464b76d0c6", x"2e8cae784cc263f5", x"e44c8f1fdf13da6b", x"befd65c4be21b599", x"1107ea2650146a32");
            when 29784066 => data <= (x"bebd0bb931376803", x"19fb4acf4c3025f3", x"2a238f1a70c46f83", x"20c42a71e771b0ef", x"463a2daaf564eb79", x"f3717d869a92ce87", x"f356133ee9d9b6a0", x"2f5f2014fdcd1e7c");
            when 13011416 => data <= (x"7f86ad99a197f1a5", x"e11fce02cc8b7952", x"720811c716ec9e24", x"21b665374fa48fb0", x"3fd0d88b312209ae", x"874989bc1ac0f68b", x"4cdebdc7bf491df8", x"7561d961d7a63e95");
            when 29074329 => data <= (x"eddad36ce46dd8ea", x"2909670c18abf507", x"8094ca9ce02875f8", x"f5096c02e3fa64db", x"21b02e7e84518fd5", x"bea2e71769bc3724", x"15812408e31f208d", x"bf6b645629030bd7");
            when 31768217 => data <= (x"5ca5d424597ec4e3", x"0859004210b9d8d6", x"a52f05ec0c44c73b", x"dda0ee6dd99917d7", x"a5cdf70bdaffead6", x"e067472ce00974c0", x"fb14663f0b4d8946", x"5a596c0c8292d139");
            when 8968889 => data <= (x"648d6165af7e571c", x"cd068ebb722992e7", x"6255287b74ee7a5e", x"fd72296fb7697ca9", x"55f49d8fd573f6a1", x"eb080cbc49ba1a2d", x"262a6c0d2a33184f", x"549c449ad79c7881");
            when 17800852 => data <= (x"489c580ef5f62f2c", x"f0b048b6d2784f93", x"fd34b2bacacda079", x"84950ce652a81bf3", x"cfebbf2b18a717a0", x"83ef6f3347470ba5", x"90a2f72585be78c7", x"f83e1a6af1816e4f");
            when 14132274 => data <= (x"2cd3aaa2d1416594", x"654d667fbdd55942", x"ccaaa9199edfa41f", x"ed87a94de701b764", x"5342873bde7c38c9", x"27815f58dd268f15", x"2e985f9665b155f6", x"324d9170d5ef18e0");
            when 4905071 => data <= (x"e94a719f8222fd87", x"02e70f3edbda47f5", x"f33a583f204ced59", x"286d869da169e0ad", x"90acfb61d46eb998", x"bcb43523de791b19", x"34b8db516a902550", x"4d19f6fc092bccf3");
            when 22088808 => data <= (x"b7a615e53ffa6d31", x"e9d0ce3adec3a768", x"fb6dafe7e6f0a3bd", x"96bd0119db354dfc", x"4170172781307e4c", x"5674780907ddfed7", x"616ef7c4cb7caee7", x"de4390c5d0bd9f97");
            when 7475537 => data <= (x"f7f41760f14a10e7", x"eaf0c3deeb0e5cf7", x"c048663ab36d92ec", x"208106d9cf2d750d", x"acad57dc2b44110c", x"22009881fa6b0e57", x"fb1ed0ab96452f1e", x"f973b1525a407c0b");
            when 195206 => data <= (x"ecfe9d6e3e6d4951", x"79127917435a5ecd", x"37c8b81e97e2555c", x"79fccad4a6c1df7e", x"b5842825af271231", x"7269716ad3d059d9", x"bd05dca672ea68fa", x"de50513479ec9f0c");
            when 12578741 => data <= (x"322484d10f6fba1c", x"37b441296b774879", x"a03e03903701bd1e", x"e391fefddf6d30d5", x"6382ff63f077b972", x"7303cbce960ffe18", x"b27b5f872078af41", x"a65335a01d4ccee3");
            when 874071 => data <= (x"7bd09c7b212863b3", x"af9cb695ba9ee2fe", x"929c1d61563502d1", x"1cd903ffd544729b", x"594c00c5e739a7a8", x"6b95b50fd23d22a9", x"718ee0b36da9baf6", x"17f57d20d8810402");
            when 7774929 => data <= (x"0f650fb3118c0001", x"7ba95dafa8f4d3b4", x"502c7dcd89f5c9ea", x"3d0528ad0f49edc5", x"01fbf7953e2cdbea", x"bac40f409930a10d", x"1c8abedab6005161", x"88df595b374484c7");
            when 18339135 => data <= (x"9e81c6fcc33eee4e", x"6f089397f5a1a6a6", x"57f35386b97425db", x"3883db25508510e1", x"0f9fb5eb5601927f", x"958e509bd5d408b6", x"0d76fd71b34dd6e9", x"19f1773be4d6e91d");
            when 6493295 => data <= (x"8a6c9ed892d783e4", x"57777a7888745f14", x"09c0575f92bf5078", x"19ce2136c67252ba", x"e47464106dadafaa", x"8aaea3fbe161447d", x"28181311b19d891d", x"7126926d260cdea1");
            when 1545255 => data <= (x"884a22387126c53a", x"853484ac3b4f3e6f", x"3a022158b61dda12", x"11aa09209e5f903c", x"45a6ade59e855273", x"6210fc42d8b9e2b7", x"d270164a5978cb09", x"9d6d5107f3b96a20");
            when 13762283 => data <= (x"e1677e13a25a8f41", x"1cdedaa1fad56029", x"0a3149905ff51e47", x"44e9f9376abcc6f2", x"e5bf8980178ead47", x"34c3c9ddb378f4d7", x"4231054d77ea980b", x"684a4148fb39b9aa");
            when 13308566 => data <= (x"2a92fdf8c2155258", x"82b6557daa36398f", x"853bee8b401e414e", x"7cf6b20afd97b126", x"0959d86b4283b2fc", x"08b93e38e05eaa8d", x"7300bc7d8b3f1501", x"757a9cc9951b6bf7");
            when 33202881 => data <= (x"515141510c43e1e2", x"898944c477e2afa1", x"e62bbfc7f2917bb6", x"4ef6ae5e1cca253e", x"6a23577ffc69bac2", x"a4c07edc4cbad25e", x"96ed2b0015385782", x"e3da7ed963efdd08");
            when 21337713 => data <= (x"3f3e630b6a340496", x"be4a39f3305f5179", x"d6f292ae5b8bf9cf", x"d0ce5d88841a0cfa", x"d3014df3bfbb1dda", x"72993c9202633c1b", x"e27d251d257eae1b", x"dae853cd89791da2");
            when 1830864 => data <= (x"46ee21962d12a06a", x"4402d416965d4e4a", x"ca1c172860b1fbdf", x"0ff69763c3d123ac", x"4a13d226fc6ad240", x"acdc100b91c78761", x"902dfed725436c1c", x"2ef9c6a292d0df38");
            when 20517233 => data <= (x"02ebfa7f7f22c9f4", x"633d3b3510fe86ff", x"a891ff988d2716bb", x"5b126750e96d8e33", x"98e28406137792c8", x"751096091d4c91db", x"ba35893eb9a36f4c", x"521507d6648b01b9");
            when 19228580 => data <= (x"a975576d3b9734bd", x"beea45a84f7fc097", x"1aa4a9dd5d250f5d", x"13ed95423d4281f5", x"98ac4008be519885", x"2b4c507855b23aed", x"6cfbaeefdc7a33c1", x"1c5f43626d4cba61");
            when 22674083 => data <= (x"4b7f88c2c82ae191", x"30053f1dd7edfaec", x"994a779788ece6b6", x"098d084e758e83e6", x"229cba4f718429b4", x"3dcffd35e5540c67", x"89848094fd9aef6b", x"983bf93f1f9b0fe3");
            when 18549709 => data <= (x"77a88961e7ef99ff", x"47c8265a91cb4ae8", x"3e7d3300479b676f", x"0366a56383affddb", x"e89d0b8c2d6470b0", x"5c57f029465b9c1f", x"74b3e3040d3516fd", x"ebab32ec6e24952f");
            when 22125448 => data <= (x"d8996ab92aeb5060", x"f72155f4f2c0a23f", x"ee57b1d160c43bf9", x"512f4d90147be209", x"aa76a18f94fb949b", x"45a68fa110256e39", x"b4dbca60ad9effa5", x"00bf6bcdf95fd294");
            when 27342535 => data <= (x"8a00905e9697571e", x"729c066745563e75", x"012d8fddb7edf920", x"2233fcec55be6230", x"574b2aae8d568eac", x"a79f362aad6d9740", x"c8616512b5ed52f2", x"24fd4f2eb87fb872");
            when 17655898 => data <= (x"d1d45d984be92e5c", x"51642e12a3f85658", x"4489b0906ed742c6", x"9b24399cb10e4264", x"aa3b9919394609fb", x"c7fb75b1069d799c", x"b07e036b12357793", x"96a42b2875846a81");
            when 14792444 => data <= (x"d1f2cbb05e9e7a13", x"54a73ba2bbb5f767", x"354fd3df564d25ee", x"d1b9ebba4a3a833f", x"2dac7f732681a2c2", x"b22efe517b1795fd", x"67d8bf68b8811eb4", x"76ae85c7fd59295d");
            when 15211065 => data <= (x"ee28ff5db3913cd5", x"aba8243a3051b5d7", x"6080710ab006dba5", x"1499b6598d44be2c", x"f22ad8775dd94fd3", x"ffa4ecfbfcfd8f6b", x"a658ec159ea051ea", x"fb36a7e68c4c25a5");
            when 19389845 => data <= (x"b7636b0f8fe51ec2", x"b8922ec84cb9236e", x"8d583dcd6ca92787", x"feb1649842a86d87", x"055c3e469b4808d3", x"09e73e310468d943", x"470c297352666ffe", x"a90122948dd5b235");
            when 23238976 => data <= (x"85890714d3d0e1df", x"ebafbef5dcbcce9a", x"5a9c15a63b2561d4", x"2545d7447cb35e0e", x"8829ae87c36a7b58", x"2b782bf1dc35ebd2", x"eba35bca62e1949b", x"54aefc276aad3ad9");
            when 11421585 => data <= (x"f44ccc15f6938179", x"e6b6bf13eb79a4c3", x"8d8be81c5e599b77", x"b4a5c706680bdcd8", x"1f50481414be4b2d", x"9efe870d20eaab4f", x"47a097e473719151", x"711528d790f22b33");
            when 1376635 => data <= (x"36697f5fb0524cb7", x"c8f4abaa92320e93", x"72e5a433a5d15000", x"a3d8db26a433b5f0", x"28f87985862cf9dd", x"5373407d16db7ca4", x"f8eacac13363a5a7", x"2b178904a2dd4db5");
            when 22404444 => data <= (x"6053c08446db6d08", x"50bec8068c85d2bb", x"06a144f5069325b9", x"348ce34964f8f89a", x"b1718f028da4e28f", x"a42e41539e2bb09b", x"105611f1ebf53bb4", x"2d9ece6eae6f9ddc");
            when 15370562 => data <= (x"ca1f3bc69792b8b7", x"04f07d26a61148a9", x"d700b9df4996b645", x"89c4aab77296c8e1", x"eb38021453304d51", x"6a678e505637f02c", x"978ead049123ae2a", x"1b1358623b99ee2c");
            when 502846 => data <= (x"a339a9f527728a4c", x"0bbc036e4c18523e", x"a5a2f9ffc05a6d72", x"41735986d84e6969", x"259cb50391154511", x"25e6edfd601da5e3", x"8a9b76565351fe3d", x"5155d07d3e45822f");
            when 23560202 => data <= (x"4e51ae0b8e4f4060", x"3c1c4a140d1818f5", x"59041ff388c7c1e4", x"9cae35958f1999e6", x"dfc1a733af926e60", x"0f1777ae188a93d8", x"f0850e19d4c7a5a3", x"ad7c9a6641c422b3");
            when 25976861 => data <= (x"9082e35e825012e7", x"2364967cb2f0d79f", x"17595e03ce2b5512", x"67298442b9fc23b3", x"4711c65e8a9abed3", x"6c86889ff19dc727", x"4004d043cd80cd12", x"530a941e5ebc6fb5");
            when 21514912 => data <= (x"d32833e00380ee1e", x"b103d8c079201fd6", x"80543fafc29c2c60", x"58128150a9edbd74", x"7b8c0cc287a51e92", x"7bdf8dd70eed6854", x"eefac4f6ea7156c2", x"a232170824903745");
            when 28477849 => data <= (x"cded050121f214b2", x"e36444b2be199ee5", x"4cf811d843a3ee8c", x"33b353ecadc9002c", x"f952c5cbbd59f117", x"8f6748ba36437d02", x"3e459ab36b57d295", x"278cb711c519a0b6");
            when 33555656 => data <= (x"d20b279e56609b9e", x"cc1d355b1beddc3b", x"156e2427883be759", x"1a3c03e3f198a54b", x"1d74f8dbd9ff7848", x"8bea5bdf3b2ddec7", x"fb799bc4809ee7ac", x"1eea3b63b9ec4854");
            when 25113096 => data <= (x"974685b126b5d240", x"cb1b0d3b62011ac3", x"9758336f42cfc94e", x"53021bce72bf8261", x"b3e5675f91bddc51", x"a1bf91c72517a156", x"4dc8c724dd920964", x"0bf1cd212e5b7c3c");
            when 10859981 => data <= (x"19010575504a3a6f", x"22bc48361cc41e5e", x"c1347774f478ce03", x"0bc9cfdce95110ec", x"5178559e68343914", x"76c72b41fb0c3afd", x"0443baf75d99aa47", x"afab96257012bbfe");
            when 7877756 => data <= (x"0f7126b296d42b40", x"57240b7db610b150", x"e0991d13e8ddf8f2", x"3c576e53961ec175", x"abfd0a339ada3cf1", x"edc2d92b14745915", x"d02ce549b562c8c3", x"d64522e4551f6ee3");
            when 30455976 => data <= (x"4a970417756f4c9b", x"db6a646df1092df3", x"6cecbe7f92b50106", x"136ccf530b2dbdf3", x"206c65dd1e629c3d", x"2bc97fc7413bf2bc", x"e3eb2ad3c3b242c6", x"d92068f32fbdc1b0");
            when 1223255 => data <= (x"eb9ee674de56f6c0", x"3fb2ccd52002a7ec", x"3969c3571dafa9f5", x"60dd2f613297eb62", x"849bb41a89b45162", x"64cf487ba6c3c538", x"78a54fdd99ba5797", x"8dc950ca3ba610a6");
            when 16671611 => data <= (x"e9ddc561484195b7", x"cc0bcd7161b5813a", x"37559ee238ead89a", x"f05f80e2f8efb663", x"60cfcb92b7f24f4e", x"8f7b2af40aa45c51", x"26b3a700e24d5634", x"f17a44072a546bc4");
            when 32845386 => data <= (x"378156b8c8be2174", x"9b9aac2f7c9a3442", x"04d363e19206f6a0", x"d4e9e857fd563dab", x"af138e231abac5b2", x"64b7b1bc475ac16e", x"9503a1ddd54225fe", x"38f61abd10e62481");
            when 20813111 => data <= (x"3ac783e9fafeb58f", x"1c8affdd8d2efd5b", x"c7e4edf458a2ce4f", x"8e19d69103b14b78", x"9b884917a3713d0b", x"76c2939d431bc160", x"64e13adae2dd6dc3", x"ca3fe2ee46c07b8f");
            when 17350763 => data <= (x"42bbcd40ab89c3cd", x"d70e51221f6ed987", x"ec66fce4ffc4073e", x"bf62dc07c2240d51", x"c05b18064fc9eb8b", x"5e1285ca9f74ae13", x"c3bbba56ba896d0b", x"c23bd1db48792248");
            when 23809504 => data <= (x"2ac55185189c22f8", x"72a5b086dde5ef4f", x"f8daf76f3573805b", x"cdeb4744fd110421", x"6abe6b3fec7cbd49", x"b5eb627d6af07abc", x"9dabdcdf89e9a76c", x"b0a0e4a49e04c51b");
            when 22117844 => data <= (x"712affefd90e87a6", x"9cbc619b7a9b299b", x"e06b842f5032e914", x"67f97b62e57072d9", x"18b994d83ba2db46", x"c1ddf11fa2ba15d7", x"46948d27c67acabf", x"471eedccb3f651a6");
            when 709973 => data <= (x"2fd2e81c3d4f4c9d", x"c326593e474614dc", x"ccc13eba285f6d9e", x"7068e0e40471f09b", x"136f691a1037df98", x"ebf064fccdf48765", x"d186677d6e6b34cf", x"a093abb3790c4cfd");
            when 14122498 => data <= (x"67900e4424377a76", x"63cde57a8a4ec627", x"3782434240183166", x"167deebc2a54ebc1", x"e827e3b957c88186", x"63a75817058ef41f", x"5201a2b00b55bb1a", x"782a9555f5660de5");
            when 8644331 => data <= (x"c46cb0b86374f4c2", x"6f063b251f143518", x"e10434686d61d0d8", x"84b1db65443cf7b3", x"977fcde4a98d735b", x"1234d1abc3fc187d", x"2155b6675ef4cd25", x"fc71a41306b59007");
            when 2341098 => data <= (x"cdcca0f7c0f1c94a", x"68bc601982ff9aad", x"b02873aa64267b14", x"83edfe707a78baf9", x"2edafb2f62ac2172", x"d671e8af885f950f", x"60ab6d3d7092d8e7", x"fcfdfa2f24bf0f47");
            when 32979373 => data <= (x"ea103ae14e0945c0", x"87e0d09485892ce9", x"3fc5e3a718c451c3", x"306df06fa5047d80", x"ba5a8f7206ebcbb0", x"d90943aaf01c77fc", x"956f23132da01f41", x"199503c8a8537a1f");
            when 399319 => data <= (x"345b6cde980cea57", x"cc359ee9438cd408", x"1dc65f4df16dffc5", x"32fd88c58ef9182c", x"baabfc86de1fff66", x"865d424b8d82ae01", x"3f274a9328395a2d", x"547dc85a33d8c971");
            when 13627730 => data <= (x"f0c3430d6a7fc9b9", x"056290976b279bfb", x"b3b46cb2f0f03c3b", x"2a3918025d0dbaf2", x"e9e5f84f8c69a508", x"0a4acb640e25e91b", x"f095370cfffe7ba9", x"eeeee7b4ba75873c");
            when 18697547 => data <= (x"602b880d74b3d031", x"b4fa95272b5e19b9", x"5c9fa6f11cd7334e", x"b96ac047ed74d77d", x"a2f6a52450d3b1d0", x"682f1c4cd7dd3d55", x"c179b952d91dd80b", x"602de357668b47ac");
            when 32072920 => data <= (x"85c9d40e2a01f0be", x"df4da254fd41b5d6", x"f3d3f1ad144e540d", x"153831d95315c870", x"6d5fbbf2b001373c", x"7829bca5b8fd5095", x"217b6b1f7e09749c", x"30f6e079535d0786");
            when 6525732 => data <= (x"4af27f76d769898b", x"22fd91bcc6a5f54d", x"f3b0737ef973edae", x"b2e33577da8fc539", x"808a716f0e894e38", x"ac8bf038858510b5", x"eb55214247c2fd1f", x"2519f4e69f6a4dd0");
            when 11958268 => data <= (x"ea85907595b580a3", x"e256b0d2fde67c62", x"07db5d73a7154584", x"869328bd66e53271", x"fe20a2f51f46b90a", x"f8729cc4b108345c", x"b1ee39b77536fc82", x"ef3370b2f6e14a8c");
            when 26677975 => data <= (x"53c13e7eef05f6f2", x"720e009a845edc9f", x"fc31a7479231541c", x"bf71aafd28538cc7", x"bb2c731c0d879adb", x"d1636296ac9097ab", x"0096e6e786b97eef", x"6f7e97efe403c141");
            when 28736193 => data <= (x"60adf9769b2de9d7", x"e900b9b5f1f6d19f", x"57554495703e87c4", x"0931d5848dcec2d7", x"a2c83bbbb627b4f8", x"03538a3715bb77ef", x"8865107ca527c8b8", x"1b8ea5a8784e1f01");
            when 957371 => data <= (x"bc2fc6bf34058e2f", x"96e728a7186e5d3d", x"3a414862438e93db", x"5566bb41398b62a9", x"b5ab46fe19952e27", x"51a60f3c6b22d720", x"39dc0aaf65bb8f00", x"554fabc3cbd08f9f");
            when 17588077 => data <= (x"4343abe30a6ae913", x"3010506bb84364dd", x"9bc614ef7c2777e9", x"9e9682d263046e7b", x"f8f68a36c259b17f", x"2b9afc9fb357e505", x"c61e9eb59e50dabb", x"1f9122947cf7a358");
            when 33195277 => data <= (x"720c123e56dbe074", x"0cda34e70cf54127", x"77c21138ce6acf60", x"4ae325acae51ed90", x"4ae3167cf52a0a7d", x"1b0d087d0e7fe75a", x"2b9ddf3b6c79ba60", x"6e055ec33a30cdb5");
            when 28639865 => data <= (x"cbc085d2dc81ea71", x"470edcfedffa3e37", x"da8e4b042d59f464", x"2a829a8acea54f73", x"8f8bb20905506968", x"321da0d0eddc30ce", x"924bd82fd38ee1d7", x"225814b321b4cb6b");
            when 19050724 => data <= (x"69332e5dd87d34a5", x"58737a8e5231adc1", x"12e1cdcc2af01c6c", x"c8bd8e865d9b0e04", x"8f66c7ae2fd0e220", x"aa747e4e33d10ffa", x"0a7d410cbecb0f22", x"693ffe5afb9c0508");
            when 32149750 => data <= (x"59c305b836a769fa", x"d18d7f02ff777909", x"4318a08ddb8a1461", x"87109139b3164ad2", x"dd58324eaec2e27b", x"f7ea5a03cba6eeaa", x"8eab06d29f8eaf21", x"2fbd6a8a2363182f");
            when 3117979 => data <= (x"c404151a2006dae4", x"5c100736b339b1ac", x"d457a4e84a557417", x"f9504ade7f1b6dfe", x"27fe074c9e4f60b0", x"14f73c236bd8bfbf", x"b3ae106cdc825201", x"6e17365e702d17d0");
            when 22748851 => data <= (x"a0aa835b2b1af049", x"899631ae37161a42", x"a74e8b93636278a3", x"1a30859ac6911392", x"bee7ddc50ac70e24", x"87dbfc23a0f00560", x"d508305d83cbf548", x"bd724d188973a9f3");
            when 6426221 => data <= (x"67dbb817d7dc8014", x"a6a841e017e69564", x"1f0a91dd035b8893", x"cc85bcf8dd9c7e9e", x"b7308d3deb64cba0", x"78bdbeba40a35a82", x"3011630b360c3805", x"3c29efac57ea58b0");
            when 19399321 => data <= (x"9c3bb85e966273f6", x"a3f20edad95827e5", x"0fc3dfddc5965897", x"f8a89d2dc0f3ce74", x"41c97ff2331a5754", x"76c5ae261a0cfd84", x"bf7c0ce3342fbd5c", x"590922615e3f1392");
            when 16569743 => data <= (x"d62a7e13c1b5d23a", x"fc33a94e1ac5880b", x"c95a307cb1baf5fd", x"55f88771a5f9bec8", x"327d70c3b100db13", x"fce4aa49f52fa1fe", x"22293d68917cacd2", x"8bda4ca7a8229e5b");
            when 6582414 => data <= (x"6de2f0aaefd231e9", x"618a54d0abcd07cf", x"167f5de31224737c", x"fce1e573cf7f5297", x"1cacfaad144c1eb6", x"a7cf924345d55dd7", x"9a8a7d9a983f6b45", x"3e58faa82e60b841");
            when 9043586 => data <= (x"480f7794bf0305fa", x"52625cbae98d9c4e", x"8b17b5c2a084e5a5", x"d8bfab694df30144", x"4eea8645c564b2b2", x"847a39184647c9b7", x"0fcaf5c6f369dabf", x"14ae6d3aa4b4e995");
            when 18276979 => data <= (x"279febbf9b19cc12", x"77d4ed681a26e316", x"f5f5b85632a7abd8", x"ec5ed277e0172284", x"967b2b476c3c6817", x"238b2e062605d53f", x"a050770e3b0d8a36", x"c9f87be38165302b");
            when 29219144 => data <= (x"960ee57367c40096", x"efb2984f3024892e", x"14dcce2ee48a3811", x"0d9280b1c66be059", x"0089c832a4b416b3", x"60e3d639a1aaf7df", x"7ebfe1aee1a4f5a8", x"77132295416c15f1");
            when 10081091 => data <= (x"cc11e5d7bbfdb49c", x"51f87d11fbf160ff", x"27af2f96b7dc44df", x"610d959ef7255c33", x"a80ecda0808372a7", x"1ff49c8f7229be2d", x"06a88785bd2aaa5e", x"31e6fa2368226b4c");
            when 28504587 => data <= (x"9333b1ed9ec3e6b4", x"384fcf9667161472", x"a03c224b136b0de0", x"419416ab9b77d7d2", x"2cf0fac01381745c", x"3ac821f3b0dd5570", x"80b44f553e9097d3", x"cac202802540bf2d");
            when 9762885 => data <= (x"d4555cad2045107e", x"ab969814fac1e3de", x"65281ee11b09bbfb", x"1299d55ff313650e", x"14954a336be4affd", x"de468a672bf41429", x"2204b5e7e4b07e7b", x"f8232c635d4c3bcc");
            when 11531608 => data <= (x"b7c8c107c6aabe25", x"43d3f2c5d1a8c5ed", x"e93837605f3fdc6f", x"fe50d7938008ce87", x"f454a269bd30cee9", x"7d3c83191ae228e1", x"588ad261190a1b98", x"e4964774199b3565");
            when 10385062 => data <= (x"dac30fd804cea47b", x"085a04d1fd4a830b", x"c42544bc7c6883bc", x"5469a7c040992a75", x"33d97b8d98d3e0f1", x"326b07a66eaa4024", x"3205cb7edce8c5f9", x"fb7ad7881128460a");
            when 17342760 => data <= (x"34d50f914f82f2a7", x"f7739b9ba65e1e2a", x"5cdc7794277d1cf8", x"a3366e718595e8f7", x"51742f177ff8d6e9", x"c3e07230e7121f19", x"daac2bcde91d2620", x"aa3cbd26f3c663b2");
            when 28367614 => data <= (x"ede651e586393e56", x"ed76dffdd4b34946", x"068d1d0c8dd186c4", x"7e412d9f1d9a53e9", x"6a6c4728cc129c84", x"5ced8d43869ba6cc", x"7b107b387e1fb24f", x"72dabc73f89b925f");
            when 13258337 => data <= (x"f480a083898df264", x"2f9f448bad0fb8ca", x"20dbf569e559ec1a", x"4f1affcd9d320ca4", x"71f1b62b93684863", x"99a026af377c6516", x"3131be8f4d6a07af", x"308cbdafd9d03fc8");
            when 25772667 => data <= (x"1d9c33633753680a", x"8b72078d66b056b5", x"c7558366fc3c4ffd", x"faf709adfcf4f50f", x"814ddd997aa58bb8", x"04c8a38c8fa0bf05", x"8502c754923159d2", x"69b849148e197154");
            when 19072305 => data <= (x"c32980336defd3fa", x"9e9daf88ce86f358", x"764c32c38db9a172", x"25835d185bcf49f9", x"1262020efa91fa8a", x"01f1db8ffda75445", x"5b045e9041f03b7b", x"fb68705929dd5f17");
            when 30294952 => data <= (x"55cf93583bc91ee7", x"9b21284b24cc102f", x"700741ac90a06c1f", x"d8bb8ce9ed0fdcde", x"76d5f55262ef6d4d", x"f6b4e6710c7835f7", x"ed5746e3357befb8", x"43165c942f9ee38b");
            when 31422587 => data <= (x"430a2b6b671b0e1c", x"67d2a0fd6b2fdb83", x"5f086ea9d3f6b76c", x"fe7c644795ff322b", x"344b5126c6e6a15a", x"55f747917edc11a3", x"9da9574cdd416b29", x"4a1ecd9e92c8cde2");
            when 14590733 => data <= (x"7462fec24c23b3c3", x"51170591314717f5", x"e2c4634a455d466a", x"ed83fc4d8a014e10", x"5ccdcfbfafa82fd2", x"273df9f92cdd1dd6", x"06b0868e7fc0e6eb", x"53a52be3aedac9f1");
            when 20326696 => data <= (x"72a324bbdd8f2aa7", x"f8e7ec01ffc3903e", x"8e9feb3b75f554b1", x"25d952dab2e37389", x"101e81c48b76ef85", x"eac3ed5bfb1dd21d", x"827f34fd60b780cf", x"c24b175d7957972d");
            when 12349940 => data <= (x"483713fd30fbf57c", x"9bb283dd9f43b22f", x"43addfa54830482b", x"537d3bb3e8eeac13", x"c58056227de4b963", x"7bdb2f50d183aa66", x"8cb39f488a3b1549", x"0fe43791063c82cf");
            when 26563656 => data <= (x"e133cdca9b399bb3", x"120cf377e7f6014b", x"f08d8635fda5fe75", x"cf0d9490040d2929", x"32a514f0757e6643", x"6192e171f65acd9a", x"a0028f4d6e3e8bd7", x"94bbbdeeaa9b2aa1");
            when 18429144 => data <= (x"f2bd040dad9435da", x"41c9cce067d32df9", x"7e499d2802c56166", x"8126ed93d3dabd6f", x"760486e4cc30f249", x"cf1c05d1b7826d01", x"6ea55e2f4494fb5a", x"37b44f766f82361b");
            when 25228141 => data <= (x"c64ad94922b93f5a", x"56d764edc5da0e2a", x"d4a6867900156874", x"7ea05fca4c22be74", x"f232cc4939e4bd54", x"bcd440fce3a6dbb4", x"10d58a81df68059f", x"899a0755eea9d9ec");
            when 17601968 => data <= (x"008cf79ff1d94f51", x"a1e0ca6a80aab6c5", x"51866a0d1190d74a", x"182b37e4b59f29cc", x"0aeda568fcc6d697", x"8ab1c9cb23630f58", x"1b990842034bfa11", x"1b13964e960c75de");
            when 23181221 => data <= (x"8de1ceb896611337", x"cd59cf5846bef710", x"61e3c74b628bfd42", x"489ac14e55dcdc33", x"026f17414aef2f94", x"3d6486df22602714", x"dfd4b569f934a55a", x"80814b08bafc6427");
            when 18217625 => data <= (x"2d525c6e653bb994", x"95ea81c9e882fcb9", x"6a73749408f0aa48", x"f1be9d3315b1dcc3", x"d968fe22448116ab", x"c6c88f7055be1851", x"fecb41793147f4fe", x"f0b60882af4faa1d");
            when 9666098 => data <= (x"54d6a5916d614b91", x"08efa5bac44e6811", x"3743bc6bc03585bb", x"84426b72f1a5d0b7", x"419f000e491ac012", x"17828a6b3bfc802a", x"0affca604eab15f4", x"29d01e9f4b7ed0d4");
            when 19192175 => data <= (x"cdd0e92f7e282b14", x"48a1cb5accbebd7a", x"df9e8cc6ffd1e270", x"710afab8f3ecd55e", x"24cf6bd15641ddc9", x"a41ac719022ca6dd", x"09f64bfdb6705b6d", x"8e08406673666183");
            when 22849575 => data <= (x"cbc049a09b845472", x"3b0838adb5ffa259", x"ec62e6f8d83a175b", x"bf999dcc5a3657f6", x"96118efb88cc9240", x"8859bb82113c33c3", x"faddf4d816eacb95", x"e7afbb2b5bb9111e");
            when 27132900 => data <= (x"51f190157c32c13a", x"d93bffd650d6dbef", x"8f34f3cc138328fb", x"290c250f43b5587d", x"309cbfcfb6c3050d", x"4142344a7ba2ec76", x"07c9a58602a2ce53", x"c3b2fd2338c8b9db");
            when 9841214 => data <= (x"35a4a4447f0522f3", x"2417fba90060501b", x"bc009935b6d9ada6", x"c878585107e5f239", x"b28dbc1a9d4320cc", x"96e054562445524c", x"c9fce404c6f4eaed", x"77d1fdf8b2f1477b");
            when 30429605 => data <= (x"a09c418a065ec781", x"752f3b9905157a2e", x"53fbb31678c0b926", x"2496c8c79ae95ccd", x"0e45e79e85711e1f", x"58eb948550db4eb8", x"e29efc3ae5f4acc7", x"b0c0b709c1acd13d");
            when 21779822 => data <= (x"896f8262db0d476c", x"e59b505ff46d761f", x"1f3ae3a9c5ebd4f4", x"738cbe018f380709", x"36847050f57315f6", x"1325449b30be5a93", x"a5722c85de86f807", x"4b5f8bdb049ec62e");
            when 20081898 => data <= (x"1b737d0e9a50a79f", x"de814058354847ab", x"b5ecaf829efca34a", x"82e7102320358634", x"ac8d702aeb755bd3", x"b98eb97d3a5c6ec1", x"c01671519e4f5311", x"5ac760e503d19378");
            when 9505546 => data <= (x"8b0382450d662617", x"a42fcd2826f95157", x"1f17cdead41ee362", x"4124d3e055a940bd", x"21bb0584f5abf2c9", x"a12df91f050b099e", x"09e0ad4651c10ceb", x"083923c5f295aa14");
            when 11453163 => data <= (x"0cfec22df68e7648", x"120e5f0e15f1ab30", x"4553d41badd3b1a9", x"2a57e66acb348507", x"ed31bb346cd1ca34", x"c0676886111e759a", x"c529b81ef86cb294", x"4aa0bc9286f63634");
            when 4624912 => data <= (x"cbf1f41615ff2b88", x"32edecdc6e728814", x"8a89df2ba17d3809", x"32613ff233eeda4a", x"1051cf8e43874741", x"ddb20d6cc00a9274", x"fbf31ac51b0c2e70", x"87b69e9692733e38");
            when 4971328 => data <= (x"f917e192ed7f2d66", x"216348d95cc097ec", x"3a4e425f0a53b0a4", x"512450d12ebcf177", x"356568af8e08d662", x"e43500d24c531a8e", x"cad6564f308ab464", x"d295a1097ff29f18");
            when 18913052 => data <= (x"e9e8edce927b11ed", x"5ca84878637c3ba6", x"36e208aa5e88ba00", x"f8e249310eb2c5aa", x"d433854fc2c95295", x"3471bcf6c4824e8d", x"d8e70e7027791258", x"cb60cde16851ddb9");
            when 233294 => data <= (x"bb35ae811b147575", x"9fb3b34c9e58d8e8", x"2b71c62d9ec233a8", x"3ac8d5809b6f32dc", x"b675cf7c9d4d21bf", x"42c1673f68a88565", x"183c0d41403703cb", x"3355cd9083621879");
            when 29608453 => data <= (x"1364bfab4c5aa871", x"00cfb77d51dac7e7", x"0f1e06c65210a1ae", x"99ef32de2b88af07", x"c04d456fc0c999d2", x"29d6c67eb2cf1544", x"4082d5425e4bea4e", x"49a1eff20077b2ce");
            when 6206227 => data <= (x"5720ab291bd4536c", x"fea94708b9a90e9f", x"8bf62b3c3a787313", x"8bd5f0a992079f41", x"d7f9e233bba0d2d7", x"636a555d996cdbbe", x"24c76e77ab229e85", x"9feb7fb073816755");
            when 21111576 => data <= (x"c9cef78108d6dbdd", x"711a08e05336a28e", x"d81be21bbc3893f1", x"d95d57552a7acb81", x"d755f316a9d178a2", x"0f3de57aadc36340", x"4242caba6c79ce6b", x"8135b959f99e4b7a");
            when 31325888 => data <= (x"968c6ba11c4d0b32", x"53a022633adb3e13", x"4463a865b69ef91b", x"0d0b2f39365aa71b", x"ccb8b245db780ae5", x"09b3b835b2bf622d", x"57abdcb59a124779", x"fc8d2be94c1566d0");
            when 20005447 => data <= (x"73175304fab60a0a", x"2bb500a02204d26c", x"ef3e02eafd40bf95", x"d84abcbcd9a8b876", x"1185acf85320b053", x"1c07a524b94b6190", x"de359a8bf53c1bca", x"f0537b5d83279a8d");
            when 5000477 => data <= (x"c12bcfde0ce7606c", x"f1c43e43cb7caeca", x"77522cb4ff03049d", x"2b789dc832ccddad", x"3bc64be8815f3b8f", x"382b20a77102ddee", x"75b3bf32195cd298", x"cd859a1c5fb332ca");
            when 2330006 => data <= (x"95e8ebbd59c43195", x"9cf043c41e8ab44e", x"874110542aa6e94f", x"ffee83d4abc7e982", x"cc3b14ff5ea7c375", x"124a727811ebc784", x"8d32e6c26eb38975", x"95b6b6dadcce3070");
            when 17834081 => data <= (x"008dfb71898806e2", x"9486e3a6fbc05c36", x"832fb73d17f36cfc", x"a3cada48c799f420", x"0b6de7b135354b57", x"84cbb348c4495435", x"0954953d0328ccb2", x"d5b98a570b62d421");
            when 10096976 => data <= (x"4be2883897f67f88", x"69d30cd41db61a52", x"a1f043ee0183afe4", x"a48e8b7cb0eb3f98", x"62bad6601e0af6db", x"ec6a321dcc3f3d25", x"76bd88de447748ae", x"f213ecc6dc9244ee");
            when 25215957 => data <= (x"21136792e83a297c", x"e8b9eedb16508c71", x"195a38e9ad9b65b5", x"2f0d5e71ca6cd764", x"798374923cec5c32", x"585bee701f32ead9", x"2782d8a7f4763416", x"24a34c7f3b820580");
            when 21645852 => data <= (x"157e4775163c8224", x"9eb71bc230364ae3", x"cd779bc9ab3358ea", x"d6bb4dfc4d1724f4", x"e4b6ae51950f754b", x"10aa1136afc132e3", x"124f74fb045726b7", x"50fa9e2d6e0a8fc4");
            when 25573484 => data <= (x"027ed53d2b943f32", x"d8d9c8b01ce4b6b6", x"4b1137aafaaced65", x"c0bfa27894eabb62", x"37f97ba84f47a8ae", x"9ab8864a09a244ff", x"e261862ded4cb1c6", x"451c4e1affa6a196");
            when 19945315 => data <= (x"0c832c139ac4bb19", x"e380c8587c179c44", x"39d4432b82bbc844", x"ea2f6084b4363ca9", x"d00524c06305127a", x"97b83c72d691ab5b", x"9ca74f5f35549f93", x"231a87a7e4e0b46f");
            when 4802645 => data <= (x"a40bcb916b85aa7a", x"688ee031f19007a7", x"f6b827f4b1d65d84", x"72d3894853ccc2a9", x"71fe2b656cfa63b8", x"ff13f5efcfa6b06e", x"541aaf8f763f4508", x"57f44881d3321207");
            when 30379959 => data <= (x"b2818eabf0ff2133", x"9b60ac479128d963", x"ec62c86045d68afb", x"4a3c799ce1b07d27", x"d17ec1420c54606b", x"b531bdf8021d4d51", x"d44478f95e8b5b1f", x"7e272f7422e23b53");
            when 8946509 => data <= (x"6fd2666666bb2526", x"41005ad6573ce498", x"b27c6bae1c7c85f9", x"f4b3bf3e237fb4aa", x"e64de645b5e149e3", x"f2b4bebb59faeef6", x"c98a80d5f0b7afd7", x"13fa6d09121c7d9c");
            when 30143755 => data <= (x"60bde2566d1e6060", x"c8d62f6dc9bd20ee", x"19352cb7beff5fd9", x"6f0648f1ff4bac65", x"d28954b11c462b29", x"c0ce1515132efb9b", x"99b5f5e11b8dad19", x"03c85a160649bf63");
            when 13651220 => data <= (x"9ac5e7fc95326297", x"ecfa7a38f317823b", x"fe19e2d71448041e", x"757012456bd94290", x"25836c7d759bf4fd", x"c3ed7b021ac756ef", x"a17aaeae0259050e", x"e1edff8e882ad0c3");
            when 1451206 => data <= (x"4ad2ca184f3ff3d2", x"854290779d3b193b", x"d13461790bf39af1", x"06609996a38b7c9a", x"467178fc1a3272e8", x"89bd7e1bda6c30ff", x"b7281b241c4f73ae", x"5bda5384a3acf755");
            when 16560773 => data <= (x"d0a206431e6c4330", x"909903c56675a3ab", x"ebcd7bb12b52bfe4", x"5102577848043426", x"cb81933a013504fd", x"980424c827078b1f", x"29b9ffbb4fd9c4d2", x"8b586c57e1f4bc6a");
            when 14426860 => data <= (x"bcd48676eb2c638c", x"2c149586e7f589cd", x"b56999003ff1ef12", x"682e9c427e26ff2c", x"e5232e1a2e7e7447", x"7f973482a0a01acb", x"8285e3452d9e8af0", x"fc4c78685f95c857");
            when 9759386 => data <= (x"a2f63c76d27b942d", x"b035c8a5efe86258", x"1526032c5c1e58e7", x"467ba29065bdaa99", x"609d44d17ec181a2", x"861016082abb14b0", x"0c618f8514b7d892", x"1bb356e11af9bb40");
            when 17155943 => data <= (x"bf7baf64fda05eea", x"76fc7bad9737a767", x"eb3d3a8a20908152", x"1c231734ebe6e2ea", x"bb5f73569b6496ef", x"f25e0b45e7af6751", x"fa3bd76bfa09fed7", x"b59a6b168aa870b8");
            when 11482685 => data <= (x"7e7e8239edcc23a8", x"f343ca5c5268fc59", x"656d946fc87609b1", x"21647624ee100be1", x"66e5c00c60d4484c", x"ad78d7877639ca24", x"0b5b17c597788bd4", x"fd542209731395a9");
            when 18256415 => data <= (x"611b642a393a4866", x"e7e68422512f0444", x"ae5363c45c0cde7c", x"79c41a13e9f62d8b", x"b7a01a8968d4acfd", x"7443e2e6a9389573", x"1aee1da20183d64d", x"3da97d37549c7ccd");
            when 17580705 => data <= (x"eb095dc444d1c66c", x"4fcd5c8ccb3acb27", x"6778fbea5dc32691", x"4cd7566dbee459c7", x"b56248bb4129f496", x"19a59c8ed20d41c4", x"9a8870c27410c961", x"ba8ce197de03d9ec");
            when 18468239 => data <= (x"e04ecb7694f8cee0", x"5d02e4ddbb813c4d", x"c1ee9ffe3d75377f", x"8bb32d688773e983", x"0af115e99b1b90ec", x"4e2d1aeadc6d8ac9", x"d2fdf78f17827fab", x"f8cf1dbcc2f23407");
            when 32053280 => data <= (x"7082aa114637cb85", x"bd4354bc0386a600", x"e14fb669ddb079bb", x"f55934a1a5d5f559", x"0c7c2934557701d4", x"4630d3d5bb9799f2", x"58f67119bce3cf3c", x"7a7b519bfddf0356");
            when 7837154 => data <= (x"60cb3713ad6b1cf8", x"b74485e7cb9744e9", x"8144b00eaeb7407e", x"d9def98c9f8ff9d5", x"42ea550c67258be5", x"c7d9205d4a2c82f1", x"35292ffcb5e59b72", x"6d35abe2d429f462");
            when 24971811 => data <= (x"89538664afecca82", x"3f176727f238765b", x"bec1752be1143d4e", x"2a8d97b1e4aa96c2", x"f2f5fb6e895a420d", x"97c2f958bb7b6b7a", x"a775cb42a33071ee", x"a53086c77631e8b6");
            when 29003853 => data <= (x"3b824c59554ff776", x"c07dc7f2eebfcd0e", x"bf0d2d951f198ba9", x"81f103ff28467313", x"eb450aa5635f8589", x"5c0dd872b6a1e4ff", x"ad7a394864ab8ccd", x"db2c041b433bb897");
            when 26682026 => data <= (x"3f1decd4d694ed94", x"d862f79dd1b9f8cc", x"a58c9409b1bd7874", x"e28dd57cb24b73d1", x"ba56b88893b49b79", x"bbe80db8c5b64196", x"166a471987b07ea9", x"cf1627ebc277ff7f");
            when 16159747 => data <= (x"ffd3f3541fac4638", x"6b63b902d695f100", x"afba8504250a24ed", x"ee7049060590afa8", x"4fe33b6282bc95f7", x"37b368c09b950d1b", x"3e90500f8ff63742", x"e86df1d48de2df5a");
            when 32818080 => data <= (x"18de481b8503e9d6", x"1aeff5c9e299d2c8", x"0d168ad5739a8384", x"7ea125271e14ce9a", x"d4fb08e3222c07b4", x"d4410bbdd4df7ab5", x"e30e2736a914dbec", x"72f96709c73b27fb");
            when 22896595 => data <= (x"53bfb1237b6e557a", x"b096f8fdb3aac6e9", x"984ff5a9b0c2c62e", x"bd2ac14811b56795", x"874b3659648f4fa9", x"fc23cee3e2ae37c8", x"4359c6f114166d1d", x"6449d04ba17aa528");
            when 32206950 => data <= (x"f0ffbb3761de7ab5", x"0f170b313e62f3d4", x"1fa56da72afa7c5c", x"011c50d15053a3a2", x"e237fc3e6cdf4492", x"3d5d68b3b77d022b", x"dbaeb0e95be5114c", x"5562aa6299c20675");
            when 14883125 => data <= (x"3a3c5ca49722dda5", x"9c859c7b7979c132", x"baefbe27d865fced", x"aa5305cb697384ff", x"0398680654eddae2", x"57627270ee24753d", x"d7c6172c24faf7f6", x"611f10c80c90cc64");
            when 3477182 => data <= (x"41160d041bc4e7f2", x"e3867dfff3c876e3", x"f7be0fed606962ab", x"74a9f2ea3e875c94", x"5f4a62b736b17bdb", x"9fda7dc50806e5ea", x"b5745d4c48440ce7", x"17f3139d127da5f5");
            when 27344132 => data <= (x"6348f49fb4e3203a", x"33f01040c3ad7eaa", x"214a01ece5846a77", x"7cdb21ee79946f30", x"f601ef84df603c29", x"a574d38737264ef4", x"5a7cfc911cf5f8e3", x"bd709c75df0b511c");
            when 30300875 => data <= (x"1288993f4efdf351", x"5950d887df6e9ec5", x"023b9fbe318dcead", x"06efe23ec96f9a52", x"4d6ff7353ccaecdd", x"e5e9ce0f0776fb62", x"e5f86dca2f4a12bb", x"14f17468527e7931");
            when 12452674 => data <= (x"570a110b33f60e8e", x"e3d6dc18b99a08e3", x"142667a3ddde8416", x"08144c0bdd8d3fb9", x"6cedb2b97b602b4b", x"eb56e7161514d75d", x"b5f7bb8ea49135e3", x"800ad23c957fe81e");
            when 23507741 => data <= (x"b4afe199e150e02c", x"e20b66dd27f2fb2a", x"4df77231147ea5ad", x"b79c932300bbb440", x"9596d14d0e6c2404", x"95725b893fd1a4ad", x"0126949818dc797d", x"379111ca61f12f14");
            when 14820089 => data <= (x"34904fd313537329", x"eb86781203ec1084", x"80ef3c3d391300e7", x"9ba0b2526879e61d", x"647c61b12b66c472", x"11334c737ca4aa59", x"dd01be6858a23bfa", x"f077a70d9574e6c4");
            when 127447 => data <= (x"9afee41938022e4e", x"7a0c6f043fbf34e8", x"55fec2f6f40e6c58", x"c51440f2fc2e4d51", x"c3e62b9eadf15f61", x"c5e9473817a76349", x"8311134432afeb92", x"357dfa65a789be9f");
            when 16936539 => data <= (x"bb3e9bb22c43f135", x"15a2cd937b363a7d", x"9cd78636367b785d", x"67da83de65bc7508", x"c6d247e4cb4b590a", x"a9d72b11dd36806e", x"8566ef31cf365ef1", x"bf6ab3171f9c6d02");
            when 11988070 => data <= (x"4d7ed44fc2b92c31", x"e17b60e1fdd1d6f6", x"e832ca4099a3b4aa", x"80878d6c62bcd763", x"f5abd1de4b0421ef", x"aa878561732273e9", x"ab459fc85819ae54", x"77bf5fa19ff0451e");
            when 23377622 => data <= (x"bdbc1c95bd157af8", x"27b62505083540ad", x"4b2ae4a229010fb8", x"b45471e038f58ea9", x"56780647ce086252", x"1a04f4ec7a80676e", x"0e044a493c9ef49d", x"0e88ed13b43bb593");
            when 28016289 => data <= (x"3473bc7b991c3c86", x"0c693c0002678ac7", x"67c1cf02e4c9a6ba", x"fd34f9b8871d4045", x"0a16bc276f757338", x"eec774af9692b717", x"f7e2c0e369e0664c", x"13c55ef5f59483ed");
            when 25230401 => data <= (x"febc083a364b276e", x"2a3beec61dd728da", x"da1658a4ad2b4682", x"877493ce6c48cb0e", x"c7a0b00fbebeb9f3", x"da5e0a99860dbfda", x"03a0c2906b7e6005", x"57d77266c7cb81ae");
            when 12507181 => data <= (x"51c0a67427e3ca44", x"55c7e2d6f6aafc85", x"f211406091e28589", x"2caf18b821f18b7a", x"d1cd9b2e49a80579", x"45b53d3d073aad4a", x"284d8d0e03f76423", x"5baaec24410cc862");
            when 5486014 => data <= (x"e046cd1f81e2e88b", x"ce4f83eeaacade71", x"286bd6e3102065ff", x"72ed38ef07e67858", x"989812fa7fff79b9", x"0bfa4f2a6c9a74cb", x"8349139b4e7d7aa2", x"4e4c89ee56f8c445");
            when 28714003 => data <= (x"5995ad145e217039", x"d285139e1841c7be", x"84c785f47b0ce1e8", x"ba5584f03ead8dd7", x"fc0ac064c96d26dc", x"ac588d36472a89e6", x"8110e1b50ab251b3", x"70b01e41b4f866c4");
            when 29533521 => data <= (x"199934536ee6436c", x"12d36e2c8cb5583d", x"d568e59348d3fdaa", x"2f28fc94906fb4ba", x"bf96602b032ed58c", x"ed687bf61685984e", x"994d20853ba3be39", x"d22af2dc01e4ca00");
            when 28761946 => data <= (x"114906c59e69da22", x"358eface0876d6ed", x"1184620f1fc00b4f", x"7f732e35ff1a50fd", x"adf4ae6b8b9726f0", x"87c881fd4226e52f", x"ccf639b40cd3d56c", x"ccbd1275c63034ff");
            when 22698921 => data <= (x"b09fe5f05f1d7140", x"08f887d53c63d8f7", x"7e6010a49dfeeea2", x"c1250a4d4a22f29d", x"7efd9b2de43d055d", x"5cd23a9072e158dd", x"f60ec6d8ed2ebac3", x"e6871ebafbfc9c05");
            when 16477527 => data <= (x"1a46daabfbfb03a0", x"e9cc80ea33dd043a", x"ad69a36c587ddc25", x"f6aa9e3d45b189dc", x"7b06bcfe0525d6d1", x"ea7d44733fa3fc18", x"c79291d5e42fb69b", x"4140d758821177b3");
            when 32440956 => data <= (x"9c352feab0ae99c4", x"1dc83645ab9aa6ef", x"346f0aabc189857c", x"0988b524884bec21", x"2c99178351be9e0e", x"6319c20ef9b56cea", x"7b47227134ba9d52", x"77d5f400d0bff719");
            when 29693728 => data <= (x"f442464f03094992", x"1cf23b4c7a8a171d", x"cac788ce0e2b25b7", x"10e014e256548715", x"9208b3ae2821f721", x"2e563fbbe1de4588", x"ddd435f81b5e267a", x"2924cf8d79245adc");
            when 6674220 => data <= (x"67d19fcf1e18ee21", x"7023fc80cdbdc6d1", x"aa5cdb41eec4e70a", x"92e451dd2de01edd", x"21b496202302551e", x"d95edba6bf0ac7b6", x"85996d849eb60a8a", x"ebe4018a6da3ba2b");
            when 17141879 => data <= (x"fcb6a4271a1a2701", x"502ef1df4d1b9130", x"8e084fa01acd2a08", x"0323977fb64ded60", x"025051e63c4e997a", x"53f65988fba71118", x"0c87e632f9f67da9", x"9c4bb688afafe233");
            when 21065156 => data <= (x"c75adc0590c250ed", x"16779450c6adf8f5", x"29c68ac082bb0f0e", x"9e17675e3f647dfc", x"d7187f2fd83c761c", x"d76a2ecc4b37063c", x"0f000a6f4c154bcd", x"f19140ca03c47035");
            when 28935811 => data <= (x"d51e8cb11f2f889e", x"2ea204df5fcea6bd", x"20e8dd9ca00e6cad", x"18819f28546d6e39", x"efd28f4827fceee2", x"d911d48393c17f1b", x"8462c01a2c2fa3c7", x"41d9a81909f9fcaa");
            when 25933694 => data <= (x"1eeccf2fb41b5905", x"9c8da7cbee685890", x"097c45c11722c770", x"c00820ccb136b650", x"06dbb58a7dd39ddd", x"ee7b02625214ae34", x"40969db44f798adb", x"4ffeba03eb67d833");
            when 22726405 => data <= (x"a9e6b8e23dfbb49e", x"42281d50ef3d972f", x"bf341624a50ec913", x"f753ae80ab13c236", x"b8e6d86e68e61298", x"8c49106a214ce373", x"1e85d0577cee9e1e", x"3f843109d94de93a");
            when 752146 => data <= (x"24a28d562bec18a0", x"b7908a21d15203b6", x"29b3dcb57bfac2fa", x"c30c5b1de72b9a2a", x"9821d5f7146feef2", x"43181146c07ac9ac", x"98182a5b46d7f872", x"094a7703ca19f5f6");
            when 30775703 => data <= (x"d5011cfd48dbb099", x"4c5e2a33687778e6", x"0a2823df7a83f811", x"540fbb1efcc659b3", x"6a32b387f0b3f64f", x"50c682ddd4af0955", x"59aa88da3616521e", x"a780d9a755d975d2");
            when 28482488 => data <= (x"18f0b3992b5ac125", x"7be205c3b01d87d7", x"6f8905a88e87bd16", x"1f778833933028a1", x"d1759d32d1482105", x"5761f1995cbeef6a", x"3f539f97d12f2a42", x"d7dfe6f1c6254536");
            when 5319114 => data <= (x"34aa2567bc3ee2e8", x"ef2d860f970acb67", x"f7afd1ad5efa1cdd", x"c9c87774f253ceca", x"68b7dace9cd5cabe", x"239a6dec8d176ffe", x"413f71a533419c3f", x"04cf6eb0d36fa7ab");
            when 21658642 => data <= (x"301dfba03d08f0eb", x"45fb948eeede5e81", x"96bcc0e8b4d9bca4", x"26be1f9f07b0d330", x"7e2e274ffcbeb463", x"84fa8923343cd7ee", x"0d6725290833b545", x"65b1a1fcc96afa36");
            when 4541693 => data <= (x"9f9bb13aae4cd816", x"0432b4aea537d2b3", x"5c1e5f7bb05f67a2", x"8bb310cc23e054a8", x"24f68c631b3bdfb8", x"5e16a57417db4940", x"871d63555dd22a4c", x"d58370a75c848beb");
            when 10055196 => data <= (x"382922fe3fc57276", x"a2c2f40a22207e51", x"9f41cb299314e7c6", x"b2c95012dcc93dce", x"d0ddabdf925b2d2f", x"fde4cf49040b93fb", x"d197c2ca0e5573f9", x"2765ac53b6fd65f4");
            when 3392596 => data <= (x"6167936b5a7fbbdd", x"ec77e1bb92600a31", x"701fc82f21e55da4", x"5a0be3cb78c300e0", x"7dec71bf9c615a03", x"606117e75c592369", x"23682e2d9e66f66e", x"fd233ec144a90399");
            when 175919 => data <= (x"e572941621eca1df", x"6f8afa6794ef841a", x"44ee4607fefd1f06", x"47ac571ae8c5117b", x"b88041de7cff5e2a", x"176cce8e3da846f2", x"05ba15186cdb4a89", x"3264162a865dc4e8");
            when 32854675 => data <= (x"a74a35a925ee7f95", x"9db76995fcf3cf1f", x"d4478165bbd7b6ed", x"064d9f5779f6b5ab", x"47f374c20bbcf46f", x"3ad1dd37619c8a78", x"984e093c724ca6d2", x"b2d9a61c9ee15cbe");
            when 6224625 => data <= (x"439ce5c487a6277a", x"4fef3fcdd615b674", x"fc120ae2349ef8e5", x"84ded26f79d81f57", x"7cd17c2311a8a612", x"5b20b42196baca6c", x"6477b2797104e4e8", x"43e74e6e038f356c");
            when 16412181 => data <= (x"231ef657c4fbb56b", x"5821ba8213e8ebbc", x"e1d7994ca95b3bdb", x"a846ef6d9cc07f5c", x"9f29926469217bdd", x"ef65c0f491382779", x"edc963cfcb943c1b", x"9408dffa067c2aea");
            when 27602764 => data <= (x"da5c3763e09e382f", x"0a2f7a621f4b776f", x"1b0151a4e88193e0", x"1a2754d09d6d28ae", x"05ac390e12d8e781", x"564566051562877d", x"b19598897191b09b", x"926d38893a0f6741");
            when 19398592 => data <= (x"7a4fa631280cf70c", x"9e799580a92266fc", x"3a248f76b32f0291", x"e6562b1eb7f1827a", x"f09012ab5ef68816", x"4c7536cd54360954", x"6d871020df62808d", x"21a50655a1d549c8");
            when 3404605 => data <= (x"9d9ffb5e6b2767d5", x"9dba118d06c7f885", x"d3a32d19dbae6778", x"08727ea36f5b21ef", x"d603b15a5e659082", x"20eba10eb168ae08", x"d326a7d7faee2cee", x"9c9333af47098975");
            when 9350614 => data <= (x"2a59ae42f5fbdb59", x"7531bed017307fe6", x"2263b198be669567", x"7dac884778ef68ff", x"3d3d7662c905b739", x"eb7de8fe507a2fed", x"f834340c5efba678", x"3b97a5d4c3914779");
            when 28561056 => data <= (x"e75671e105a6ed2e", x"87e8fa496518c3dd", x"d2ca2927881cc384", x"b3e6690a15a83887", x"f4d23a195f3a6998", x"799da3c1be5d69f5", x"27e0583ad4fe7997", x"89fa567a48c25069");
            when 12379735 => data <= (x"c8214bde24e63740", x"c51e928484483511", x"7004b73bb351de59", x"23d7439eaffbd996", x"016dafa3af691d3c", x"428edc463c05c5da", x"093d96f2f16faced", x"cdae4699c42accae");
            when 23126031 => data <= (x"ea2dcb31a29f760f", x"a428e15696b21a95", x"5e09ac70609b733c", x"2b2176fe1bffe314", x"e8a21e2c58c9fa8e", x"8f3ee573245d69f0", x"cad851a64edb5efe", x"d6b204b70fc07268");
            when 30618621 => data <= (x"5fee7a2be4032709", x"e754853169be2aed", x"615735ae2ce10f44", x"4b689cca7b275de8", x"38e97d3c624e0e83", x"df92c1d3525cfad9", x"ff7ff5b61300b3ce", x"c2cbc1c470d74e20");
            when 4627261 => data <= (x"323b5179bf02ed5b", x"011a406348060afa", x"120216f80bdcacff", x"5f1a6509da1d8acb", x"eef6ef3100e592fa", x"0792a0952f850446", x"78e4de79dd5b391a", x"59d4e493d8845835");
            when 21297913 => data <= (x"98240e7d2c13550e", x"4610cc7abc634c41", x"54162d689c4bed97", x"e6d18dc002f55424", x"a6cd8cffc6d56770", x"a5af4b8327619580", x"d6e2fc6b6ff55db5", x"30535431ea886d71");
            when 26840490 => data <= (x"6d59333905438bcc", x"169cda996862eae2", x"080e54d019b6b4c8", x"6a20cf239f622002", x"824c31b1bc7011d3", x"bee0e5c56afb1d60", x"d9905dbce656ec46", x"9a9120ad57ebde7c");
            when 31611564 => data <= (x"18938b88c37cf41c", x"e156e3173a1d0b7f", x"e04641aca956975d", x"ba1b0940f9d736fd", x"ac4db7945bdc06be", x"925ddc01cbccc084", x"b58c8d7253e538dd", x"93f477b8d1b312c3");
            when 3914093 => data <= (x"b8cb574a91a7ce89", x"a183d09e34f34cc4", x"79630efb8d81281e", x"2d59f4998e9844e2", x"5aff0e27cb7a77ea", x"987ab98d4794ce14", x"e1b359bd9dc237f7", x"5074cd28cb79d20c");
            when 16432491 => data <= (x"95783e52d1372f94", x"c30de3fef6fa0487", x"d2a169b25c173287", x"8923b84e9441fb8b", x"981af70b0aaed93d", x"7492d42ec57bbe2e", x"8c6e0050a338e4b1", x"72595c663fdf96ce");
            when 31247711 => data <= (x"4eb77e7d00417214", x"46ab0c021d007594", x"066badf1f386df8d", x"1c0aed848bf2d4d5", x"cd6bd9aae49778ad", x"63fd508a9d7844ba", x"33acad8303bb9ab3", x"62bd2f786c77bf71");
            when 14935599 => data <= (x"00f299a3a1d65684", x"49f7323b5822240b", x"ab653cc38bc53838", x"aec004fa9d41a788", x"540a1ccee3951824", x"1f02957672a7e96c", x"691b15ed36702daa", x"252bdc396cd540c6");
            when 2689193 => data <= (x"6793db22f45b2710", x"7f15e87cdec5946b", x"d492b607076abc9f", x"f8bde756b05dc40e", x"40587b8d3181865e", x"cbd7681f2a7f48d1", x"3d085624eea4f6be", x"969ead6abaefa431");
            when 4153560 => data <= (x"1ddf0b302a94848f", x"e6dcb17b532f3b6d", x"a6858cb57b5c0446", x"8750cee27e065537", x"d282152b10dc43ff", x"1dc0b6a297bffe8b", x"9c96a9248dc5c198", x"45c826eafcad02d2");
            when 9721850 => data <= (x"cdecf580d16e6d33", x"c0007a5b398120b3", x"ce343748447bf8ce", x"f67ea778152c1318", x"f0c7cade749f74a6", x"bae0051b8ef2a8b3", x"656824f3a3271b12", x"2b7fc4fa9bc2e492");
            when 29449325 => data <= (x"cfeae3703dba4623", x"84602c8512009385", x"fdb1ea562c166014", x"b6d27d3a8440302a", x"d27c39895a670aff", x"9407f006b127197d", x"755a1e61b0a593b4", x"015c08e00c83d7b0");
            when 8277394 => data <= (x"604851e0ddea37e7", x"9367aada6281792e", x"e754ab5e2cc86af0", x"4f26b93d13a352ef", x"9f4cd2f961a65bfa", x"b0d1bb05c6c7ce77", x"f34691a5f7fddb16", x"93375edf73353ceb");
            when 24168253 => data <= (x"923bd2109fc7aa3d", x"d3019a5fa0c1aaa3", x"b5c560061d7ccaf3", x"d8bf2f922c40581e", x"2d52d743a0650ceb", x"d7117d588a9a15b9", x"104ecc98f282da07", x"2187bbfe2c07e6d8");
            when 8633730 => data <= (x"22bc684ef5fa115f", x"0a6adeef16ad8835", x"c26b9f7a3220db69", x"66c3cdb456c215a1", x"84f918d04d5adedd", x"cbdb547db842c328", x"575d79ae114d36e3", x"0442a0246f90061e");
            when 12650671 => data <= (x"f4b0d1469ed6f3d3", x"419a0b6af527a245", x"1fd34c842252e2e0", x"1a2a59c117959f3a", x"70541f2510058b16", x"10c75cbe075a86e1", x"60e24d50eddeb019", x"8c0d8d061bc3776e");
            when 609109 => data <= (x"d09ef9ec6f3f245d", x"82f0c339a521c748", x"a45bb32a699d6b09", x"854a8ad6ca6faa21", x"58a9e615efb302de", x"a5de5eb7940ea105", x"f567ecdf57fa0ef2", x"75e231effe352b90");
            when 7977288 => data <= (x"79665188ff700df7", x"ef6d6d862c62ebb2", x"df92262c93f1f6f6", x"b00716deabb23ce2", x"92b2fb3d274444c3", x"05317ab48f9d7190", x"b9e9bb1e60e23ee2", x"31f2d830d6abc1cf");
            when 11660162 => data <= (x"8fa567acf8388d6f", x"de5e930d36739afa", x"ecc2ba417731720b", x"9a9e06ddf794dc37", x"c4a356b245fc65f8", x"5e2a4c9fea8db1ee", x"ef7717420e348830", x"312f801bf7cae37e");
            when 13628157 => data <= (x"fead8f21e82a1a58", x"d391a6b3cfdedbf4", x"cd6b1ed1052ff8ce", x"72cdf51cee79da2d", x"1be8e9aefcdc73f6", x"4601759d5eb78ce2", x"3f51a2af68877af6", x"670c432f5320bd34");
            when 9488955 => data <= (x"4e7b276f83c16a4f", x"12e09261f84231c2", x"2cb94796880882bd", x"473c29188a6b0212", x"dc0287463438e54c", x"5a13615d6b7a73c5", x"6d86de61ec9106dc", x"ab1f82690337e27f");
            when 27875635 => data <= (x"5b384a82e7094738", x"8c22bded9a5e4e54", x"626686273066f08f", x"04bbef41c46d0fc3", x"9bcb82ee873bea22", x"10f6dc324ca819d3", x"f91fb5f18450acc9", x"d3f1e609a82ee345");
            when 1905767 => data <= (x"460615a5bb4724de", x"a1e1163e56c61340", x"aa1b6040309bbb3d", x"b079c55eb1ee94bb", x"b0930427a69a4a5b", x"9d9787f7ae49a744", x"e7d80410677356f5", x"cf50e527eaa81aba");
            when 25764372 => data <= (x"cb68dbfd687568e2", x"75ed961db3a362ac", x"0a49f0864606b918", x"c6f0a7ab4356f917", x"36d38ffcb025c1f6", x"61807739119636f8", x"290f2879ebff3fad", x"da72204652a02a45");
            when 5055437 => data <= (x"cc364f4b0214217c", x"ac0ec67f0106a9e1", x"d7b13b6fae456ab3", x"2795042c19e1d988", x"948e28e952b15a97", x"55a72bc8892a1ca8", x"70cd1434800e1e2c", x"eab97be6c4ddc725");
            when 7161741 => data <= (x"7d21999509b56b55", x"36b4f070a9f05505", x"e1745555f4c1aec8", x"4103d1c2971464f3", x"085d2117f5d9dc19", x"30120e34a45f903e", x"841e71229476c25a", x"485d56839d30e75e");
            when 20139770 => data <= (x"df9123fba5346c09", x"290105e4e688bdec", x"989386d3aa913c69", x"417b2e318921408c", x"3c6b67e249a1b472", x"4ee305ec7362704b", x"8798da82f3d07bbb", x"f36ca11e9877f513");
            when 22728474 => data <= (x"5bf59f54c458f193", x"32a37eec1701ea6f", x"4d68739718b0603e", x"d8e99a905c2d6cad", x"a096a3325983bf10", x"ad5523d384ff063c", x"61bf4e6924722384", x"b6aff9329f24a07e");
            when 16167873 => data <= (x"3f8b8fd491e26065", x"a1f5a99c1b74cfcd", x"09494828987a497c", x"22d8e78ca655bcdc", x"b237165cf89ee837", x"0188b93f8498c753", x"f43252d5482197a0", x"81dc87d4dd59109b");
            when 27153716 => data <= (x"f27c14cc6bf957a4", x"21f36867e441bbb3", x"ec871ed46359a62a", x"9bd4de3fa4e5cdf7", x"e5ca8fe4650db42f", x"328a21188e6bd649", x"88e851bfad1f184b", x"6574a4f83e74afe8");
            when 28285872 => data <= (x"05249e49ed179d58", x"ad0477b592413f0a", x"292183dbed5519cc", x"f5cd7f427c06de69", x"361ca61fc6644d52", x"b2a578d82bbb1fce", x"2191d60d2b40b3db", x"7865db3014d27521");
            when 29365305 => data <= (x"44c255d26b4881be", x"9fd5bc3b8238023a", x"be5f8c0b95b9251d", x"27353c7845dc6d86", x"4234b9e346125bee", x"537cd551db9ffe2f", x"5e956006a1f5e780", x"de6b1ce16f2afc53");
            when 14274789 => data <= (x"9f4f39db04dd1b4b", x"a48e0ef4b118b5c6", x"03b6ef99dcc6b352", x"d39e6481d5905b37", x"7925c40c919eada1", x"0252fd0910c0d3b7", x"06fcd9c66c2b3f30", x"ac888b25fd39c91c");
            when 2746326 => data <= (x"52cea786de280fba", x"6b62926f08a90e5f", x"d33c2a5da887c75c", x"9ca3a033501585a2", x"8d7355d4573b4ee2", x"8583e818c5f8b987", x"4854abb9fcf846ee", x"9199c40a70921c9a");
            when 26447896 => data <= (x"b0776b4e4920a992", x"095aed34fb71e0d7", x"a54314ea04fd2b1e", x"d9652abd82018d79", x"645525c4e28abbf4", x"83e766f0df3c32af", x"3edcb4bee17d8866", x"8fae9c54a5d0c3ae");
            when 569241 => data <= (x"d3a421109897fc07", x"4049192cb1d8264b", x"efc47eeaaf3b8d44", x"0f0df56d733819b8", x"06d46d2ee2585ae5", x"5e55780edcac084e", x"6dbfb5902128885f", x"c55b51422db04477");
            when 24561665 => data <= (x"20f4cd3abaa1fdd6", x"5a6fe4efdf3efbe0", x"e963c129f20d1b20", x"90d04372b3f8f212", x"a95d73787607cc2f", x"3d47a5e3a6febba8", x"a2cb19b83b8e050f", x"9904bc47957c613d");
            when 4281348 => data <= (x"2284f79eb12b8421", x"f5c83a22536726a3", x"f3aa7856318f5229", x"a016e98e7bddd574", x"2472317886a6f1f3", x"453fc15294fe505b", x"65cd6b38bf0adb5e", x"dc8cf82488673c37");
            when 9069463 => data <= (x"52bd1f2ee8f6e194", x"1d7f8e02bfe58a64", x"a9c77e322dbe6386", x"bf5e9cda1137513e", x"d4a4ad16f830f385", x"46f1e8d5ed1b9eee", x"03ac22dd94acb875", x"a6bd6fa387f3e4d0");
            when 27484790 => data <= (x"025054b433fc4752", x"2bafef9ccbace089", x"45b20bec804dde28", x"36e9d255a6b765fc", x"577fdfd8291bc51f", x"c3d359a43a198e77", x"bd7cf42f2b1b2ef2", x"c1d00030c9d8977c");
            when 32948412 => data <= (x"f8cd5d42f3bccbfd", x"ca7e63a9abf3e336", x"c4e92ecc7af88020", x"6a368fe00ad8fc26", x"8fa2fce430b8be96", x"903acc8a7fb1ddfb", x"aa2c2d288481e435", x"44def767b5dd1412");
            when 14473511 => data <= (x"c4e2789427f5ce99", x"1adb7bee973dcdec", x"8ec93247dada1119", x"bcf91a13609e961d", x"157481da59491d02", x"f422a1869020a1fd", x"bb8a6cc4c3612e3e", x"e2ecd6d47fed75f9");
            when 12562154 => data <= (x"141517790179390c", x"cf80d75ca0492bd9", x"691c09eaa86ef443", x"e364b42fa0507bed", x"256bf3fae3e9aaee", x"7c8550e9d21de935", x"be38641cddd1d405", x"2dfef97deb638c2d");
            when 18548696 => data <= (x"b4d4ea35e803bc82", x"a40a894f6e45454d", x"b718309d97fdc76e", x"147f1001404d4330", x"7d02c8e5dcdb6f50", x"7373504d061fbc37", x"9bb93b889d6b1394", x"02272f06f9f73288");
            when 15074929 => data <= (x"3dde83958cea712f", x"9209ac83d441ded4", x"b8823969f83c0940", x"e9b51b9d1a417326", x"0fafc158feed3e6d", x"1e7ef4026a8d0779", x"cfb1c30a8b3ca689", x"3eaff862cbb56158");
            when 9596254 => data <= (x"4a45f6349b6734f6", x"c020c0e9a9abe750", x"9c0d7b7ffbd66a8f", x"1c840ee196ae6c66", x"dc2c307428b09ed5", x"c78c6c7e17a83520", x"4d4c40598862659e", x"9119da948d1c58e9");
            when 10759989 => data <= (x"3d55ea1bed6fa1ef", x"68261ed529e9d2b8", x"5ef0414a31671f88", x"de7d950add5415e8", x"465641eb16c41b13", x"dff445817f6a88f2", x"24e2b3624e73940f", x"b7cb3c7059e6de7f");
            when 27055604 => data <= (x"4d0c3402cfd42217", x"557c66165ac35b26", x"2ceda90a0536e741", x"7df53c41dfb0dbc5", x"d725a1717e992d9d", x"fb5fd29a3b5bc7fa", x"c408ae828227905e", x"4346561a29a0286a");
            when 11055641 => data <= (x"32426a9c5aa4aa65", x"f95275bd3976877d", x"b6612c7bdc768a0d", x"dd62d3b87121c73e", x"1dffbbe5bd0c1028", x"d2a65c94f626b650", x"d6ebbe7cf1eed4cd", x"0943e243c3590007");
            when 27716722 => data <= (x"025cf37de3b2efe7", x"4a9b3ec66524ba76", x"2488eb3d877553a4", x"eae2bc9d77ff7931", x"20922fc19836855e", x"df4b0dc5b6d3dbb7", x"01e62bdaf7d8ee3d", x"620b0f95a237d235");
            when 348832 => data <= (x"2eae1a277d22b8f2", x"1b2ffd644790a6a0", x"177dbe820929ddeb", x"7e658e324f8c8547", x"55e41ffad7cceae1", x"7660d8876dfdd946", x"4ccc7af309d7859a", x"2c7f0da238e13c63");
            when 1547044 => data <= (x"e1d0b85a40b2e965", x"c651bb3cb2713528", x"58862f6172918702", x"29ea98bbe490fdaa", x"d7ffcc62b5f2d069", x"5dd01d11c145cb41", x"58948deb92655861", x"e6fbac3d4ef04801");
            when 16202929 => data <= (x"1b4338d6cfe7c720", x"94fb0ef01e68e29a", x"8218a718c0178949", x"84ca58b4292ff015", x"d0d452bff1a6a177", x"4ba5feca4da4556f", x"f12635766d176662", x"f5f8fff25b3e2879");
            when 14241533 => data <= (x"1597529795a2bc54", x"6ce3776d12b7d6a2", x"578d4c94a02010ef", x"d6f8209850f6bcbe", x"cf2ee14fc80fbc76", x"fa71b963785dd7d8", x"5d1c2f0c00ab0841", x"2426da0414bbd755");
            when 6423156 => data <= (x"6a9ed6791f364055", x"5e94fbe3fe47a6f4", x"01a1d56b37a02839", x"557ce3e18357222c", x"f44ff45849afe40a", x"eab1bc2c3aa09229", x"797972293bed8541", x"63479fc05535ada2");
            when 32354768 => data <= (x"c8e6be3ed60c24d1", x"97179bf66095c63f", x"62bf05d46c9fec55", x"d218073d0320af9a", x"2f1b118614d4c25b", x"c84d0ea8e105dbda", x"1ad7eb70f785e7e2", x"b0ab155c65951c58");
            when 2723151 => data <= (x"7ec7c2d94803fc8d", x"8b66642db1c3be1a", x"05afcc5530e5881b", x"b4bb2d1719e2f350", x"8714d2fbf65c47cc", x"5d8508b0fb43d137", x"301fa554979d4b12", x"970a13e147c706c8");
            when 25105451 => data <= (x"880bd0a969a57a6f", x"49f9091205571792", x"bca1fd5e06075298", x"d4f494ba34dc94d4", x"36cddd4ae96b3646", x"d2d825434420bcf5", x"3ff2bc76703333d0", x"db2f96bf8f5ed30f");
            when 33537111 => data <= (x"04c6ccc8c9cbebf6", x"a027815cbf5937d1", x"f051dcc1dcd4d5d9", x"9f62775a10712b16", x"85412285f8462607", x"7b8571d55d95c863", x"40dcd2ce4a9c3e51", x"531ed57f328e3d72");
            when 578683 => data <= (x"4e936f3e7fe957af", x"80f633c91ee3168e", x"58f40f85f7d78bf7", x"819e88c6daa62306", x"cd5567274ec3b23f", x"bfc9640fd59058b8", x"b182bec59b2462a9", x"3eef3b07d113f1d2");
            when 31831512 => data <= (x"2bef1ca737e624d0", x"886fb75ba1f2107b", x"07d1b05146ea9c9c", x"7256ec1e79d40154", x"91f92969dcf0ba28", x"eda7eececc412d03", x"8d13a97fbe3d37bf", x"3e0dc26a9cea8b99");
            when 5493286 => data <= (x"272fd724a9c0eb3d", x"e51a57e115e42ef6", x"0e947a5820c993b5", x"4c97bc1a6898d01c", x"311a486bb8a3ebf0", x"576efd160d8605cb", x"7feca3448655bbfa", x"94faa086fb0d19b5");
            when 143290 => data <= (x"f2a1e8af150bee73", x"d7016ed06cef4d99", x"302fc827f6d7fd9e", x"871dd18317405f44", x"a5525d5ca8d32cde", x"4a46c2700d37b674", x"d3d59ef8bf5e5382", x"74fd4cdd3b91085e");
            when 22778168 => data <= (x"4837cfa59f6b7ac3", x"c85fc8e8c86efb8f", x"78c06a16c74a9db2", x"0f33d7ca2d8ce96f", x"1289bf49dd0150b0", x"ad37aeacb2b63f83", x"3cd486388ffcb07c", x"2d65d783328322e8");
            when 13093099 => data <= (x"5b42019040b0b03e", x"f5e7f5797cbdcec4", x"2afc80608506a2e7", x"ae5a71efff456550", x"6b62fd1999aaa221", x"5b785abf658f64d6", x"9274ec78795c7db4", x"c55da42ef46c29cf");
            when 25921656 => data <= (x"568005a18c2d707a", x"cac72ff8e6b936e6", x"e0e4c646bcd1ea35", x"eddfbdac9da7e6a7", x"fd5bc240a93a0d82", x"861a0814ec7c5001", x"167db138ebdeea4d", x"8139cc3d6ee11cac");
            when 19835364 => data <= (x"d699dca91bcb1b48", x"285ea9272bcbc4a9", x"ed1ff7f66c7d21fa", x"8482334dcbac0bea", x"2db302d79835f816", x"3e08f846c787e192", x"3e71308aee6e6890", x"940ad893c13e77b9");
            when 23326403 => data <= (x"e3db3874fca4625f", x"28a98ac672576d80", x"0970308a52331760", x"1d9b6aa26e5a0149", x"b055c94c9163a209", x"d85b190de5ac3e20", x"4827dc734618a8dc", x"d22d90ecd2a464c3");
            when 24181901 => data <= (x"8694f327448f5c22", x"92293bc11c9778af", x"23fd81eba09bbb10", x"f64b859949dd947e", x"9dda44f10808f4cf", x"2b7213c1662fd7be", x"cefe0d8dbe2fa943", x"650b92282d51c9a5");
            when 3261488 => data <= (x"c28ec6c40d04b14e", x"bded2590cf6a3d94", x"cbfa1f1c3b26cf98", x"9eb088d82a478ecb", x"57e960cfff00ece3", x"a7fcd4c8d0e7e260", x"499fb23603de8179", x"64b0ddb247241712");
            when 15771043 => data <= (x"f8e993315940806c", x"6ef6297a4f122b5f", x"1c54011de92ae88c", x"0c1482d88364cbb8", x"c21bffb61f64c96d", x"16630bd9f407f93d", x"2ea2ba80b9721309", x"5c7769d0232d8524");
            when 9625704 => data <= (x"d652f76ad8f3dc43", x"f9e33389c1fefa07", x"dd83178269221645", x"2013908412bc05d6", x"c2f2c25dabdb9ad6", x"b512905233256955", x"8e02f7b139998586", x"0838105d61ff9520");
            when 11398095 => data <= (x"bc28f68e8ebf32d0", x"40e8975fe9b5c462", x"0023bc42b18ec275", x"3a04ede9a0e8db34", x"4de4e9f5a934b968", x"0f334ac9fc170f60", x"3b89268e1f680be9", x"9f372041c9f224c1");
            when 24536519 => data <= (x"c02ab98b15b2620a", x"baab743896fe6a6f", x"60d738f0b6a55543", x"1bd58a984d323f11", x"457860ae1a684490", x"b0846aca986aa41a", x"c4b562c4633193b5", x"5d30848fb13c91bb");
            when 32983960 => data <= (x"9498b1c77fbadae5", x"e14bc90d1fd08dfe", x"76a2944308dc8f7f", x"572d9b72d33ada0a", x"93a977599df8b34b", x"adf9774107424111", x"d5add94934254163", x"e7d5254bdd2af770");
            when 2685290 => data <= (x"7c637f14818de6e5", x"cdf5c76a5db2186b", x"c8cdf87bfaf7f656", x"b97496e9bfdd047e", x"aa692299d94c6b8e", x"9affe109778fd087", x"a467301e3fdd5a41", x"c80b896a769b4ae3");
            when 32532854 => data <= (x"6fc2531dc79aaa72", x"3da3e3d7fecaf4d0", x"810db5e69b0b3764", x"84cbe42f919e7e91", x"47818efe3da99be6", x"966cf5ce6a7b1da3", x"a8fa6628afae4c6d", x"d42ee41f5e0485ac");
            when 13494968 => data <= (x"a684a258577f1715", x"35c30b15d46b294b", x"1441485097fbd370", x"25455a5f0ab9cb15", x"27b78255d812ec99", x"19866df9f4d3d862", x"a973df32c8a65dce", x"f6c02640416848d4");
            when 30491318 => data <= (x"247c81f93cf4fe52", x"6cd7c4bbe9077d53", x"3b2c336313cf5853", x"93f45974ba0e2c60", x"b6400e15fa736985", x"0df45850eff5ca4e", x"afec34a02f501b01", x"e01c94e36c1aa36e");
            when 1744381 => data <= (x"462930ae283ea22c", x"e262f16b7ed3eafc", x"7c8468d65a41376f", x"c30f3ad8492b2e99", x"6a24f4ece9389203", x"484b56fb101de126", x"ff8cc797dba34834", x"9abf74d8e9da3698");
            when 21901686 => data <= (x"c654fde2c1dcd583", x"a4a05ae903d70d49", x"3cbbbe994d7c0aa0", x"5bb74cf4b454cbef", x"e20e68b4d074ff4c", x"d14b9d1a4ba0d817", x"3a8637d7a29b97b8", x"2126656eb82deb4b");
            when 17148493 => data <= (x"359a7634b3942920", x"c19f707bdd601e72", x"4708b4addfb8eff5", x"0b60bcd9d488bb74", x"26f25bbb38fa4158", x"98712a6673c33e32", x"4e0621b2ad40c534", x"a103dc28059186a2");
            when 6604179 => data <= (x"9b19175894e6574d", x"5ba312472e214f1c", x"eb0891187293fa78", x"c7a6c1fa6449c1a3", x"906b33cff7b9b8f9", x"a4e908f1e1741445", x"3dba4ed4b180c2d4", x"d1a25f5a671beb67");
            when 25989844 => data <= (x"69c05f9d3859c09e", x"9f7cca3054ba2968", x"402d8bb053f65eb3", x"0350106d483ba95f", x"d664e4f2e4a4051f", x"f91b94c0d271bace", x"b2bc86bb62a556eb", x"4059bf5e7aa9558d");
            when 4644463 => data <= (x"13387dfa779cb910", x"b37dc34ce8c360cb", x"2f388993f7e6ffef", x"be6388ce394bb5ec", x"1abb1366166273b3", x"b065024c16282d50", x"0ee83208c3d6d10d", x"9f3bba7d65cbf301");
            when 3691587 => data <= (x"daf7b5c9ee34efc5", x"c9e25e8e0e612484", x"8cf8da307a69d337", x"b7cfb5508339f898", x"14ea47efc571a6cf", x"e22e118c1b8d97d3", x"9800d945ac974d05", x"f07ac40463e1f9e5");
            when 30080383 => data <= (x"d4713873d7e70623", x"1a31532bc80f1aa9", x"3d6e6d69be03b375", x"51a778912350af87", x"708dd4980855b6b2", x"2850922d7d9ff931", x"7a70c3209586f2dd", x"634ab12e899a3092");
            when 4080703 => data <= (x"80a0bce3c1057f7c", x"c66f96cf8b622db9", x"2a6ce4b9d2a40f50", x"0b42904727de5d41", x"55d9b420548027f5", x"bcf1d3a662d84924", x"d79e124f619f022a", x"ea579b346f140948");
            when 33544278 => data <= (x"95d70e561d021b0b", x"64fe613cff8fc621", x"a0cc9f6e1ed9fd95", x"8da4cea84cd3e320", x"c41f83d779299782", x"be7b21b08e4b2edf", x"d89eba71a47e7ce5", x"b8dc6d0be0082840");
            when 29818877 => data <= (x"ee13e60c945cf162", x"21706217657f70a3", x"6edfbc6fa18e85ca", x"05ae01c762288129", x"2ac926d9b99d67d6", x"3950240dfe95b7d6", x"24e48614e8a75a08", x"8c57f8c987996e8f");
            when 10863342 => data <= (x"2f130cba78787661", x"cef25964a215c947", x"1e11694f6aa3a6aa", x"e012c13d066991e0", x"44d5dbdf65aa04ab", x"621cdd212c6d30e5", x"fd58398d63d580d3", x"e209141704c04b13");
            when 20578260 => data <= (x"0c383ab570bd7998", x"b305fe37a11e06d8", x"5e37a296ce9d3fc3", x"362b718cb0d3c001", x"31c396599dfbae42", x"2634a1248ac84a1c", x"2f6b9b2860873b41", x"97e8e2fcbd9313e0");
            when 21290827 => data <= (x"dded6b7423efe532", x"ffdfc55f2c4e56fb", x"f73547ac7f53bc43", x"5fb9e83b020a5787", x"b3400cd71ad18e98", x"c8de65a1a9b83041", x"f9b65043b11664cf", x"b5bd664edfb4d9b8");
            when 22560855 => data <= (x"aba6d6256e974405", x"777b491c3e860793", x"187a6a02b8b14b67", x"a90d984a0e70f4c9", x"b274f9b86bf6f9ad", x"1ab00b06b1df85c1", x"f305605d6853c6b9", x"4a5a572d8d994ca5");
            when 27823124 => data <= (x"14512bf4d43341d6", x"64f60381068f5a64", x"9fadb5ef591916ff", x"3b0439e12bafeaa0", x"036cd25aa1e9934a", x"8bfae0f8e635adf1", x"a878e04c23839b9c", x"44ec1d1f05d690b7");
            when 31834667 => data <= (x"f3712d68b43a7432", x"a81b8560af5271a3", x"3992e39458b54171", x"2e7c53d8fcf0a910", x"27825b600365ac81", x"97af3d4741bd3610", x"ce6ad57adec2202d", x"1f5efcdf26fc6d3e");
            when 503338 => data <= (x"aae8ae8608bc27e5", x"a6a32d21f1ca74e4", x"43ffae0abb9c0d5a", x"29f7ef703fa4ec51", x"ec1a4d1ba5da5331", x"d3c9ee145a82864d", x"d645d7417a4507d9", x"0f35b8f02eb93875");
            when 18455406 => data <= (x"bd6fc7cc36bf11b3", x"d10d6f3c49f17258", x"ed3f6553a1b6e64c", x"fdba20001f01d28b", x"c973b31362a79c72", x"61ed7c48f6e1c519", x"157acb66068a6718", x"0284489d2f575917");
            when 13296354 => data <= (x"d236ab2d9ace1575", x"64ba79c36e1d5e73", x"1ace4bf9c30e9188", x"d72eb62d22e8a118", x"7b353e985881e5f8", x"a3d47b0c4a669b2a", x"148c8e80b78c9143", x"23e796754d03020c");
            when 4031974 => data <= (x"022d037417d75d43", x"b604bbdaa1251150", x"534effe75d8cfc54", x"1cbbb313914793db", x"3bb76d243af31555", x"fd6aa8fc88b80638", x"03bf546eba8c4fc3", x"6ea66ca1c8664c0c");
            when 28365394 => data <= (x"23d2a8eb4c367a66", x"1d4fb9fd8321d617", x"1a6a39c58c0eaaae", x"2a0ec055b6199f88", x"10a59bb17f58afd7", x"418534fc785135d6", x"b453a0c29de99c11", x"dc5c18b2e5727032");
            when 32845200 => data <= (x"8df631d21f956f3a", x"b078de071673dd4a", x"8054a6696b6a7f3c", x"3f03ff7e7103d7b7", x"d460074fcac96dc6", x"f45687fe8aed368e", x"7ff984055432f60f", x"00c00e69f90382aa");
            when 4464092 => data <= (x"a07eff9524371f91", x"db7f45d60b5342e9", x"854786deb2bff850", x"3e10cd7a99ff7776", x"f54504b09a9feab0", x"02e1a8d30b2365e7", x"6c2f6f3bd87b11d5", x"713ef6016cba6ed0");
            when 3715652 => data <= (x"6a88693bb2ecc667", x"83d6d64b57066c67", x"6438cd0d8b2de895", x"ef4bb85c7b09b936", x"b689c50c8d32ddc3", x"628ef7e1499ccd3e", x"d6f47b7fc7fe3e84", x"b99e11e7e82d64fd");
            when 10756860 => data <= (x"6253f5ae8d9aca04", x"a6c91cbe1849fed8", x"e874ad393b48783c", x"a96b81287ad53639", x"90d1a9d64d096eb3", x"bab6abf743cc7624", x"d6ca14b63bcbc547", x"21ebc6b92b710be1");
            when 24634131 => data <= (x"9e0ee1f27a0ab85c", x"e6e34c72c1fad6ae", x"fed7779f2fdab7ab", x"4cab5df8620d352c", x"d34d5e1fcac9c47f", x"da6c4176daaca0bc", x"a8e83ac456160cb9", x"35897a049734f3a7");
            when 11145390 => data <= (x"d4cb263a987aa0ea", x"e3ad57da51641d1b", x"156430dc31db74ae", x"23a5df98f8eeb5ce", x"d6294a6798f7bdd2", x"840af632acba6311", x"e166a521e5139d07", x"289b4a5a0399a743");
            when 7163262 => data <= (x"632d6af0ad0f61e4", x"20ef3288636b790d", x"4df86eceeab498f5", x"df890f9ddd2ce5a9", x"c566c54b07966272", x"e36b06e4eb4fba55", x"1860995c0a801def", x"f251f9091f5cdbbc");
            when 31221607 => data <= (x"2dac7aa1c2b7bde6", x"373e4b101a24ac99", x"0944be669cc9ffc9", x"c1183e341c79fa75", x"67bcec3f317a117c", x"98ad9b3856919191", x"ee10f6db76acc606", x"5db157495f8eb1d5");
            when 14723323 => data <= (x"e3f1980cf57e0242", x"5f52541ef8ffcdc2", x"8ca5cf14d9e5fee2", x"b61cc47c84030e1c", x"a25f00c784c6e03b", x"a51abe5548571308", x"f11559101de4af1b", x"bb9aa40055b232bd");
            when 22813550 => data <= (x"c4635b1fd3be38ad", x"eb4fb746c1744ac1", x"40e60f8a9d167b60", x"24d55181cac6e576", x"41bbe26883785b0d", x"e9f694610e663a35", x"4d7e86c1126f332f", x"eaced0ce9b92edf2");
            when 31904467 => data <= (x"ba31ac1e07e556e6", x"e2542366a1ccbf60", x"aabcf262c2b6cd98", x"261b4326059953ce", x"79b07120becf8a3b", x"52aefbb4faee1826", x"94983c1bbefde5cb", x"bfc2b0ee21ef0217");
            when 9432147 => data <= (x"78cb39533e98db52", x"97e84b4940fe9ec5", x"53b9da4ba96fb37b", x"0e438c05eb9525a7", x"19cbb51dacea4942", x"0a2dec5351e85188", x"46ec93d9ae779812", x"384765b4168eceb1");
            when 7802337 => data <= (x"3a1db12d127aaacb", x"e1053f935f36286e", x"b9d50bc14e23c994", x"1c69b8efddb97308", x"c3a69d6af5f827f7", x"dd288a4135f2ca59", x"95c68154c7ef4568", x"6b0265fcc50f2d86");
            when 17000769 => data <= (x"50e32c5817aeb2fd", x"44d4680fa6a996ab", x"d378af34d337b6a1", x"61227a40e16d4b7a", x"49dca4cd95bf3632", x"a98a9f498e24ea0e", x"f7e37cf6fc665b4e", x"6267250d844ebf80");
            when 14280773 => data <= (x"9031c6d60eb3fb11", x"843a01de2ca9129f", x"47ca9336827b2542", x"220912a893cafb87", x"d05d37ae95a1127c", x"534ee095bee6f8a9", x"3e9899ca7038acf8", x"01f77ce846510534");
            when 10194617 => data <= (x"d59f81f8e4585b4f", x"dc57cfeee765c60f", x"9be6cbb6c3a5f186", x"68d6f5565ded5cf5", x"d817e5106ecd7690", x"fbfdcdee59e11879", x"c6d93274ddfce7fe", x"c52ced93baa134e9");
            when 22154183 => data <= (x"db2d6d2a5a9c0a38", x"59f0870bf4ec4360", x"b210a661d5e26de8", x"4ae8fc251e765565", x"c5cad86962a9a74f", x"7e7e5a274893f3f6", x"34e926ae9243c540", x"317afa5bf7bc4bcb");
            when 11871082 => data <= (x"c24812dbb5aa7b2c", x"42d4ada4fd718a50", x"048c16093e5b7b66", x"f43079492f85cffb", x"18bc6cf757f875f9", x"bc2a9e9771f2e2a9", x"432190a5dfa64848", x"0e99ee6b15ff7e6c");
            when 29544524 => data <= (x"639dd6259c5431bc", x"a8e639cb3c687091", x"44f32318298901f7", x"0402678685317c14", x"5185633f6bf5572f", x"bfeed937fd66fda0", x"d7db9e9504a3613f", x"cea0d153e4215d6f");
            when 29581856 => data <= (x"bf5aeb056ecb574a", x"f4a883775213e833", x"62f04eb4642860af", x"dd0fca41fbc5601f", x"30e625a2158fd065", x"af9e1001ce41866a", x"50f96a84edde2050", x"79110199aaab4f98");
            when 32373082 => data <= (x"10521f385707af33", x"90decb54fcb4eba0", x"4fce82b892049b02", x"213c9bbbd99c2e91", x"dfd927cc87c61d4e", x"a9dd574331ae2622", x"c1bbe66f6278dc55", x"45e91417b011fb35");
            when 7798782 => data <= (x"107ae7dbe393347a", x"7ceb4082a5ebe6d3", x"1018fe249e556de0", x"83c59d5dbc60715c", x"25422fa63bf2d7c3", x"e9c3111186a1bc49", x"2246be9e713e3346", x"1f6920cfc4d94135");
            when 18660735 => data <= (x"d58a4eb6eb6dd5d2", x"1ca7265ad6dce0b3", x"04ed30a9edaba854", x"3940cf93ab675ee1", x"d4f9fd7b2f219d2d", x"8525164acf743fcc", x"619e8a04bda4eeb4", x"3209c377046fa628");
            when 4749909 => data <= (x"92ee4215b1ed3383", x"9d882f687c29a36f", x"92ede13b0129f3ca", x"1440b097ccc2152f", x"b9ad1a8f77472c6c", x"09ba405dcd6e3865", x"80ea3fea16d42c50", x"d0000a2a6e7eb034");
            when 11667057 => data <= (x"c50080b88f2b1e82", x"ec69493c5ef87d62", x"ebd23a1c437185d8", x"5cfd59058c0c6a01", x"f90a3b8705c39705", x"a9faece3fd40dc82", x"715a6699604f13cc", x"b679f25905731598");
            when 20116957 => data <= (x"ec6983fe611b2cbf", x"7fdff9808f0c8cfd", x"bbb1dde3fe59df8f", x"5c75415c7445958c", x"72d36411997d016a", x"a1231d04d4cb5374", x"ebd0428fb6ab4529", x"63301ae931a473f7");
            when 9365883 => data <= (x"817b41971155fc90", x"2865f27a67a74d14", x"a81d579a5237d14b", x"b30143999d7c2d0a", x"3889a32780f6abb7", x"26e10948e1d270da", x"ee72ee3e605f1bec", x"c5428ff3f573c5bd");
            when 17258373 => data <= (x"b42513f424b2aede", x"9f8f7ad90f192ad0", x"cd91f6693b1721e2", x"4dae32a1345b8a2f", x"78aa29840a5b4bad", x"4d2eab89f845719c", x"91337e21c9337e56", x"a7205088116feee1");
            when 27833760 => data <= (x"023e5bd247068d7c", x"a9837aaa73f9cdd2", x"0ee57ca45c2aac14", x"d88ff9dee92fb06d", x"59956b259ee20d57", x"b1f918bb1694640f", x"ba8bce1759dd9b1e", x"8b1efe0b9ef86e58");
            when 21197741 => data <= (x"31875c8b2a75e5db", x"109a05346c4f9589", x"076f1c51dd38417f", x"58cc795a9f53b03d", x"f00b92dba2d4010d", x"95084d83729d5c0f", x"815175e26db9ec77", x"5ffc7d8e0190100d");
            when 17436478 => data <= (x"58ed4e13b755b4cf", x"5ef98079802eeaec", x"ed94dd168f43c161", x"ebc3f2ebbec798c5", x"7fbec1637b643028", x"d29bf0b1dc68bf20", x"b8dda3db03ad7c3f", x"cb3d220b0847d81f");
            when 27556440 => data <= (x"a2b9f898551234f6", x"2982027e9dc04d3f", x"ae47484de3ecdb79", x"ad9ef1aba516c80f", x"7a5de2a9bd1b740a", x"f87133d24dcdefeb", x"d07e5641dece6b80", x"8a12798918a36833");
            when 5130799 => data <= (x"de0a3b891bf62a3f", x"97e3e3346467a009", x"cc2a1972f4f16e87", x"9dde377f0506d470", x"b1828c800b35823e", x"84477c2305c0b966", x"dda8e01b8bcd02f7", x"e880e40d3b76a560");
            when 1857135 => data <= (x"a03ad682ea5324e0", x"1bce02b5b7f8d0ba", x"19d00f8509bf32af", x"11c7d4cb3fce84f9", x"ecb481fd2b869bd0", x"126287a3d8ad7d87", x"9acdd9cb941b300b", x"65cfd45a04ada649");
            when 3335680 => data <= (x"155fe2f1740585fc", x"2afa2ad1ae330f7b", x"cd6d33d247129d1b", x"db88021bc286e7f3", x"1dfdff43cd73bf5a", x"d327917c518d2571", x"6f0768789e0b22f6", x"6a791e78aa8b9390");
            when 13633015 => data <= (x"935fd761d8b87798", x"c2c3d236fd4523ea", x"0de24bbb6166779d", x"5e370c90ebcf80d0", x"6ad2e228382954cb", x"ddff2772673d30e7", x"604d276f59c635fb", x"ffdc46531a0fe71d");
            when 19634095 => data <= (x"afe8356f7d2b9479", x"897456dbec4e7dfa", x"06008dd95051060a", x"4d872ae0f5508249", x"49a6e94fd733d066", x"81c5e8900c25439d", x"ec5044618f3b9d54", x"3c58a515575d3fbe");
            when 10534679 => data <= (x"99ee5d47e86211f5", x"c48d0f5736097e45", x"ae5ba675442258b6", x"48ad9ae56c066681", x"d6b306507a1d6ddf", x"7176e8481053ca8f", x"31fb150fad234045", x"c95fc1c7c2424044");
            when 931116 => data <= (x"e1322cd0a41b7bf0", x"20b37d524c94a836", x"731a2bf0b3aa94d3", x"3c083fcb14a73777", x"70178c5ea5df4ddc", x"32268e0049f5ede5", x"294ecb0cca4cfc9c", x"49af5584cd36e010");
            when 28742765 => data <= (x"af867e3ddd6266dd", x"6c50696ec40ec82b", x"27267e356eb01c60", x"9350098673ca6b75", x"87bd0199b8953d87", x"b79fa91ed44846f4", x"949ea91123281ad3", x"aeaf553874f3af3f");
            when 33215902 => data <= (x"b226d456f20f5355", x"c93a09335927982c", x"4e52de753a3c2861", x"5c37f2354f6027d1", x"274ef6901182bc1d", x"1c708368d2fa0a89", x"36f90025d03ed86f", x"8969ecbc8a8df369");
            when 30010039 => data <= (x"77a3db2b635ea4f4", x"eea35ab58fef611b", x"05a9775ac258b9e7", x"264b4a77896994bb", x"e63a305876082bc5", x"9c6f6cb51dc4ed03", x"4ff1f69ab26e0421", x"e22d94d0e3e0985c");
            when 31430046 => data <= (x"6a5939e6ae2a10cc", x"be5575e166787909", x"c0a2a1f095a81f3f", x"842b5efdadffcd9d", x"717ac30f44acdf45", x"9eabc570ee54482a", x"715a43737e859413", x"da0d9edf14ab7e08");
            when 2135221 => data <= (x"a6a8a45dc068fecd", x"76fca5867f27cd7d", x"db6a7e0e2256a8d0", x"9b77d75278a59cf4", x"e8d10c3f553f536b", x"fc928b9214fb5af0", x"65f75aea915ff2a8", x"aa625321d17858c0");
            when 7599358 => data <= (x"1424051eae4b5953", x"2673e47e9647d93e", x"e96e43357b2e0d39", x"a412947cc8501d5b", x"365e1ba011bc4bd7", x"8c1aa34c5c7bb217", x"60ccd3714bf70722", x"70bb7dc12d4b33b4");
            when 3218924 => data <= (x"84279ac43a08b6cb", x"14bafeeb881cc40b", x"df6432971133c9f9", x"ca122acc224deb04", x"a1c0f58212f52b81", x"7fbe99e38eeec1bf", x"eed7e3dc25a4ee9b", x"6858b629a9319e5d");
            when 29351379 => data <= (x"a6353b5df39ebc51", x"268cc08a2618dd58", x"757a3ae5dded5566", x"064ba3604ca92cf9", x"3d69a1232d26109b", x"00bb47d94fc59af0", x"f16140da9f037298", x"ce683f8db830b912");
            when 32899296 => data <= (x"ecfba63df72bfc77", x"cd41f5daec30a04f", x"edb6a217843580da", x"d204c7d789b0c190", x"e55b67e6fd1924e4", x"778ac244478bf9dd", x"563b9675a77d2b00", x"0cbdd11ce07042de");
            when 27097806 => data <= (x"78f7f2f7b522a3e8", x"b8b3161cc48fae3b", x"9f43bb1008942d1a", x"286bdb9dc564564b", x"658d307efb2e89b2", x"e4428b56f24b000b", x"4bc09199e123c6ca", x"a1f9435003d41061");
            when 6274207 => data <= (x"a528fc36163e134c", x"715383b6eab71654", x"346f5de53d713874", x"b624820deafa5c70", x"249045121b576a97", x"be01be373481dd0e", x"83a3ac8f7fa62080", x"6062dc69c2e99a63");
            when 10173387 => data <= (x"42488d69fedbd973", x"f8ae68318e13338c", x"9a48ad20ee6134ec", x"1749d3b30dce06a6", x"e4141c26e4be11ea", x"d6bd9c9d3644ad94", x"833ac088d909595e", x"743570ad3cd23827");
            when 2939863 => data <= (x"ab2dff62401313b0", x"4a5a049d0486248e", x"9ca94bd974aeb5b3", x"6cd0f82d38363819", x"f9bcc6d3afd5b535", x"c468b3a3154d1255", x"05a6a008c6d0a88c", x"dfe36987dd5d31cf");
            when 23847303 => data <= (x"68f3d725e25c2de4", x"c2ad64127f126555", x"9298e34337c7fec9", x"a8c9e1158aac38bf", x"3bbcbb9dc2382ec2", x"a86ca0182521c444", x"3fe29d1af7320441", x"40a2c282e5fe475b");
            when 30444518 => data <= (x"6ee4ab081c058bb1", x"639a36ee48a8b68e", x"f82c407bbf439e3c", x"4856086e6d09d793", x"bade26942f0640ce", x"ab2cd753435266b6", x"af013fd22377d9c0", x"5f3c32f106ad327a");
            when 5196034 => data <= (x"1713728641f07c29", x"cbdb14041d1e806b", x"732d8179113917d4", x"26dc2c62ff37c627", x"90def67a8c5ba197", x"f1429d3028b3af49", x"ca0f088e7ca76ff0", x"2d4f1b2893a193db");
            when 5417271 => data <= (x"f625b393f65788dd", x"d18959b5e2d3e6ae", x"2e36b8a1c4d35647", x"55637e1de67fb277", x"c817d9b4f1645200", x"4f2308c7bc76b5da", x"35d2ba5e208edd44", x"ee07a5403503eb9a");
            when 4704551 => data <= (x"b4f982255334c4b6", x"33a742bbc2517615", x"79c017e422c6159e", x"092df09dcc4d7c6a", x"595388eac91c7931", x"97ea0cd00633bf43", x"d1f75927adfbc720", x"4185bb46bd153239");
            when 11506919 => data <= (x"bd4f2f2306cc3caf", x"0d213d66d2f707d2", x"428ae49d3b026437", x"2949a0df1ab3d5c1", x"671411542451b9d4", x"47cdbbd719d39ace", x"92bb595f4edc4215", x"106f79eebd684707");
            when 27080049 => data <= (x"c1e07070c878ee1d", x"c4bd8ef2fdd9a70b", x"f8ec2a98ccad2747", x"dc613be549a389f6", x"a34439a2323e505a", x"279817cb329778d3", x"743b2ce6a231f0c2", x"ff5b636a493dba19");
            when 24570935 => data <= (x"946cb0f5880f4bfa", x"9d552e32850fc039", x"dbd194e3fce94a3e", x"802c8787e7a0b8fd", x"e20ad13144d3f182", x"02c0553769aebedb", x"b77ec1c617b5ea71", x"5f351ce0e6792bc1");
            when 25782852 => data <= (x"27c7884f62bc960a", x"29083feda0535b44", x"ac8a16cb213ce13a", x"68f65bbce57dbd3f", x"ddb4ea32e5667dbf", x"29b7e17b0d6ff729", x"d8012b8734bc0642", x"92655ddc7d881164");
            when 16752332 => data <= (x"547a551874307fbb", x"7e5b7befc15ff6c3", x"83b62ab98526e2ff", x"491be69934c0365d", x"90847a8f8531c480", x"036042b270105fed", x"0c61b9815ce7976e", x"41ac3020728e64e4");
            when 23617018 => data <= (x"9a8ead6acc7f543d", x"db1cffb13b16e7ea", x"9c035a2ab799ed47", x"663488e96dc76046", x"6645c5e29df588d9", x"5116e6001801bfec", x"79e58d2cd4a25504", x"c324b9115b5d65f1");
            when 32498803 => data <= (x"25d26199f8899f17", x"d188514d76618fb0", x"1f88624f4c5868dc", x"70c1c09e660d1e7c", x"9280a1eb2e53edbf", x"2c544dcde65efb72", x"f1abc5df4fe63278", x"d52a6e13b10ace62");
            when 13767172 => data <= (x"d8fe2af9c55e8c89", x"21b53d954675e735", x"92f25c1978f1c4f7", x"17a244a91fc47404", x"26660800179a20ad", x"1f75dcc04814b244", x"1ee2ce2bf3551f94", x"9f24d76c7db9eae3");
            when 20844524 => data <= (x"9b5273c711a83b35", x"7c624e0cb95560e4", x"6f8e0da65d6ec735", x"75355b7336a1e91d", x"0d91b291ff23324f", x"b2d750506bff6475", x"ca8b0460691867a5", x"b43e16113bd498dd");
            when 5004614 => data <= (x"aed2b519505b9197", x"e71d02745d70d1e7", x"954770bec0271f66", x"67694886ed3b70f1", x"af1976b0f1519425", x"6877cd654441763b", x"86a64e9bfb8babf1", x"807216c32468a9be");
            when 13572339 => data <= (x"c3ea8365371e8f57", x"6490e626f11f9240", x"c0105a64cef6ab1d", x"bddbbd306c1543b4", x"d054ec916ab3c447", x"b4500992dc2b1cbd", x"ac64087340f8f57a", x"7b5ec84a22b66081");
            when 33553946 => data <= (x"b15e412e34696eaa", x"55cdac31815ba420", x"a3ad8261a802da17", x"c8f3e09a4bcee752", x"b9ac254b1b2961d3", x"9360a6bba472ba25", x"992ad75c3cc881e3", x"24be8363b3a10ee6");
            when 9027843 => data <= (x"e4903870044bbe4b", x"e31174a35b7875f6", x"1554f60503cfe6dc", x"ab6dc7aaacf77b57", x"64a70696a195c178", x"b90c43d3e7aa8dba", x"06da6230166d1643", x"35a46b63184f8db8");
            when 14375153 => data <= (x"e2ed8c83cf2aa78f", x"6b823b399c6d9eef", x"ff878aef0ed3835c", x"5073ca452ecc3c35", x"ba68dbbb760a0442", x"2292699afd0cdc58", x"932a8d83133c0a47", x"49c4fcb70bd8e5fe");
            when 28014258 => data <= (x"e6c7fb382b96543b", x"55adea7ef7c773c1", x"7a32c1321ae21479", x"8cb2c9ccdf3222cd", x"64b90314d230a216", x"93137323a7282e4f", x"06695d48a8445842", x"68b2e7adce4a012c");
            when 9579494 => data <= (x"e37b054b69488ea7", x"cac16f709cbac6e3", x"f5d6e21264b4969b", x"f6a234c60f0ae34d", x"f4e859d3ee5e5025", x"a7f7b373b46e7b73", x"6dc90fb22affadaf", x"2d4aa58d1bb6e406");
            when 13701525 => data <= (x"10ab6c1dcff026cc", x"dd81b760953026a2", x"b82b9394a2008fb7", x"68621a208bc0768f", x"b423193951ac6408", x"3688e0c501c8c839", x"ff4a4ee60403ed23", x"00ed49c0293fc7cc");
            when 10057665 => data <= (x"1d997cccbc1b4d86", x"4050ad1a5302e381", x"cd68550fdf28592c", x"375568f26546057d", x"e70389b87ef1ae67", x"f1def06a92bf9df5", x"8cc7b2b8df544c9f", x"9d3d0fe154576a9c");
            when 31709287 => data <= (x"7f24c5abf1fe1d68", x"2138b99389e375ac", x"5fe872051ce9ce03", x"5a8153261c05662d", x"179478dca4351fdb", x"9bf0eefed5bbe0cb", x"22ca7930925dd14d", x"25c7fe8859c9ee5f");
            when 6613448 => data <= (x"38c96ae9314431a4", x"85a0ac4646d06701", x"12e9021d8da03873", x"8cde07fa21930c87", x"d736bad5062f49a7", x"be97c77cfdd01157", x"363031ee1be16bee", x"285ec53d84976804");
            when 758832 => data <= (x"af678a1877bf74b0", x"678ab5ea89a20cc5", x"f4c091e79f89f560", x"d24e86ccef2b6fac", x"119c8562c6cab368", x"a5cc819bdfc5799a", x"b8c4c4628c87cabf", x"b8fd0ad2b8a8e672");
            when 28592429 => data <= (x"93358cf81c80d5b7", x"819ef8c29efab71c", x"985554110b5dc4bc", x"27347ad57621f1fb", x"a0e799daf22c1de8", x"ed66d24cef142565", x"47caf821a5e85240", x"dd641786c767a07b");
            when 24480425 => data <= (x"68974e9234f43fed", x"56113bf3d040f25a", x"c6dab71d13cbc28a", x"c1f6dead9d7447b3", x"13da85553897de14", x"9819cfb7b926fb09", x"f5f344a262d21281", x"c578af51d721803a");
            when 17531998 => data <= (x"fa1682a6a8efa49c", x"fdc10bd62df0d416", x"5b4577d4bd484ff7", x"9a89a898206a9e15", x"e06a468b31dca7c2", x"1817e1ef87990f6c", x"bdf1ef1614fd9b10", x"ad03bff1d10e7d29");
            when 28304149 => data <= (x"0631781c122fdbc3", x"e83f3735e7adf480", x"fd099f2518b7dd78", x"c59d75f724140e54", x"ba561809d5696697", x"8735827ad8042842", x"7efeee71c5e00f5c", x"818a72ff198635f8");
            when 12500550 => data <= (x"d2fcfabbc859556c", x"3bbd1e83e4008cd8", x"854f9602dbc7b14d", x"a4a2ea1632dac2fd", x"a2927cbd35aca73f", x"9738901b6a3e63ae", x"5819f0d79ff10f25", x"85211b81a8325d84");
            when 12444880 => data <= (x"55bcc5bd354fcc70", x"65bd2cade6c03577", x"c590163cf2749245", x"4a01c9d3f8bf0ed4", x"763aed23cb61262d", x"a0f3c80be4e2b359", x"fa17bdd4417cb8a4", x"956de8cea569a65f");
            when 29915381 => data <= (x"41d2cf8617c6ed8d", x"deeed572719dcd46", x"234209d538612d91", x"1747f202bd7bb3bd", x"12d3c6051473d2c4", x"30e62f05cdceef8f", x"90887484b23705ee", x"7070eac16d2489f1");
            when 17883987 => data <= (x"4480977416f0c711", x"48afd7b2720fd653", x"e211a39abddbde65", x"f79abc5847a8aff6", x"6460b4a61dc8969a", x"28795f99828b4e9f", x"0d34de8545360067", x"1d16ce6188d077b9");
            when 19711229 => data <= (x"336c37a00a16cafe", x"9eda1a2de72ffc82", x"7dfbfc6b371992c2", x"409681a45b1ad5db", x"b5ad1bed53b67174", x"4739e97858baaca1", x"26b4e9df95ede033", x"d92145cc0056e5ac");
            when 23906963 => data <= (x"f7c20b05147368a9", x"9f1d73e4c5e6fb06", x"81e97e1e412198f3", x"a23ee786f4e6e841", x"9cf4094b22fd0a12", x"7fca325cd1574216", x"ffe10c4b259f5e6d", x"561fac22d73b7db7");
            when 13335521 => data <= (x"011494b0685745e1", x"b39e6b298bc9948e", x"356cd2fdfcad226b", x"50fa2a4fab36547e", x"cd6fa7127f7e97f4", x"d64ecf735fe8d4c6", x"44f8e8a3c02f98e7", x"011cabc324da0afc");
            when 12362792 => data <= (x"0543ae6bc6821294", x"da2983315c0b54c1", x"87025b6e6ab828c6", x"532c17c2fafec870", x"88276586075b7efe", x"5c8fca7600357081", x"9d495fb930f05b8c", x"27370146c0ae08dc");
            when 3297116 => data <= (x"c46bb4cfff1c7a8f", x"6c7c003658ed188c", x"bce1aa2d642df421", x"c9aaec07147f7174", x"9ee3bc74a02f8973", x"9af4309707d526dd", x"d0339b8270a856cc", x"3887e72a33b0b2bc");
            when 2007462 => data <= (x"9171ba3c2d860a73", x"a456b85beeb82808", x"f65125333e2b6837", x"4451a60f5fae850a", x"a36f0135a309f895", x"953a21986975e08e", x"d6d440da89ccc63e", x"caa23481c078c911");
            when 18033055 => data <= (x"4141891316cf2b38", x"f64491d989c7dd83", x"0eeb4ff3db8321ca", x"bee16b512ffc2e37", x"f2e86f5a0464824f", x"218c1f870fe6bb43", x"8a6e4d47e0b966e1", x"b0eb9514ea36c493");
            when 24704453 => data <= (x"019e3be8ee7ad71a", x"6c23a888a44b01df", x"3d1b83cc9cac1ae7", x"1476a98832cbe2bc", x"6f529345a8e52719", x"a37ead89cbd7317b", x"42c9fe5ec5f484b5", x"ecd0f43b01321427");
            when 19176385 => data <= (x"545b6c492e3a0459", x"76f177fb1e087c37", x"f2b2bc6c6a80bf7f", x"b84d23b07d48e3da", x"f6bf5ca1fee60d7b", x"89c5d708fcf91e4c", x"4c869ca09882e62a", x"ece7ec7849ddf3da");
            when 28700173 => data <= (x"3240459873cf22cb", x"0c293538e2666c01", x"3038ade06c2869c6", x"3b2fdf5b5953f358", x"760e965847ae3971", x"460974d62ac1597f", x"f2be045f671e6cbb", x"330513087224cfa9");
            when 22022275 => data <= (x"0d5b190be411c485", x"b524daf55cdbfea4", x"ee0e3f995e519b80", x"4d1a7ac809ee25ff", x"bf6a8f93996acc14", x"4871aca742dd9548", x"35eb602f2eeda7bd", x"668766bf84321c6f");
            when 1839982 => data <= (x"a56955396af0d057", x"6db50ddd34a191eb", x"7ff9f4b0754386ab", x"0b6ac3ca2db0d521", x"9250b888655cfe2d", x"88c4a8865e1af5e3", x"080f74dd269d0483", x"daeb4f3d76200aa7");
            when 3530168 => data <= (x"41fd58d224f21eb6", x"e9f19cbffaab64ec", x"fc7c218013dd23d7", x"0563584172dfd2e7", x"3dbaec21581bcbeb", x"03dd744e44ad9201", x"faf57e40e6e4ea5c", x"4a785d05695d3097");
            when 9402596 => data <= (x"fd24b9134fbd7d05", x"47ed799f4ea0281f", x"5d35034037d7e7a1", x"2391e9c3d0580430", x"7ffd395e5d717bfb", x"818668f07b656b16", x"ec146e44b3039bda", x"d3e284f9eb7e1930");
            when 26260188 => data <= (x"df429f8a36cc5b87", x"c2fa016e82c30823", x"c0d176799671ec8e", x"30858c7515af64ba", x"687dfa00be59c236", x"fb99777607b483e6", x"a176c3d4a6ed53bc", x"25f31366f280d95e");
            when 27052890 => data <= (x"9f7b1415e8b8c850", x"4855dc859097ed25", x"43b8f63d4eb56ab4", x"49b01292e3522d59", x"4f7d7a7089e80ccb", x"cdcc544534f484de", x"a39c9a93e9df5393", x"6ccd6c713ee078ba");
            when 550987 => data <= (x"16a083e043276214", x"e69734c70a255cc6", x"2028e43dc9201d6d", x"41bf54f5e16b8704", x"abb781bbac003eef", x"66c0406be2db3680", x"b3b07de3b1f63d64", x"d99135c533f6ecf1");
            when 2251112 => data <= (x"803ba624f2b2a12f", x"704c7416c0f0f880", x"645de2188167834f", x"992c7b960ead8815", x"21d5a2fd5c8f2ff4", x"a43f1750a6d138c7", x"be66087c3702f1b2", x"1358e8d761bb4d68");
            when 16932703 => data <= (x"4dfa3b83c9eeb61a", x"d5c0f1bf9706c322", x"b395a61b77121662", x"2ad73262fed3cdcd", x"7034fc8a15b64933", x"87f71585233941e4", x"99bfc7e8e2158cc2", x"c54949bf35a744b8");
            when 23351987 => data <= (x"15d1d78f80e4ad1e", x"993ad2dbb41d37bf", x"d60d52388527e6d6", x"989bd3aa824a2b47", x"5f6fe000c2d5c985", x"d21c6a7ea15f976e", x"a899502607c544d3", x"51891c854a602889");
            when 32551038 => data <= (x"8c2546e875acc9d2", x"afdd6e6fa374d9a6", x"c55456dac965a91e", x"43ebb0a4385c50cf", x"a90e8ec116e36dfc", x"5f3fbf0e1d8ae068", x"492ec9b964012323", x"68d5265c8cf84bb6");
            when 20913358 => data <= (x"75769fb1d3132b94", x"6c66e51b53c0f226", x"5778965ac844770d", x"caca4e82b183f456", x"1441fd97b0f8e13e", x"f75282c0473c8b12", x"dd3683932d46a57d", x"40ebeb8210829c1e");
            when 15060832 => data <= (x"b130aa010391bae7", x"e077243539bd9854", x"2b3f151bf675fd8c", x"ec79f38a2234fcb3", x"de8db0e7918d7e82", x"f3f2ffe969d157a3", x"7e2e9aa9c8e6c67f", x"7ea9eae2a5175fa6");
            when 6526842 => data <= (x"cb30dab9eddf6c9e", x"c9d7c8b88973247b", x"8b7e10a8926bfd31", x"d98514cc477f82b6", x"e5de2168512e17fc", x"8bc45160dc17eaa8", x"5039c963457d1de1", x"2913232a70dd1c5c");
            when 4339999 => data <= (x"fd451d8807d969f6", x"cfc8d945a6d19ecb", x"95fadfa05af871a9", x"ea70d4d0c92b5a4a", x"dd621b0054ecdadc", x"853290d2fa3f87b3", x"2af0b4a0c2eb3694", x"37f29b453776a180");
            when 30306161 => data <= (x"51facefa79bb3ed5", x"f4c08bbc9cb4c050", x"64ed7b88c6d8cba0", x"92d29a7b03693a87", x"6868e4d83ad80c90", x"ebc22b625b9b0093", x"c2b96f84bfd1586e", x"6eee1289739c6555");
            when 27653486 => data <= (x"dace172548f5481f", x"7d9f02c8e46cdd6a", x"9bd1abb9c1f57c05", x"c8a1faf3bb25ac23", x"fb5b7683f0edd3a9", x"28347c9ab1368df6", x"f8938d19628ce58b", x"f8d7289a7b549be8");
            when 8507828 => data <= (x"2ab1367799de1c33", x"a334ae670b7d7245", x"d41e0c1020642555", x"c430228a4b9f493f", x"f02b68bc36f85e4e", x"1fe0eb77e0cc7622", x"0a6e29bc3b11bc4d", x"b5ffd1ec55a8a35b");
            when 1496831 => data <= (x"6f3a16b1809306f2", x"042ad95a36e3eed4", x"f377c658de23a941", x"6ff974331a345554", x"e2d7414301d2122a", x"e26a383eb365b178", x"54ff65d419ee44d1", x"13bd7a2df0f15e3a");
            when 12352167 => data <= (x"42d51900a05cf3a8", x"2f429098d89c5b44", x"300d3b71e8ff7953", x"cd1684d35e2226d4", x"1c3fe821c41d7627", x"d3daf52f02c79049", x"3f32763b266865a8", x"4d65b6d80392712b");
            when 23212879 => data <= (x"21a4289e5ec8688d", x"3b36f2b61a553157", x"f876c1449d3ebb78", x"110dff9c8412cf8a", x"eb4a1a635406c821", x"43266d65a7f577b7", x"47325092eb3950ab", x"e3af6179709133af");
            when 20816736 => data <= (x"4c9423c755771ada", x"88c87323b1c25145", x"52ff2258fb70a7d3", x"d158ac258d537ab6", x"234a5a1b285c9ee6", x"a40045a4ca7b1cee", x"f8a46eef42657b5e", x"9112b663c3beb421");
            when 21551502 => data <= (x"c7e6c74df9677e7f", x"9967b4847eb7d8cd", x"e8c03b82ee922d81", x"6ac18cc75a0c6cf0", x"a23a57ab37f1d2b6", x"8230fa9326a92d6c", x"d895382f42bb4ea2", x"5f4f2fe020177c06");
            when 18033133 => data <= (x"41671b141986991e", x"aded30e3cb8520ae", x"d77139af3b8ecd4f", x"8031b1c39d04731e", x"df6535c93171ea83", x"dac4bad71e6be743", x"a40253aab1cdc481", x"41e5a2909dcaddad");
            when 26600573 => data <= (x"4e5f3e035864ef8c", x"1a4031246deb675e", x"e6063f6b9a3c09b3", x"23a362e380515a02", x"53c65b1580c19cc8", x"5d49646a51b997fb", x"c503c08cf157603f", x"e9841f6ba5bad019");
            when 11960197 => data <= (x"afa1e16a162b1191", x"115088943e9bfb4a", x"d02dffc598209123", x"6961155f2b7ebf5b", x"3b2acc5437395507", x"701bef1d04d04c51", x"03a2bf7c617ebb6a", x"ae2136eb3c59970a");
            when 32595764 => data <= (x"4462f77ffd6a81d4", x"287b861e3b42128e", x"1fb3b6c3314bcec6", x"af249097f9de9c69", x"5f13fd4796e540d3", x"0e68c03370210206", x"d57762d2d5eaeae9", x"b02b30b67ac06b12");
            when 10578960 => data <= (x"93eaeebc19fe0278", x"cec3d5224eb81ce5", x"ed06b97249d0ac9c", x"aa13a2d816d6e66b", x"531231f5a26adf59", x"0485080a9aea1339", x"1c488cdf65e1b168", x"c7cf181d18323b5f");
            when 5355156 => data <= (x"fafdd50a372cb2e9", x"44dbc1c2989b5906", x"81ddbfb9abaa55e2", x"8eca9c593302f34d", x"6291732bfde46228", x"fdab42ac37701073", x"5b6ab20883dadc50", x"8238dca36498d36e");
            when 24071225 => data <= (x"b64d7eef6f663544", x"5cc453faf5ce8b74", x"fdf449b5156c8cef", x"2fa46eeeef364e05", x"87d8b16c18fa30f6", x"92d8f64a15bff6df", x"5c051fd1eb256ff8", x"1c9e548f74c9017c");
            when 32048963 => data <= (x"c76b4a1e27894228", x"4029ac3c4b00abbc", x"dd3ea2575f8b34cb", x"20d162a59915aae3", x"5f820f0ac4ee3574", x"25f78bdf37f1681a", x"652de2a639421885", x"8480284b2d9f0560");
            when 32381430 => data <= (x"7d993b49749835d3", x"1e02a2700691d2cb", x"b2eb38aaa52a8cc4", x"2c17ba50c3661da4", x"6c962030a2479eb6", x"45d679a2410b456e", x"b4c5552ab42ccea8", x"54ae5e6be9f83db4");
            when 19635002 => data <= (x"e8234fa41b3d22dd", x"5332c7534088114f", x"1af10bafd4c44339", x"8b24f23343fc0765", x"3792a484066636d6", x"e6326552cbab6355", x"6ed681049ba886ee", x"ed4b820e0aec9831");
            when 9819848 => data <= (x"f22c39b93332f28a", x"68d8a483d8e46dc0", x"d497ddbf29946969", x"64e8a595b6a6d080", x"05e3abf4b698cc05", x"7283cddd0964bc1d", x"0df2886c2dc5f502", x"019ef1f4110bb5d2");
            when 21588904 => data <= (x"988f076b788e0edb", x"19cfdb00962c8c6c", x"78c6b1f18900ac6f", x"134f1d95d08b2b49", x"3ccd4ac2ec47a8b2", x"7bead3f841e9333f", x"600fb67c89daa18d", x"6e210b983542394f");
            when 8494166 => data <= (x"ca09d69bb3f0c5f3", x"18bcf19b32612de1", x"287e382e30640bf6", x"ddaa4f6bd5227300", x"48e672b390895551", x"c52a0a6d2bfad543", x"c7f4ffc035979fed", x"91aa7ec00cdd9e64");
            when 9975186 => data <= (x"a070c715680f206f", x"162505bca2af8937", x"c4aa826f0a8c6b77", x"3ffd22d6e05f8b28", x"225b338b92e5bcbe", x"66add3ab4eb7a485", x"9b9befce37997172", x"1acb7e0d0f1a231e");
            when 5810482 => data <= (x"2963b710e7d0bef3", x"1123b74e5a436b40", x"530beb077cd6027b", x"751621420ade330c", x"ac7669e78a00c1e5", x"cbd9767493670cdc", x"f6414d2446b45578", x"96e43894cfc3ad7d");
            when 31142430 => data <= (x"c9fc069c7d0eba60", x"c0635d5f58bfaded", x"118197f744dfcb96", x"4dfe84965c4ce810", x"c4a66b0250c901dc", x"32dabbc0967db092", x"b96a6d4378b1de54", x"036336482e78ecf0");
            when 16185607 => data <= (x"bb0361e682591225", x"ee70d3a0957920e7", x"59f27a2358545765", x"74fb603544f64080", x"068abdc0ec30a087", x"1ae8cedccab9237f", x"d185999f1c296df5", x"252e9e4f4d9dc57f");
            when 20093686 => data <= (x"7c4223083e55086f", x"fdc741d4d0a19821", x"db8715e915b62f4b", x"fe0a669a2b388e17", x"f00d117bdcee778d", x"552d1536567a6526", x"3597063fa446764b", x"85d85f18c14991ae");
            when 17247504 => data <= (x"31b72d56482d9efc", x"f6370249c273b0d6", x"a94d018bda0615b8", x"5d893f19ff299728", x"6db15d44e096a526", x"6bbd26e279cf197e", x"a84ed1eb50e50e58", x"a3ec68b7a76ac63b");
            when 15727202 => data <= (x"594f9db114b2380d", x"b4c547e9788a859d", x"021a896f2e9f7777", x"02f77f581c38639c", x"6099523f272f1425", x"e026de015d837199", x"2ce42edc9b4a9592", x"f34b5387e5d5df82");
            when 24310249 => data <= (x"817723c978859eb5", x"351fca7b7ecf7b5c", x"23b3ad8d0693ebfa", x"a4810308c124b640", x"e0e9dfbad038a151", x"58c957e2972cf9e9", x"2c92399d12d91c21", x"ef3a5a6c6418e5e4");
            when 24580696 => data <= (x"4eb97ca8896b77f6", x"7e00723f64a1f7d4", x"1c0a4fba8ad0ba76", x"6bae8a1ee8c9e71c", x"625f7ef10de1ca7d", x"b9e38d2bdec8a88e", x"84c6814e9e661666", x"01ca15d58aa455c7");
            when 31595475 => data <= (x"a1078df885bebbfd", x"d60da14344e4394c", x"3bc248205c73204e", x"b085a7d650e9b1fe", x"627db12591856f38", x"4a17a31936d3d049", x"91377b80fe8251f9", x"d2385e135c7f68d0");
            when 17447900 => data <= (x"2b3c932fe1fa460e", x"1bdaecfb65e9b0e5", x"d77ac9b512e044ac", x"b1be5c5530d1ace8", x"47acbc277b9b4f48", x"6ce1f6e5ec960077", x"c31689e6e385d2f8", x"9c2b8bafc69b1a66");
            when 32089248 => data <= (x"031a69d3f44de36b", x"2185c7589e8b6644", x"080efd7e95f8d1ea", x"7da963f016fcfcd0", x"dcb572dbb5aab1c5", x"0717cf7748d84869", x"115499e50f746502", x"4ea5ab310777ed64");
            when 14291855 => data <= (x"515b026d6269f572", x"16efe43b585983c0", x"9c29da9486025a68", x"2fb1429c5b52b334", x"16859b28c454b784", x"f7a6d5476c3e149b", x"a016cb01c011e4a6", x"80b4fb1c14b4fe25");
            when 8825579 => data <= (x"6163ebd781090471", x"130b86e7c8e58dc0", x"84dbebc7636f2f5d", x"a92d7a87115bb0e3", x"2444b02be29a1df4", x"38f9b27ed552695a", x"0ed329cc2a218d91", x"83015a158f345ce5");
            when 27220364 => data <= (x"5bc8276f432641c5", x"835495e7bff1765e", x"3d4f24f0b5eaf1e4", x"96da4058f0500dbc", x"a85abc49d63a4183", x"e4c46f2d2f8d15c6", x"4e29b6098c1c9fc5", x"c5ac74eaeb64cf41");
            when 16247226 => data <= (x"3c855905b0ec07da", x"806b01c794487170", x"1c4d1e0cd6d93c48", x"5a966719815e0e76", x"c8117f6514a8317d", x"d93099896646c2bd", x"e68d4c08c1fa3564", x"704763b406ff4b6e");
            when 8897544 => data <= (x"661aecaa2d785ff8", x"12b6c03927d88173", x"b6e3c95da0c3f4e7", x"33cc5f6b4c262734", x"ae423ad293fc90b6", x"da7b73d89372d413", x"e94cc72ebd73094a", x"86ebee60fc518f41");
            when 24236819 => data <= (x"3a966fbad61d5ae5", x"9cd05a11eb2c7007", x"4d4b6d11bb8d2950", x"b9cdcc1d407f01cc", x"a44a121346c1dd9d", x"af9ddd1ec6a32bb6", x"2436cbe284a936a2", x"83b7c1102e711326");
            when 5099151 => data <= (x"1ef2eb7b7e1f3310", x"bc82c25144153f1f", x"26609e16ddc456b8", x"f68e6f97ede1b931", x"09baf6fbe66012f2", x"58efe8797528fb10", x"fae739c599406016", x"b02617d933661afa");
            when 9861705 => data <= (x"89f8501d17d4a101", x"027ddf4812dcab3b", x"45e52498d35bae92", x"c9dddd67352eb4b6", x"ed0a658c5cadd768", x"fe05367d7a286077", x"0cb9e5f828deb807", x"028ad0147898d62c");
            when 19303339 => data <= (x"e3ab86c981416383", x"7b34cda199621c09", x"b5a0e20d42f76842", x"7efdc2faebbf9f25", x"c43368acb5fcff27", x"871ef8b468625eba", x"bcf4c83356602a1f", x"3cf54a4da84b6a67");
            when 24844815 => data <= (x"597ef20e06882285", x"4b5f1b7079a26205", x"a0266fb470f084cc", x"83e4f8a0815706ce", x"cad0409929fecdbb", x"744b6a85964683fd", x"f0c6f4c9cde2c250", x"15b26d808f37c6e2");
            when 30168977 => data <= (x"c03518ebad8b6a4c", x"4665293164c87857", x"40f0ae892bd0cb80", x"ba052cfdb6b92024", x"2229864178b51342", x"69552bbb683ed1a0", x"56c2112cb9d9c9a9", x"eed6587d016d9723");
            when 1418943 => data <= (x"6df1b270101de3ac", x"d2bba25660a974a7", x"09623e9abaab1cdb", x"4e502fe88a64642d", x"545aa597a2899b77", x"4b7ddef5e3c45b00", x"d63ca86120b83be5", x"662e00035efa20ec");
            when 14550533 => data <= (x"ee82daf69b3427d9", x"9b624a1a292d44d4", x"92b158227e09d2ca", x"d9aeea865edc4c23", x"7000f36c00da2133", x"ef14ee5a14b48cb4", x"98ad0eb959a73ae0", x"2983d899dd7dafd8");
            when 18572219 => data <= (x"7b224e67be7c1ad9", x"c33245c8f5711de1", x"1295d12657cfffb4", x"0ff6e6bf0fb95cef", x"ed2ea7b7ef9ec308", x"0af7e8374908ada2", x"4c4288b773b8efcd", x"c96beeabfd2e9163");
            when 17691223 => data <= (x"caa3d47d1bad9f33", x"274306e7e9685d16", x"825dab1c7b0183de", x"b9dff33995aff905", x"dffbbcf962dc6373", x"270aa00cc762340d", x"1e868d9028a29119", x"236927c05c8fa806");
            when 13580999 => data <= (x"fd208e9fb7770efb", x"a007754903fea7a6", x"1a5e30fd653241e3", x"37c71c4839647acb", x"5f08478ba2edd25b", x"543787eed07d5cc8", x"8ce4e70ef6a9bd2d", x"35c77a069eab2ebe");
            when 17603173 => data <= (x"a8c4ada0abb37894", x"5ade6b83ef9508e7", x"1947fef16a06c53f", x"ec81c5f9f5686d6a", x"1078fd5d788853b2", x"294f6ab8a24503f6", x"f0c8e78ec28f1663", x"44acd30a4271cfc7");
            when 16402429 => data <= (x"5e61b1255472852d", x"4ce56b09ee2b0bea", x"c78d4db3d3b73091", x"ed8e443d085fc845", x"881db84fec3f849b", x"a118cf80b8942808", x"b686afb2a83600b3", x"4412f0786ddea8ec");
            when 29057022 => data <= (x"17c9328140564951", x"52e57bdc3a2e502a", x"ef9f86d69f702440", x"c288637b962fa3f7", x"80b2b3cf689d0058", x"e2fe78976211ab0e", x"3e038ff91bec7500", x"d04fe0e4e354de42");
            when 6478372 => data <= (x"cb845546fdf54bc9", x"46ccf27f908bb9af", x"6e396f497301057d", x"843912c50486d432", x"869392eb9ef25c3e", x"f00cc3b31cf76caa", x"4f12e25f5bbc419e", x"acf966e7297f7ed2");
            when 32244518 => data <= (x"2cc714c71eb8e573", x"3afa82af25c44195", x"dfa5f75a677097e9", x"d818ccccba13bdd0", x"41be86f772cb4712", x"1f4bc6a5c7602343", x"2ce37d2545d2b525", x"56f2087e3624f7a6");
            when 30596756 => data <= (x"d1d9df9ab23d2489", x"8e47718ca7078004", x"19beb38fb0398871", x"9bd698bba7588911", x"10109bd6e17f43fd", x"7aa1dac582850804", x"3927c2cdd3ca47b3", x"429ba08ba719111e");
            when 22659298 => data <= (x"183a2c7a534e8c22", x"2ffb64a56e9cd363", x"3fabd33f3237f5a4", x"f5c808ea79bc3c16", x"79073bbf5e2966d1", x"52fd9f72f2f6acf3", x"58496e9d53a15fe7", x"95f5a6edfb209cfb");
            when 31097365 => data <= (x"bb0d0f6d4651adc2", x"4f5bfc4784d75974", x"f7634f8ffef50f70", x"f99f74b87ee5dad7", x"e5dedf19b4713fdf", x"e133b21f31e48015", x"27b367e0ba793947", x"8fd81715f7d5d348");
            when 12214792 => data <= (x"4a45727044144169", x"a9b657bedbd10de9", x"766f0b70e48aba4c", x"bd7a29aadbb7187c", x"fe19b572b208f8d2", x"10a417c8d9ab0c79", x"ae40e518271c9608", x"a41fa36b6e9bda60");
            when 5761601 => data <= (x"d8971f484be5fd8d", x"07543fa55ec5e58e", x"823f042ecda8ed7d", x"08a0b8cfedfcadbf", x"eeda71993de79b47", x"ccb95629c1a0000a", x"b95501f0082be110", x"31e81f6d4a86f3d5");
            when 14451215 => data <= (x"48bd9e922fb9b372", x"7977484e3fbab559", x"aae399fb4df8092b", x"a19dccd3f7f982af", x"526dc8c587df73c8", x"23bf21f49ba9d213", x"0bcfbdf7e926eacc", x"96dd80ea954ed159");
            when 13546087 => data <= (x"152ee03f96010e28", x"b45269f11fc1fb59", x"cd8f1513731f5d46", x"8efab3dc42e4663b", x"43615c3db5b1d5dc", x"bf0f75c7f9c06b82", x"70e3d73beb976a42", x"d8072db1891b1efa");
            when 4844252 => data <= (x"10c3d60d75834af8", x"ec1e9d147eb33c0a", x"7dd2c734cbd94c40", x"f5cd18078780887c", x"97410e9be36f6a05", x"d4a5b6e6703f6148", x"ca1ab4af877cd680", x"5a14afb8235ecf73");
            when 7414747 => data <= (x"8aac888f06b57728", x"fba69a5d15ef258b", x"7b58cb8bafcd00e3", x"671ddf2bc8be33af", x"086432956925c1a1", x"a29d82eb0e63c3bc", x"507ce5603a384a7d", x"5a20bb8f54a36595");
            when 28679558 => data <= (x"65c7aefe3a156525", x"5f9f34028103b43f", x"61895259e241a9f0", x"3eae9fcd373dee0b", x"0832113b34d4fb05", x"43cc0dc508843bb0", x"003615d1ebc03070", x"535af2148b059927");
            when 470483 => data <= (x"56bdaeda7ac4fc49", x"47da17b9cbd2a633", x"bc8eecce30e2de4c", x"68a0ed2fb30c249d", x"601a4686b2ff8011", x"b49a492d78c826e5", x"4f19186934b5c409", x"b79c775b5269f473");
            when 23559427 => data <= (x"067ef4caaabc07a0", x"ed469f6cb73378ce", x"f533363fc144bde8", x"34a71009119ec911", x"ed49e8092ee8e4c2", x"7e456e2a744b2a6a", x"04d6418da0329d11", x"b9509a6b1b411d9d");
            when 28337126 => data <= (x"9b2dfcf16bd0f0b2", x"b61beb0296c212c1", x"60dc0742207473ff", x"528610d238900cfd", x"5b1d5a60df50e0c5", x"d135f34cd3aaa0e6", x"e211fdbd0c76876b", x"6eecc5434a4c006b");
            when 10570392 => data <= (x"fb59ab07b98813eb", x"eae75fa060e6c270", x"cbf88ff9d8d28f9e", x"1b8d173762b14e5f", x"9065652af6bcc9b8", x"3964d4f299bb57e7", x"16644b68007454f4", x"5375c5b3140a7be7");
            when 14587581 => data <= (x"0f4eed75e7658236", x"a54bd87e7926e11e", x"6296ddd0d13216c2", x"d92b0cc5d61eaff6", x"96b15d668712be72", x"5dc93947571cd28e", x"7d8f513b39a1a62b", x"c3d5faa19e2c3411");
            when 24043886 => data <= (x"a547968c61ce026e", x"f9fb938d224f2f77", x"1cddf1e30f97313c", x"c6e7b72a29205020", x"8a6c52820e2040d4", x"163dd117a49bc14a", x"c852c74c5eb19f92", x"80dd7d83030ef071");
            when 32575471 => data <= (x"e0ab2a2822259f47", x"5a6351ca1385cf55", x"5e5694509587add5", x"ab42bd94cfffa539", x"7734c0b309f0eca2", x"f4c882fa94757574", x"61a7e8126aceaee9", x"4643e0d5f9e2ddde");
            when 28092636 => data <= (x"b8765a0b172fc3ae", x"c7bec0140af492d1", x"8cfdefcbbfbff9d7", x"52f79dab2b22531e", x"b3d6ff1f71de6b00", x"5ae7c2042ad3af84", x"93a797d8ed0a3dc1", x"22e0469dc6c93a62");
            when 9233618 => data <= (x"a020d8c9db3d9cd0", x"8da60c9ab64d0c89", x"be3e81f64a1003c5", x"8f430e66825941c3", x"21c3142a53356e06", x"8b09b28b46835fb0", x"e0d8d2c0b419c74c", x"0eee0391cf3716cd");
            when 4805775 => data <= (x"df3c9d74fca56092", x"909cbe68ee0a1f72", x"283efc0fe8f97447", x"ebdf5a7c84178df9", x"cfc123c5487a3e08", x"52a81123401e1454", x"f46ea1139501fe70", x"17b3f8dc340f8e42");
            when 7514125 => data <= (x"30802920f9e4770a", x"c53c8ba312022ed3", x"60a5ae4780136913", x"ab786823c6e11ac8", x"647218af9e19904d", x"4ce7991f69f451a1", x"f45f8df8d7c7eec0", x"8656cd17c1ffb491");
            when 23819412 => data <= (x"36e39c89fc162963", x"e3a0f7b062e0209a", x"ae871b1a7f71851e", x"9922ac9789e87721", x"2eece6b6ef3b8794", x"4d4bac77d990f37b", x"9dca0cbc7fab6d0f", x"59cbc487ee46b4b1");
            when 18065685 => data <= (x"85348a9275225a25", x"cec8c7a39fa7a74e", x"26a268330674db05", x"b580a1a23b642792", x"cc5e7bb48e90dd99", x"86a8f8b07e0d7b8b", x"3ab1d43126f7fbdb", x"ac0651a298d2afbd");
            when 24275065 => data <= (x"331385dc6b88998a", x"feca8edfbf9e3950", x"7089b9dbf3839f94", x"85a369d61be15910", x"97883b4e3f07cdb4", x"71429c6866584df0", x"8b047881f71855c5", x"86a63241542c51d4");
            when 2507122 => data <= (x"cd863386ec02f363", x"90cef4d6563d542b", x"650bedb9db4c25b0", x"47a5d324f53f1085", x"a750a3ba6b559a56", x"bccbde2e0b43e80b", x"b0a68f5d07a27f98", x"9fdcc9446a5062fd");
            when 16587773 => data <= (x"1c731b9c16c3cbf5", x"5e7fd86be24e6a6b", x"3c9a94c4f8ce8605", x"876255f1642ae679", x"953d4937882f11bf", x"0ed55338c679f4c7", x"b4d7e0777c596728", x"710e86eb70052773");
            when 29681599 => data <= (x"90a79afcf46b6dd1", x"134b70756ad94453", x"89691da8eb68b354", x"8901fc5824c72cfa", x"f92d767902f14f08", x"8f83284d3b4ca443", x"b522062f92fbbf38", x"e7a1c56b7876604d");
            when 28094972 => data <= (x"16c5a125e9a74e4e", x"d87edeeca711c26e", x"2b45b54c748b03a1", x"7dad748eef0ca70f", x"c930b33ec6ce362a", x"ba928c1fee29e333", x"e1ce5a7cdb27de70", x"2be767c1b5937f68");
            when 8803411 => data <= (x"b8beeeb536dacb78", x"eba8810dfb4b4433", x"316b4eacfe074eec", x"458464e5712f28ac", x"364e5a0a5c635fbc", x"aba2f355451c3d43", x"3711f32e88f3b015", x"4e1a25fcca19bde4");
            when 8432199 => data <= (x"0df025dd1aa83546", x"5fd3f339cfcda0dd", x"552f75e74c47b8db", x"35a8848581866895", x"ec0555ed460e7edd", x"f34b930c639aceab", x"0b359a14a5cbce95", x"1bcafa3b3591d3ab");
            when 5077020 => data <= (x"c08c4e1e99bc932d", x"e30329c9d49db024", x"3d93401b683c309b", x"d03d4f7e2297c853", x"5a79b81808bb6af6", x"6f449f5c3cd2c810", x"6004ca5c87a18ccd", x"79f44013f71a7eb4");
            when 2704149 => data <= (x"7a7367d003e3fd46", x"e93fbfaab349128f", x"2209ebec7c312327", x"09567964a70317ae", x"da382b4bce5574e1", x"2aae94959502694a", x"12ff147866e894ba", x"66e4515409429bf3");
            when 28796474 => data <= (x"eb9c728398e55418", x"06018c9901df4691", x"e179bcc4e9b4fac1", x"821bc67947ae2f6a", x"1849d1144a09312c", x"3ac61748215bd864", x"7f8c3565fa546d5c", x"7afdefeb01b0ef32");
            when 30530492 => data <= (x"d7d85bbbf6e08930", x"abe7c63afd72ac76", x"1fae97be79aa6616", x"adbc19a78df00613", x"df3e3039ef92714a", x"427cf80eb8daee62", x"b4fdee39adffd59e", x"cc8fe6a311a1196f");
            when 2888505 => data <= (x"179c00585b2899cf", x"079553a522762cb2", x"831c64e5e3ad7723", x"ffa4d6381811d18f", x"529c85990e4427ac", x"21c9d2d4a0187ea8", x"7b0707b9e629ddb9", x"d2e9c18737d89064");
            when 15458306 => data <= (x"4d2ca07221326179", x"0297f9d8ec75ceb6", x"d152d633cfa4c516", x"72efbad3d71166f2", x"5cd95d6c1fe1ede1", x"6c9cb35b64ba321d", x"c59f64d2a4475893", x"0f333be418d6f255");
            when 5361672 => data <= (x"dd40f060d812827d", x"ebaf8b1214d10c45", x"f023111564e15fbb", x"72c92652bab9f2d3", x"376d505f5bf90364", x"e99c818526c55db0", x"23d8078dc8b70fc8", x"58a5cc0250ff5620");
            when 31304783 => data <= (x"7425e529eca00edd", x"960e10c283bff51c", x"033dd812d0ce4f86", x"05aa955d7c179d1b", x"1496325a63b3f0c7", x"8edfa17622acdb20", x"edb113015ea62790", x"92bbd0c364da5be9");
            when 3657858 => data <= (x"a6d4fb0cd4f58e89", x"34671605a691637f", x"3331d4e1efc09298", x"510b9e2ead6dcf35", x"c76373421093fcb7", x"e597baf4f70fb77b", x"847513fd177cfdf9", x"8334cf47a22d9661");
            when 2101108 => data <= (x"e78e155490dd7bb8", x"afb785fa37f020af", x"eb5b3437c296740a", x"490830b61a18a8f6", x"72aac64857898cae", x"cd1036efc4387ef9", x"15cb17be62bdebb7", x"c337cc55bdf3593a");
            when 8507294 => data <= (x"447dd7f402529aec", x"6daceaec9f7744e3", x"286122c0cb70c003", x"3214bc2902d8683e", x"81732c10b4261860", x"d1832ae3582022e3", x"64eda6566cc5d3c6", x"d13eb3aeee6b1f36");
            when 32402046 => data <= (x"ffa9bde0000ad9da", x"80492a482f1fcc59", x"563970057c25cb49", x"b91c196f61e21211", x"dba3c20030791bac", x"9c95865a4bd4fafd", x"d10fee0383932719", x"895f9c6bd79dba21");
            when 10701597 => data <= (x"0195b77d20eae9b6", x"178a1827ff81906e", x"ec6867ce696bf3a3", x"60270e0eb3869bd6", x"43eb27abbc840aff", x"005d5dcf8539338f", x"b8cc77aa343a1f56", x"540aa6c355762210");
            when 13820367 => data <= (x"439edaa7737b0a7a", x"72ca02dc6c0989d2", x"f582c9d1ab3308bd", x"29099240f858c912", x"b2110b413749f53e", x"dc2ebcdadd6504aa", x"4e8ae26e0571b4fe", x"d291eb5b3f541c29");
            when 8376560 => data <= (x"cfc215de0efea10f", x"0ca8a0db92d11d34", x"0b3e29d95b3b4da6", x"19aa579be5e67045", x"759be84255499532", x"258db19ee2d1ade4", x"0dd6f4f67b8bd8f9", x"6a5387bb1ab8db2d");
            when 33554658 => data <= (x"ad4782cb5fa2a74e", x"e61c032bd602a686", x"19169fcc68a74147", x"411f9e76363203aa", x"c3c2d786915fdc1e", x"1b13b0768b93eeba", x"6444e499aac4b0dd", x"7916dc678b8206a4");
            when 27819241 => data <= (x"b327a76a049b94b1", x"e64cd4165ff18643", x"1a479e96c00a49a8", x"b5f7cc5f7e4db4bc", x"d110bf89ad1c92bf", x"469a6ea09e514c16", x"47d34e0b7adec074", x"362d0f3c0c8e6d3d");
            when 17032315 => data <= (x"5f6946751e49d790", x"f331c6274426b6ca", x"c87eb127f4e3ec17", x"b3d9bf04ad9a7bb7", x"8d821a58ff98a61f", x"7961213b0f0d5be1", x"ec618fd6d292a10f", x"5c1bea58e00575cb");
            when 11756162 => data <= (x"c45be1b3b180bd50", x"817ad83dd9c4a565", x"bcdca21908b3943c", x"748963a4f9d2b1ab", x"c472af2b880d804f", x"b8bd36e755d924b3", x"1c1338e472d3863e", x"3f86f8506768ea99");
            when 10864377 => data <= (x"ec78b81142aef288", x"7986883006d4ce47", x"7435eae57a4858c8", x"f9221e7859a6ab51", x"48aa89a00e1c5019", x"dd710af0f8206a82", x"4f78fede5662bef9", x"17603308ab832b3c");
            when 3140314 => data <= (x"2daa96d06a0e77a4", x"ef943ed48284562f", x"37690b4a8f95ca60", x"aa7519acadd2c5a2", x"3accf21e21500eed", x"311d4ed9053b62a4", x"b184119674756740", x"1440c1338112842f");
            when 3729758 => data <= (x"1324eb1b19a7ae1b", x"de229e68e64afc33", x"078fbba4309310a8", x"1f751a730f8fff1d", x"e7b09bc3edb23bf0", x"d3efcbb3b867561b", x"dfb62676838f3bd9", x"5273ccea6dc6a343");
            when 27690262 => data <= (x"7d0e87fd0841c262", x"2836e1f984077038", x"29cc8e662da36213", x"5c16e6747ad1450d", x"271c7097a562134a", x"f5b84250f3bbf026", x"a618398ec2d0818f", x"8ec033b2e59df5ef");
            when 5488947 => data <= (x"51d7aa2989cd1bed", x"ce22251c4bc2223f", x"86ae018980132a79", x"2663891dd4404574", x"bbd9cf76baa398ef", x"c3a22a7eef63722f", x"a968ace07b8d7ecb", x"5194c2e80e1ccb71");
            when 30408759 => data <= (x"1bced5cf8b7aa996", x"b1ebaabf9cba2ad7", x"e11c87b6e689c7b4", x"856ecafa708822f4", x"7a329421f2c37e09", x"0b881febd13680dc", x"9bd574d499c81130", x"85e032877d2cec22");
            when 2217728 => data <= (x"f0b0d89c248afa72", x"93ac20aa668ed4aa", x"e5bba67b2edf679e", x"0275efc4deb240ee", x"61c6768eb24eb8da", x"3e50eb658bcaea44", x"9277713c0e27c6bd", x"bf4b40c574c88005");
            when 573736 => data <= (x"7dc42fd07d8ccdf2", x"a30f1832f50bd697", x"795a64274ca13b92", x"0775982caeb34a83", x"4bd480929bc27d8e", x"467243237af46242", x"0ecff5bf1fb07d5e", x"999d74f3c1181d53");
            when 26763393 => data <= (x"3575e0bb63881919", x"c29f5944b73b9a81", x"9d94b2f674b84e5e", x"43202cd5fa250329", x"1066c6caf9386675", x"85b5ff1209200a1e", x"def4facb4ba466ef", x"361770b28e35dc65");
            when 6115544 => data <= (x"bad8bc09c6af3b2c", x"723b8a996df48ae5", x"e2ce573512beaa09", x"75236a0035d2e775", x"b20e6aa6eac0ebde", x"a63d3d3dfaed6bb1", x"f2e774b27156edc6", x"c4cdbac1fdf6d46d");
            when 15876887 => data <= (x"a26787a0864fb7a4", x"72eb3b74c818fdd8", x"031ab01311fcf80c", x"d4216c852dc89242", x"0c55b77c12bb4534", x"ec5a56c3058d40bf", x"f440c0f6b87bae40", x"d8940d7bbf50d8d3");
            when 9800324 => data <= (x"9a5a9f7f6dd8a792", x"a39468bfaccad100", x"cd6d00a21c035c9d", x"1843c79347a9815c", x"90d9d04a4001b84f", x"1bbb48541ffb6f0e", x"2bb6a8adc0833b5a", x"a111df9d11babb40");
            when 31364905 => data <= (x"3ad0e2910ea3b2ec", x"53e06343bf90c917", x"f259b8125695bc55", x"fcd192dbc19a69bd", x"50a7ac06c9e8dcf4", x"30cb66e23d67149f", x"0404d08078925eee", x"9ab669817fca93ea");
            when 25171408 => data <= (x"14f0a0c440c70d36", x"366d498981f30271", x"81e9644e089a16b0", x"bdab151935ad34f6", x"bd8d5185f028ad3a", x"78a345ab5ca05e2f", x"23832dca24c9e7d4", x"6911e6cb9aeaa5dd");
            when 7227160 => data <= (x"a8c2103393630da4", x"abf07b9806298b9a", x"21f1361004243cf2", x"d72d3ebcdb92e99a", x"ae18ea85b9aa4059", x"d60c8cb1e97c0102", x"2a01bc1d4ddfc6b6", x"6715a0cd19dbc572");
            when 10413489 => data <= (x"8009813400eccaab", x"09acb2d965101b53", x"17c8db1d35468e89", x"42eab62acf2550c6", x"c6f252fadaceded7", x"8cd3bccc94d8083f", x"6144bda770815696", x"acf1fd44074241ce");
            when 6553093 => data <= (x"95ff096db0fb6fbd", x"b0c5be9cf306fd8f", x"3dc5bef243aa919b", x"84e47208b333e6c7", x"48d8260d5f3f6fdb", x"ae362777ee7bf136", x"727cfb99fd39f682", x"db6c0b49a294df25");
            when 9442556 => data <= (x"de81ef889d46b81f", x"4cd5df64892a417e", x"e0ea696054b26556", x"c48db20720777f6b", x"7d827e7d821edb39", x"4b34535e37ec5355", x"2088385c03c3506d", x"377599008e3b7e6d");
            when 6468537 => data <= (x"56fab568b085b269", x"ca2702e8cfc1a99f", x"d6c8e18ed823b3cf", x"a3ee95190757ef86", x"0ca8346cf8b9c6b6", x"65137b8271a0d7d8", x"d85ccb3e4d148ea5", x"0e0e80a1a69ffee7");
            when 18265054 => data <= (x"f5765514dcf93755", x"7916f9d0ee1aab2e", x"5076c7663e64f950", x"501171c6c3549255", x"7bdbe864c048325d", x"2ad3d74d18bab717", x"54ef9b3284358f80", x"169bf53626817539");
            when 31817765 => data <= (x"7c603d5bf3f8de1b", x"694e6e6a3a9cbdd2", x"9cb54fca47c2c538", x"0ac4b8abc1c45331", x"47135557b06c40b2", x"27eb00dd39f8da36", x"256e5aebbe2d9b67", x"1c0c9f364b2246bc");
            when 22304876 => data <= (x"2126fa7dc0820d66", x"f7e0f39c1e1876eb", x"aaec526925120577", x"5d716a35209e5cd8", x"cd949b80a871ee55", x"13ac32e68f2855be", x"19eadbf5f34957fb", x"09c18a74fb724d74");
            when 4737116 => data <= (x"b51142d72f224aae", x"f47df207bb169da1", x"53ce85c0be8ab127", x"90cbb41f377ec4ba", x"d2fcda7357f49145", x"3a76c2c02621a570", x"aeaed17489d2deae", x"874ad759a7ee1ce2");
            when 15491913 => data <= (x"7017e7cab7d78ecd", x"bcfef3dcf718813c", x"a07e93282b9d5e34", x"07efd7bb5fecf5fd", x"c0dfbcc7588977f9", x"306d6170695edf0f", x"e387ed67d6070401", x"4e7f3fa14825ffd8");
            when 6138866 => data <= (x"a01e28725c4284b3", x"2e190712d569762c", x"0c26a9f6738d32d7", x"51433e13e17e6ad6", x"8afb5035d5273335", x"64518e2e219ea683", x"c53aa00d04df2fca", x"76fc1a1214b5ccf7");
            when 16312011 => data <= (x"361f167d890316a1", x"6d973ea1e5a06f19", x"f0692e552c228159", x"f1989ea9105c1890", x"77f86eb887ee4038", x"f3dca5f92328e813", x"4fef10c488ee83c8", x"dd2f1add186f610e");
            when 4443046 => data <= (x"ad9d0d4afc2f5e8c", x"ccad88285f9f5f65", x"bfbc9fb79a0e3536", x"6a2b222ab8b90621", x"e172615df6cc78b2", x"e709a071c183ae36", x"61b63c4761791786", x"b718428992d54a5d");
            when 4899985 => data <= (x"6892265e872152ba", x"451bd31252d73e4f", x"3de059f8644198d0", x"982c3b1055051b36", x"688e4455cdee6a61", x"bfd2f9764b2b1334", x"04fba836d0e56772", x"bddfb62d6e2aed4c");
            when 19120002 => data <= (x"ec964a380c79e62f", x"6af841aac42e46b6", x"7f4f6052046eec09", x"cc235d9d50aee2a8", x"1abc95351e6c8080", x"1d8b80e4d3aba65c", x"59804b04ba9e1a53", x"dd328c315fe89ac0");
            when 5661493 => data <= (x"97e272c018a1b8c7", x"615e764e0bf6cb74", x"c95a93867299ac8f", x"0831637b29540249", x"f2b18430605da654", x"742eb77056fb4a6c", x"9a70f7b787071303", x"55aec7f7271e74ac");
            when 19034072 => data <= (x"17b9aac397e40a42", x"bc91b893fbd2f8e7", x"0865351cdff63fb7", x"fd73cd741ffe482a", x"629d3e78937a8802", x"66264c2c9d27b9e4", x"e279145698ae4006", x"d9ed8b2b43f567c8");
            when 24727573 => data <= (x"78b43af14185323b", x"c6651c376a00c5bf", x"ad317451c721931c", x"df99569ba3687da6", x"7384f395835860c9", x"57a153ad73894b09", x"9788f1e9a17693f5", x"efd18989004d0f72");
            when 7853563 => data <= (x"db5c33ac3ab4d9be", x"ff41581720c93a85", x"653142b449004189", x"8869e29439c4a4a6", x"090d3ae568ef19b9", x"c8d5a6df6849c779", x"18ff7366ecfd040b", x"cce9271a47444f80");
            when 373645 => data <= (x"f318972db9cae09f", x"5f6bc6527fe4a668", x"6da9cf11ba35d4bf", x"7c0815c6614f7c6e", x"45b75dbdd4ccb26b", x"6d555c913c97b97e", x"a9004781dc3a5e53", x"d2fe6d45947ad448");
            when 18963138 => data <= (x"1c34d0a52b7fa159", x"246f34d0e9f7a793", x"1d4f5d812d1863e3", x"7df64e1532a62365", x"f840d54b992fc073", x"d01436eeaae7bf4a", x"f65980984b99ae34", x"605ece52c96c57ce");
            when 29147249 => data <= (x"c5156242b334c72e", x"8992d0e89f7ae3d9", x"1ead10cf1de82a7a", x"b6a1aa96b74d66ef", x"8b088f8818cd50fc", x"045845d604d7d9a0", x"20a96ee458e568c6", x"0eb68b7851a41bb9");
            when 15698039 => data <= (x"7cb133b5f875ee12", x"d5e6c4e8c8b4920d", x"01990306f1344e0d", x"95953583b06e819f", x"683dc0a418e50c96", x"f8920370fde71f33", x"768e0d5518b6d3bf", x"8721695a93c9b033");
            when 4923555 => data <= (x"95158793f7c7e92a", x"fe8e477d40ed3162", x"a7f08da3ae358ed3", x"29502456ce7e88df", x"2346d6b3df16cd17", x"7895409fa72e84db", x"8e849aa160cd5148", x"08b10c607f39e83b");
            when 28780516 => data <= (x"5c2a0ccbfb323974", x"95e2666c44342d7d", x"6b0bf3af36367665", x"17c7473128191668", x"7253b5abc38f6d33", x"950ead0a1b673cbc", x"95b7a061cf9051e2", x"93299cad3581f80b");
            when 5465355 => data <= (x"047380f3d2f3e30f", x"6e00a10204e3c175", x"d8337cfd38a728df", x"f92c21aa5e3f0a1d", x"1c3f429e1e7c6574", x"234ab818bf537695", x"94480c3e676489ce", x"b87c11460e786387");
            when 31464422 => data <= (x"8d01316a3f3aa991", x"e776c0413de50062", x"fb20cb8defe9e351", x"f8c29022a8c31814", x"a15c1f618cc972a4", x"e1ffc71710cb6445", x"ac57d63a17272d97", x"f43388b52bfe187d");
            when 32562602 => data <= (x"34d3d23ef9de20ec", x"b8451ccb7436251b", x"509b8e37a518bd1a", x"5a1d585b1f021b76", x"faea51edc3149e14", x"e600d3702aac9bea", x"4f7a6793a3ca47c1", x"65d879e239d8c9e6");
            when 9050029 => data <= (x"ca4ade26d2d82f73", x"c827e29dcfacdb3b", x"701f0ccca0e146e8", x"97951555082bf0f9", x"9784ae822ea7c0af", x"2529d4b1aa5d2943", x"539a3ba1852f62dc", x"06132652ce672015");
            when 5389993 => data <= (x"78acb11e1b0eaf9c", x"34bb51d277c4d103", x"b953b91f73c62086", x"b31753dba576540e", x"0b0a32c86a0ad346", x"fac8fafe005495d1", x"02f0f34594632f58", x"e0cfddd583153a25");
            when 18788468 => data <= (x"7b10fc22e9919b80", x"95ff55e6e2850e83", x"ee67ac7fe3e849ea", x"9cad0a8b255632ee", x"1933ef9fc150b785", x"71fe4701f1246793", x"380fdb080e06cd71", x"d6f8f90e5217bf92");
            when 20331336 => data <= (x"825a34a50758c0b8", x"ab1c4b7e194975a7", x"8b3b4a650d9c0605", x"51d5a4a335c9765d", x"2bc2020f5bc20f33", x"6f386afd567f8b42", x"d6aab199735e5f60", x"0956e15bbb15436f");
            when 19568783 => data <= (x"fe62ece4cba4ff2e", x"76a2483488d68de6", x"4ae7a728c63c54b3", x"ea6652b76628b58b", x"bdac7e4305b3e31f", x"b98679cade460664", x"b8990847cf40b299", x"ec49a30a6b36bbef");
            when 31913700 => data <= (x"b5a961d55c6b2994", x"eabd2292448817c1", x"b6524e58454cb0ba", x"f7bd9dba6b185cad", x"599856ea90a34e7e", x"1cf69f88ec8ac609", x"87d33b489b9d1b26", x"f053301beac9ec42");
            when 25416806 => data <= (x"a62335b1d8ecb605", x"70366b31c4738f12", x"544e694093526b05", x"3af05de6745209f2", x"d1374a56ee49eac7", x"893b2ba01b4ca47b", x"2b7ebda5cf80c87d", x"8edc4eb355456f5b");
            when 2346170 => data <= (x"f141da2a4e2c6734", x"c5f630364f51165c", x"c7d9828664f40a02", x"3ce4dce9fcc961da", x"c47cbefdf2a8777e", x"e2b3aff319be7968", x"263c5ea460884637", x"4f50ab7e77302b66");
            when 19989569 => data <= (x"fd750b8fae18f5a8", x"3a81c6c6d468d31d", x"8e85b7ef584556df", x"394d67ae4e5e8c1c", x"bce961a9591ed303", x"d2c5219e34d71231", x"45dd1d399cd42acb", x"b4f54ea8b4959796");
            when 9239853 => data <= (x"d0e265e4519fe81d", x"bcf109b350b3a3eb", x"690708c552d4b434", x"85613d8673537157", x"37fb95d77138458c", x"5f34fdf7d5d9b28c", x"de6ef2288582e260", x"20ca66d829266a4d");
            when 7490193 => data <= (x"2d7ce4e03151b458", x"1a0c6addd91e7a06", x"45908af45f7205be", x"3de8e05e0f6fd8d7", x"a5c5ad66c78db5dc", x"98402072252ae9e5", x"505a6686a2f2e296", x"0da4300d738aea64");
            when 18833292 => data <= (x"74c94f423433e74d", x"622b1a43c7e0dd5e", x"9ff1d57ef7e600d6", x"a6c88e1567cba97f", x"6459daa3e4f5b6b5", x"eee76100dd514c11", x"2a2f0a3734d3bdd2", x"1426bec199e95b11");
            when 27712304 => data <= (x"a305aa962d954daa", x"75f3acf24586a713", x"01aa0500e4ee03e4", x"920357cb22b6c72b", x"9880acd01d249de0", x"63880759d6283bcc", x"1fdb1e0d61eabb3b", x"028fcaa9c9eb5e7c");
            when 32876326 => data <= (x"48d0caa7b24f0b42", x"3a12e9307feb1776", x"a971e571a7e3bc41", x"3416459ed8e8b379", x"f513a3bf713e9790", x"03e7db9c49802d63", x"07f78cdac3a4ff2a", x"894bde456892fe3b");
            when 13235404 => data <= (x"350dadd6828920bb", x"dd8882b565632651", x"144d8a21ad124170", x"086ddafd1079c0a1", x"231929a34c3ff2cf", x"6ad7ac57ee3b755e", x"23226cb237397c03", x"37c7909637e5b3fa");
            when 33362700 => data <= (x"efa6a0493a02c0fa", x"bd1a16ea43db773c", x"b4dd68b95fcf4086", x"f5d47a9d23db01d0", x"035853b574062a81", x"8991fab2fe685f2b", x"dd87ee0322b683f5", x"4f31ce2676f95bca");
            when 30997786 => data <= (x"d27bac217dba2ef9", x"da613ded0f75ff0d", x"7f6ad07c4c2f5ffd", x"c2b240132586bc46", x"883bae9a44db22b1", x"e74b785dbc2f14c2", x"fab08a769a3d32ec", x"e35a4583d9355ded");
            when 32393319 => data <= (x"04e89ea2e66626b2", x"a8f596607e9c92d2", x"46380708d5d7b7f3", x"7396c2cd27673724", x"4e85d030a706311b", x"792f04a95474ec86", x"7c79a7878cdc3cd1", x"2e882ca7a6797a0c");
            when 29714957 => data <= (x"76fecec1082fc22c", x"cca9fc9783f7450c", x"8d2fee6784ca5053", x"af22e2563d84b7f8", x"3068d84279cd69cf", x"7a2a86b6962b47df", x"b6b86e483d921932", x"742eb8d398eab475");
            when 33427283 => data <= (x"68ef7f93fb560a09", x"c2bfbb2c428fd56e", x"4c59ee2729642718", x"c02cc981f928e370", x"d2d7a074ecaec759", x"acf858327c28961a", x"3f87f36414faae9d", x"cb8d0d36908bb6dd");
            when 7239764 => data <= (x"c0147b6c7ae6de39", x"3ee22e130bbd13dc", x"74a07223f7ae1666", x"54d43be42df756da", x"9ef1b13c5f7ffb81", x"c7100c6ea67cc3dc", x"8b5672656559ee20", x"dfc79ffc3685adf3");
            when 31810750 => data <= (x"ca4e24d37bdcaaf1", x"e65ab6953ee2e58a", x"ced8d21963821cad", x"be77203c1609d59b", x"becad97a7ee1dd8e", x"c92248f56cb37df5", x"21ec84d0786140a8", x"367b991f9f030e37");
            when 15693301 => data <= (x"5b26fabc3389cd25", x"5b1fdf96c8b83128", x"221b78cf8cd28067", x"ae8f668036c4c2bc", x"c638178734ed08d1", x"74b9c697f658da78", x"c3d3e2386ccfe8dd", x"d29d1b3fa7db3392");
            when 29379344 => data <= (x"ac8578402fa59e87", x"ded4055d7d12713f", x"3e50fec55b412bef", x"e9998b8da17151d2", x"4b3058dc54b81563", x"ce79b6416416fc19", x"5073c0d9ebc9eb4e", x"a48c22202ed09522");
            when 18993591 => data <= (x"49243a9b45f42408", x"cea7588b2d1f4901", x"cc077b3a796f342c", x"460b4b946c876478", x"889fec22961e54a2", x"21947b370cf5104d", x"8284c340b121402a", x"e92848dfde7ff515");
            when 9764975 => data <= (x"8fdb18ae9d17a65d", x"507d24b63fe9cd74", x"3fd40875c1ce314a", x"104aebc37af58b94", x"5a8dceeab3294187", x"4a9e4834a144be96", x"50eba785127ec07a", x"6e8048c4baa0f285");
            when 6452559 => data <= (x"a68e1bbb2c7f435f", x"798fb3d590b10ab4", x"2c619a4a3eb4c48c", x"a461c7ab61cb0247", x"a95b823d3880bacb", x"8404d4cdbaaa1283", x"4f3aa628eff9cbe4", x"f53cf0418330d919");
            when 16453485 => data <= (x"2b9f07b39b97fd11", x"17c4893f1dd5f9fc", x"add74020f74c1e50", x"26b013e939a2c3a5", x"7043149368aab49c", x"258405ee7a5326d6", x"10d45a62d2b2af2f", x"9e6a2498c29be3fd");
            when 24739673 => data <= (x"b2bab86a135d6114", x"492e67c342d9f5c3", x"9eb78c4cd85726a2", x"fcde34afb1f8bc22", x"50f0683c5dd7989c", x"e41f284707e26429", x"825b5af6961904e6", x"c26a80bc5f1f4724");
            when 24140967 => data <= (x"2ab10c5e4679a5c3", x"6206a1519aa1301a", x"038c234e1484fdab", x"5d768b0e7e645725", x"e353aca08fe69e61", x"35909068d8b41a5d", x"beb8540643c6f032", x"7fd1dba5cdb9b254");
            when 12967095 => data <= (x"5de2cd5e3495b508", x"e28964e42a08907c", x"325ac650d67c9b26", x"0a54b84eb5e38326", x"e02527f3e4bca7f4", x"9694b13a78ae4283", x"77575d008b159d0f", x"8512cf4dcb713d2f");
            when 20646742 => data <= (x"aea84891c68f8f10", x"776d6b94bdadce6f", x"6e875aac47a9dfdc", x"1549a65e6839f41c", x"1f8c9e42ff9715b0", x"4642adadd7bce0f5", x"2cddb96615ad60df", x"263eccf9156ddd49");
            when 27036656 => data <= (x"6f73a84b8e167e53", x"78290cf947af1c38", x"be710c195945863a", x"f947c564c82ee401", x"8d9176615464eaf9", x"a93f0107f2cb0c99", x"3ab18eeff4761847", x"45dce53677d357b6");
            when 22463815 => data <= (x"6065a0a4f4c6ca3b", x"59dd23ee740cac29", x"cac1fbe3412ff691", x"66b507a1b96212db", x"865c629339604894", x"415b97536bf5c95d", x"e67df3dc55091963", x"8f1639d612a0af68");
            when 8919950 => data <= (x"3703f096003e1381", x"e894eed2d991fd03", x"0992182e48d435d4", x"7ba5d0c218b061d1", x"14754b73ca911447", x"f980728cb685d070", x"8ba83b6a26805437", x"37eff55fd745bd11");
            when 27308762 => data <= (x"460740807f202aff", x"788ee7a3bb3aa203", x"09b55ca66b58fda8", x"b9d2f3e85d690178", x"7cbf5dc6ca9fd820", x"784c6502dcd598b5", x"7d3b20d3d9e580fc", x"d63dd6c02b9db3a5");
            when 1892200 => data <= (x"b915ddd29024034b", x"ac818930e3f3a4a3", x"73f7af60eeee5185", x"76e376f0a1aa0848", x"ae2b63192fb03a4b", x"311107384fec2e4e", x"378801d3782cdefd", x"82048072815291be");
            when 28511543 => data <= (x"ce493092f16c2312", x"fbba08c454c4a0d6", x"e3dafe44273ca58c", x"429028293304d081", x"23c40dd2e5688807", x"947cceaaf43b13df", x"76f5f3b6bd58b482", x"8061f6a8fe621d35");
            when 29330528 => data <= (x"3afb961e7f46b4ca", x"e81eb339cb744af4", x"9375da01b87e580a", x"8402e28e22c5f791", x"f412fccc44cb399b", x"9a971566008c0418", x"64fc731e90d3110a", x"59b06e49123c9207");
            when 15051589 => data <= (x"a73272636c93ba78", x"afbefc684a641f0f", x"6b652b8e1a6fe000", x"d680b875918391d4", x"314dccc209f5b807", x"f46e6fadfb9e8cfa", x"5f2a603d6ecbb493", x"78839bdc10155683");
            when 14656403 => data <= (x"e53f9c3ed4f270c3", x"2241124b0e862617", x"33aade227f2d578a", x"8eb8da0de2cd1b61", x"8c238e6b07e379a5", x"03be0f80aaea76e0", x"c9a222ef9131eef8", x"be2a9019843855a2");
            when 1120325 => data <= (x"f163aa861a0f8dc6", x"780ca04e694ed114", x"2f3832128b88919c", x"1dda1699805f7414", x"9d0136aec24d0218", x"4d9671edb3778087", x"aa622d76567d84fc", x"e926d7130ae2aac2");
            when 565841 => data <= (x"3243b9e51a573e48", x"eda4718ef822e753", x"b3abe567afb94e9b", x"5fe7804a8c675422", x"c7a72a148b5c4505", x"c56af8d04d7bb479", x"5b269f6aa2873c47", x"ae2fa8bfdd2732e8");
            when 29584927 => data <= (x"e587f57da9c2fc83", x"a9ad38e52b8f3c7d", x"ebe9e82b47bd659d", x"24a24c1cbdcf56a8", x"8e414d9a04417009", x"074b32e8aeb5a872", x"c056bb94ba36ed58", x"fb000f024fdf7209");
            when 32530530 => data <= (x"40a9ff6cd470df18", x"884984e0c22c0c84", x"6024f8e40b9e9a46", x"2e213a02c24c56bf", x"567f8735c7ebd4c5", x"7a8f1cc64f735b62", x"492b8c9c1399f9cf", x"7b41ff4d00410005");
            when 23869910 => data <= (x"624a59e3ed7b52b6", x"1ae45d7b3a6f51aa", x"1200161d221bcf84", x"f49fe1bccb20479a", x"a169346d9d9d09f5", x"c9b707ccd0f9e6d6", x"bdbb769b8aba19f0", x"bdc51ba6852cbf7a");
            when 29827889 => data <= (x"ef86d73e9f78bc3e", x"ffe8dc50c8639c0b", x"65758d4876203b17", x"044059583607fe00", x"3e1594974face997", x"1370f60d9b9b534b", x"b60d9087f13d9ae1", x"f27adf1672e6df0f");
            when 433336 => data <= (x"00a1a8cda7191a7d", x"20e925dbd21cf0dd", x"fe06556665326391", x"4a873c0f910f9053", x"143a043ccc6a07a7", x"fea6552aad074fc5", x"05b57e2c325d2751", x"200959a31e7bcdee");
            when 32217229 => data <= (x"067b0f7462edb1aa", x"293c448576a0fa54", x"930b7b0e369b8911", x"415fcff435c615ac", x"fedc170d70037c39", x"a24d4e9fe7c65c30", x"e8eb152abad4d76c", x"4d6ed99505b0f3b7");
            when 21367407 => data <= (x"6ab03f3bd9161c7d", x"8c23c97cf06135b9", x"daf5901b1203d836", x"665a5c07188a5ddd", x"25159bd0f5ba2f19", x"4f654e41fa58a88f", x"1bedce47893afde9", x"6471a2882cd2fc99");
            when 432615 => data <= (x"d679268c4936c305", x"b90e5551c5408927", x"2ea8032040efabd9", x"69127abd462dd807", x"0a329b07a206b0de", x"ea253d1aae5a4f50", x"99ceccd69007b583", x"759cf16333b2fd8b");
            when 29728938 => data <= (x"8f0122f47aab1282", x"6736fde3b1bb3927", x"22843ef67d3c13c8", x"6e17872396ba4c13", x"6fbceae325ed9fee", x"1378c9fd084207db", x"a9c515c90834f81c", x"549e596d74fbe974");
            when 25442078 => data <= (x"33d23a5d3a9ce8aa", x"73c1cab9013c9299", x"8e4b5b0389879930", x"76732ef57ed117ef", x"1cc6704918cb646a", x"040e98149c2cfa1e", x"a46f9186ac89f887", x"81bc49081d36fc8f");
            when 2523653 => data <= (x"c9fbccb4b28a4e9c", x"5e6c83a9e78c1fbf", x"135f84af19f36877", x"94a1c28c0cf98f57", x"f5a06a444124731c", x"03dc49486e2f06af", x"05956b892e2de8a3", x"f3a25f740170d0fa");
            when 31150270 => data <= (x"d704c82dc0c37faa", x"6e258b3896ef4c95", x"c725abb348da5de9", x"a829c3d590587df5", x"0c551b6faac01282", x"df6571fdad629ff7", x"aa8c5d11a1f18486", x"246b0441919736fb");
            when 15232426 => data <= (x"969246d2e616e325", x"ddc7d7140f095a07", x"a5236b021811507f", x"9ed3335409e0f356", x"b60ee6bafaa33f73", x"e2ccb2549c86872e", x"28b034dfe39a1c1a", x"c3bb42dbf54a169b");
            when 13680309 => data <= (x"102e429ea9c39f80", x"315a264be4a13e87", x"f2ffe5e396f1fdd1", x"1173e224ee2bb6ae", x"06b2f3d528ac341a", x"ddadbee5b9de2fca", x"80b3e27f9885f8ec", x"8fc979f752d97a2d");
            when 10366711 => data <= (x"41e5e9f61e481020", x"c8bbb7fa074fa323", x"5d21e0cc840e152b", x"bcdb764660a5ea16", x"0d06fd2d238e1166", x"96edc087afb38945", x"7e3c697a39fe6076", x"385888328116dce8");
            when 24705603 => data <= (x"5946be93c402199c", x"b44597dafde5afc6", x"9b7d46acb93d38da", x"de5ef0bad24b5786", x"222394d547b04b5f", x"e32f4e845f881523", x"3377298dce090023", x"9063b0105c340970");
            when 12447941 => data <= (x"a8c6acf2952ec4ba", x"bafefa6f7358b26a", x"1cec812877cfb9d4", x"97431abc6cc77171", x"6a000a4d32dffda0", x"e79dd9ff8138d8ec", x"a948150cce353b05", x"55c1587145111d4e");
            when 29095052 => data <= (x"05b8d9c5a654bde0", x"e76c7439948da38e", x"4f36964a13005642", x"f64dc15c9cb0ad1e", x"bc0ee2840d3cabba", x"7853d422c5b88e1b", x"81bd41eef4a19e49", x"d662a9bba2d77f47");
            when 18826398 => data <= (x"d3a53e084fc23c83", x"04aa1a729021fdd5", x"4ccc25293087def6", x"774cb8df96a8e773", x"0343e4d32823b18e", x"26c92d3ae947053a", x"beeb556102c290c2", x"0ffc60e87fd026fc");
            when 27162085 => data <= (x"260c2eede98abe9d", x"b69ea764f8c0c2fa", x"9a82db7e33be661b", x"27233f02941eafe0", x"7c3b472abfa995dc", x"27e379470d836a7e", x"a3bde70bc6a057ca", x"4c5d6e774bffa4f5");
            when 28704864 => data <= (x"90c2cc2ac356b3e4", x"71c6ab48e2808dfd", x"c1699de9f7f2d451", x"aeb0a789a6d65113", x"80a099dd3e2f9574", x"27452fae1e03f2ff", x"177b95c624476c72", x"f7865a04fa47a4fc");
            when 12116065 => data <= (x"2c43b94bda0996ec", x"f04b5ba19c52a911", x"006115fdb82510a0", x"8c3aab60e4af9269", x"0666f86ae1cb2f71", x"3ad68feef473d254", x"bcfaf50c03d79995", x"44d1bc4fac908f7d");
            when 17788858 => data <= (x"5ec9ab6b8c459b01", x"6d21cd5d50b128cf", x"3c871f0cf79c55e2", x"11475e1cceab516e", x"514ff33c6776aea7", x"408d581da05c8f8c", x"821744e8bb46df05", x"a7bfd93368f38dff");
            when 22994287 => data <= (x"6516ac3857e3e978", x"fa4223d02620d2b7", x"2e5071371d4aeed3", x"ca0cdb48cf7bb46c", x"905a7e537d08bec7", x"0c0913d079f4d915", x"a3c7120ace3ab3c3", x"5e2bd0477727dcfd");
            when 4657035 => data <= (x"fcbf65845734767a", x"0cd6968135dc1a8e", x"71937abd942eeb0e", x"f9aa5394104e7c29", x"e3df2830426d0e3c", x"0b21e95ab5916ff0", x"81183caf464eb342", x"70d9c079b054698b");
            when 25528588 => data <= (x"8fa643dd4e627681", x"50887ed35756530a", x"a073780479746493", x"fc703040ef017e52", x"3cdbebaf0cc4524d", x"b95261801f78d4f4", x"527c661dcb9905fe", x"6efa8cbcb161938c");
            when 1627554 => data <= (x"446e1b408efbd585", x"60f59c10205731ac", x"1522e70720f1b9fd", x"8cf46cb669546649", x"4cd18f529527a7d8", x"20e64e6056b4f1d3", x"f6a6012414e0ab8f", x"97f89fdce77febcb");
            when 22738591 => data <= (x"30a12a641a744b21", x"f2ebcf9ca0c92e49", x"acf6cdba88af1413", x"425146c7c49bac09", x"a40b3c37d17be08b", x"34657977dc5eeb11", x"3974a840e8bae709", x"cbce806f4ef70b08");
            when 11910269 => data <= (x"fba369d36042b10f", x"0c521bc852bd3e0d", x"a4737e96f7f56857", x"40697f0feac04357", x"c2356e150fce2fa2", x"b4265598ba2b18d2", x"03b6827ebf049d64", x"f547f1d3c55828fc");
            when 31480480 => data <= (x"f4b6ba735807324a", x"d6ffe81cfdd5eee7", x"4413ed7133fc4285", x"896f22ecc893066b", x"1a9155eb59970827", x"2d522b07b876afc1", x"2e8dc1729e1db5fe", x"367662f8e4ff5397");
            when 19668739 => data <= (x"2eed340f4fa1aeb8", x"1a05744d460c1274", x"5fd19882caf789e5", x"dba5c11f43736d4f", x"349bf0714acc8b9e", x"491e8dbed9665c80", x"967f3df79db0ebe2", x"8848b86a1052c403");
            when 29708523 => data <= (x"6f73b3b07547ffa2", x"21419e993a5c27a6", x"93e0e3ea29272678", x"ec13bd0260e01179", x"3c44dbbb723607ac", x"5e2ba9c9ecbc84b6", x"8d705d3fad746fdc", x"b969a28c9a73bed3");
            when 17194137 => data <= (x"c920df6c66cd149c", x"3269bb11663ef9f7", x"c8f514aa8098c6c5", x"0ce351582634dd19", x"3c35e9435cf775ca", x"c8d34d3e90f8a657", x"f7ddf4c9cf14e184", x"c88fc9e682087cf5");
            when 15190823 => data <= (x"18159c6a6a5969bc", x"1f7301de58fb5859", x"8cb5052bf7a1beb9", x"c10d6abafe746ce1", x"54bd0f191993f199", x"022ca990b5baa3d7", x"6c47377ecf39494e", x"275e2ac0300c0413");
            when 11861841 => data <= (x"01d45c449dbec7b5", x"1d3dec44fc051ab5", x"7e9b4845e524a3b8", x"45619866538980ad", x"4762f122b835defa", x"36f10de8a2c079f1", x"78f537144c6c5a9c", x"bde11bd928c7c6f7");
            when 26841388 => data <= (x"43affbbc12a0b997", x"8e1dd896a76e260e", x"6511162cea120ca1", x"5f5eaf767f62b880", x"9e7690567e22f315", x"aa5bce67e4301ede", x"26223653a50b0348", x"3032c8e37e26c43c");
            when 7044405 => data <= (x"0506e0d57caeb780", x"aeb437fb06ac41f4", x"8025067b3d889a85", x"b76ad155ea2dce44", x"a3d7143666380079", x"6d7d43530f14fc2b", x"186f8e61c82b60c3", x"b0a6f99e6327e5b6");
            when 7878837 => data <= (x"4f1a73ac06910916", x"0520493e8e878e19", x"b637e91f60f433c8", x"681440dad602794b", x"e3264495163a9e63", x"f90f6572b55928ae", x"d80f22893b01442d", x"a961e3f02f9a1c28");
            when 23052568 => data <= (x"e6ec0a6654cf7ebf", x"caf977a9b6c24edd", x"9875747ab2d01ed0", x"ec7251462ff354bd", x"a5a8bf0c813fe96f", x"f36cbd6b2cd19317", x"5d1e253b90f18c54", x"4176caca2ee1e3a8");
            when 32040569 => data <= (x"cd8ffa3f3a36c9ca", x"0d73ac22c375a6a9", x"a420cb4c49444a77", x"0a1cc725c5dcf9a5", x"bfcfc6d2a9028d59", x"04272b12665012e0", x"398d42b3aa4a099d", x"76eeb3ce77fcfcac");
            when 28109610 => data <= (x"6180af2b92c727ae", x"20bf79dc20932b68", x"0bacc6162e983369", x"7c27ddef35983297", x"be161c2c5403c14e", x"19f91d5b6b9c588f", x"51e2723cf3547eb5", x"20124665e7c75909");
            when 12026964 => data <= (x"3d8c62304965e5b6", x"957d09d821150dfd", x"dcaf6e12a1be21c8", x"04e51da9ee7aa887", x"fea3d9374a18a48d", x"ab5d2096aa994646", x"8da1acd7aa90a101", x"82fefced5613bcd8");
            when 26816970 => data <= (x"2c388a5bd68f8c4a", x"4d7e4828bd899e94", x"0b2516a7db641606", x"d07c1db7fdd123dd", x"5cd93db31bebb627", x"3e0928fe6eee0be2", x"cb6cb24aa738a5b3", x"6b68de909dd1eb4e");
            when 20002580 => data <= (x"f055dbe35d7b4975", x"fc1a6b3c0bde1695", x"a1252289cd6edc3c", x"bc67f3eee9addc18", x"62c4c53387e86896", x"e7deb8021f1e8ba0", x"0b0aa20e6d08e698", x"abd12f1472a944af");
            when 24734402 => data <= (x"bbe65158a778b327", x"8e02cdc0ca20eff6", x"f11e7c6152ab7f99", x"92089b9d8d94239d", x"39846fc8b7aa622f", x"2ea381ea905cf3bf", x"fa550f5f7000ac23", x"8dee1b0399902bcd");
            when 21852629 => data <= (x"aa1ef99b335b4933", x"9aabd7b28a9a1fb0", x"f036cfaaee6eb3cc", x"4221faf62b5f0de7", x"9edfe2126bb477d5", x"52bd6ad6e0ebec3c", x"f0f61b2bf41a463a", x"f2cff5eb27eff01b");
            when 10345392 => data <= (x"b3d0e57f5de0eaa5", x"94e3d86be7c82056", x"8bc0a27d7d0a4fb3", x"022f2f37c40cb963", x"59236be51839e72a", x"4fea4d8881caebe6", x"0958421220fe2f77", x"15e071106218cdb1");
            when 23227940 => data <= (x"1b215d8c781e97c3", x"c19be166f5bb3961", x"ea6661d153345d52", x"9b770175ae11829a", x"827ce340727881d9", x"83a4d4f5af3423af", x"30e66353134ed11e", x"3b0cf01719905037");
            when 20432199 => data <= (x"e1b14bbf77e4ee83", x"7013c92bce383a50", x"4546f7d658c40e31", x"d1892e7407ef655d", x"dbe4c32452ccb28b", x"ff4f4cbcf7086625", x"68674e188d112129", x"724bb4d0dc0d8ded");
            when 30039548 => data <= (x"092df053eb8c75fa", x"0bd0484386c7d378", x"70fc28995b4e4e1b", x"6c10f4202b3db3d1", x"811134b1fb4cfe00", x"26a3c5ee6f71269e", x"fdde3a171d2d40ee", x"999ef39fada709ce");
            when 22483436 => data <= (x"23585cca18a6b091", x"d7ee3cb6aeb69c26", x"723690059ed77d0a", x"b35a785f2f699977", x"6d26e6a0dda074e5", x"af59a408d5cd5f6d", x"0beb86e2bdfc96f7", x"57334748dbaa2988");
            when 11477175 => data <= (x"971a13e4fee7fb24", x"abaabd56ab632892", x"7636f232f900e397", x"5e93eddac6a77f32", x"fb813692ac1781d0", x"b4de9839ae296fa1", x"8ca3408a0b9b0c79", x"3c32a9c05c383005");
            when 12607220 => data <= (x"5b8e33d478d8db05", x"0cd8acff1ed8094c", x"90a3523c635988fa", x"70a784c9255c0f9b", x"0757cf9454d81efe", x"689f83536008fd59", x"715f2e628d463b46", x"134282e6c9b6fe37");
            when 24255255 => data <= (x"534648ea421e5281", x"c28c9e51b0c138e8", x"85d0874dcc67179d", x"ae32a5712ed01c7e", x"be0c8916754de778", x"c20faa4f3f359c55", x"ef2fd73d170a2020", x"9f43cf043611428e");
            when 8518583 => data <= (x"03e1d967d09260f8", x"926a4335611c0cca", x"df4e79d2eb2b62cc", x"602a6ae14d72f8f6", x"13c4cf8117abfaa7", x"11036237289a69aa", x"349436168d96260d", x"885134453b652a5e");
            when 31701159 => data <= (x"fef9f8efe7eb49b8", x"34a0e073da06cb99", x"566faaf94e961f86", x"1edc6468e9772fef", x"b5764e48a0b50857", x"0b6230a9e5de1213", x"b4cb1c6d06917f83", x"86625f52fff81d83");
            when 29228307 => data <= (x"3ade6344a20236a1", x"4f270690739113d9", x"5db38d614296a162", x"79c0749998f6dfd8", x"237205d2822d91a5", x"d5fcf53b25685a3a", x"bf0e938992782fd3", x"8ef27a7476c92632");
            when 18507820 => data <= (x"f892c1603beabafc", x"08eb01db2c6d0a1f", x"2671443e671acd7a", x"8187d31bc127a6c3", x"d2d7e5966ee393ef", x"52b3486a201aaa84", x"5c50d80a4d996d12", x"489c48a62b21e3d6");
            when 17402748 => data <= (x"1fee44c2f03b07a1", x"0590918464f624ed", x"aa9f980a52ef6976", x"69e24e5c665f66ee", x"b6c5559c7212249e", x"fab23a96d82f1d4d", x"a9baa465a7821cc6", x"7961a8569ecc82c8");
            when 6112414 => data <= (x"38463b0cc6538cb0", x"fc03d626bb39eecb", x"c2bc244ff4aefb3f", x"b276f998d777621f", x"b0da3d6aa43cafb0", x"3c415f8824114ef8", x"ecfad457e661b56d", x"16c5fc4ef1857629");
            when 12160826 => data <= (x"32d0246b9d83ebe8", x"2b91fd4998289da8", x"a037d41cc905e1bc", x"8ace2269824def5b", x"d232151f9c7382db", x"98e2fd6297e66940", x"403d704ceb86f3b9", x"5641c3f6ac62a4b7");
            when 9468419 => data <= (x"1e9e33e381794137", x"e3e0ef6b827d04a5", x"72ba5a695a7d545e", x"d963e07880eb554d", x"b1fe7cbd5107226f", x"55d5696df63d1186", x"ae37edeb62cf7afe", x"71bf9dc8e6962279");
            when 9479989 => data <= (x"73618f483af77cce", x"720b297a1a55530d", x"4cfdc2148cf02d5b", x"34346d8e4b80d91e", x"7d15f78f2adf7186", x"52fe235cf265f109", x"9053e1e4de2b663e", x"51a383a68b6dc4ba");
            when 30222790 => data <= (x"ff24c078455d799a", x"49e5f13d849d61f1", x"69e0d900ae97dd98", x"6c4e3723507aa6bf", x"86aeaeef7b72848a", x"eb5a7bdd0197bba5", x"dd3a35efecab506d", x"53274b15fcc6afa8");
            when 27383654 => data <= (x"9b79c9419abdc179", x"54164d6bc3cfb091", x"b47e0cef821c8ecb", x"64f927695b6d8f26", x"c2c241c068678d80", x"a7de812dd0dd32ff", x"45704a099cee3756", x"cd6328981d239db4");
            when 3938523 => data <= (x"59dc9f3bb08aeb7e", x"a4f1494d9ccb1942", x"dcfd3f021fe00598", x"02e4f7f9fe0126e8", x"7976c67023d0056a", x"adde25bb8a896e8b", x"7084d0440bb7452e", x"519ca683d1f7e492");
            when 31237071 => data <= (x"a63264d12821b99f", x"97d3b783be297e74", x"3f2273ea27a8a279", x"e8f57cb9a03f28cf", x"cc4b4f824e25d2c4", x"5325c702398df2f6", x"f1189d6a66a74bce", x"795a6fe2db365af5");
            when 1240880 => data <= (x"b95fcf674ba669d5", x"5ec4283b0d5ad036", x"baf8fd540d0c5d38", x"be21c9a6009e6fd9", x"efc7b02efcc02e86", x"843d3904df9ba3fe", x"2a994fcdcf0cfd47", x"ce5bc6f27a3a4163");
            when 28939387 => data <= (x"77d5299cb7e6b996", x"40592f0b3d4a35ef", x"c5752a13649bfc6f", x"016d18d7347a5eb6", x"ceaf34fbf363ff74", x"cbd60923eb53c943", x"c6b04175ff3be24e", x"e0ef2cc9bf6a6aff");
            when 33357682 => data <= (x"57a43784b2b4e210", x"83eb53538e7bbc8d", x"f0532249ebcde8e3", x"5a62a92fd59baffe", x"1ace736093c91d38", x"fbbaed858a615623", x"94030899aa530764", x"cb77f43f254b41aa");
            when 26172860 => data <= (x"c43b9ce2d9e6b9b9", x"0750fc1bbd3612ac", x"99cc2366895add32", x"88964f6fbd7622bf", x"1a27f3a7910f2928", x"8f72c04b5b7f36ba", x"475547df72a5c7a2", x"f558b489311c21ec");
            when 8135826 => data <= (x"4574ca986bc77b57", x"3be4ebd1c487689a", x"d8c368a40bcb9635", x"71d7f5f448562b48", x"88ac987e487dd1fb", x"e33a05d2470a3a19", x"53bc54ee349dddc9", x"07e46b5426fab62d");
            when 5864718 => data <= (x"1fd4fb265ea046fa", x"668b956ad9bdbacf", x"4c23af129392f872", x"28d6c73261653e2f", x"cab5e4682cafea4d", x"3d16e2f4d415e65a", x"9a8747507af09085", x"6e2f87da8f57e9e0");
            when 17813518 => data <= (x"4d2cef913c3ed48d", x"f9c51ff958451614", x"ac7f576f7408039b", x"01607862fb2ef0de", x"111de3f5af4eb0ce", x"bda592769930c571", x"cd0b06e869e9b6ae", x"9618ee43d8564ae9");
            when 15284346 => data <= (x"068cbc57a0808dc2", x"ada69ac3ea0e6d37", x"c7e05972b7056427", x"15579cf03a072dbb", x"61ea096efcabedfb", x"a6021ee0c958ff3c", x"d10e991e73304a9b", x"984eff16a3cee865");
            when 6350785 => data <= (x"5d94c69bb8e4f68f", x"6f91acd03ec884a3", x"c6c7164dd3c5a8db", x"a9a9ce76b53fc6c1", x"f8a11d11fbde5ae1", x"1651f836baa37ea3", x"416db2528b61ab4f", x"9899ee2830beaebe");
            when 15472430 => data <= (x"bd6559f1bdd0a47c", x"4ef429fbc3f33dd0", x"fd6b32786db7a521", x"a05c0c6dd9a43a66", x"198f207e047f87f5", x"2af61eaa911365cc", x"3dd233ea86da5afa", x"7286efc632f3f7e9");
            when 22319456 => data <= (x"b428ebc1c9c5d1ae", x"1b0b9f429ad50c28", x"f3945fe21d635f66", x"14f9921f8db85ca6", x"df3948a8b6e6a7b6", x"80d4a5c898a11ad5", x"1dd771e8f6f16b0b", x"b32e00548db1bf1c");
            when 30945950 => data <= (x"ab40dad4935bf703", x"6d3347e61315b20b", x"5131f2e776500968", x"f0f89f0013a16bdb", x"71b8e4c1dcf86c06", x"7f0ad85e566baf4a", x"cee3b59f0701f6dd", x"397518bb3a64c1ea");
            when 190899 => data <= (x"34bd3c539642306e", x"6f293423eefb7740", x"37771b041bb12e6d", x"50b4949e62266761", x"548cef3f68e9ff8f", x"9da20a1c1a2f2b43", x"3063aa73e06f4956", x"04b0e676eb339948");
            when 16627847 => data <= (x"76148872ba3735e1", x"1fa11d6711f74d95", x"05ffd549fd69b5af", x"9c05fc8d939ec69f", x"980ebed776f3f04e", x"34fc2cc9d2db87eb", x"3e4d76e54858a8c3", x"34a97a0341774614");
            when 6333522 => data <= (x"069352308cca09e6", x"17d4e0c39ef95436", x"36ae1a57a9aaaddc", x"0a5c10ab57ad814e", x"2d8e75f009fba4e8", x"7b7ce4c7fc689c56", x"ca8a36b99e0e0dbb", x"3d95aa8d7882a4d8");
            when 15754998 => data <= (x"fbc6fb03b2551509", x"22073ab3fe4e4041", x"d72c8e57a10fccf3", x"70ea31d4699ac7f3", x"c7e6876e3de3d165", x"87af0cdf1b8e5b1d", x"2d54449f1b17791e", x"8e9acb46731ff1b7");
            when 29319029 => data <= (x"b7aad36117310951", x"61bc0ca0a50c4e0d", x"839c78c486c2cd4d", x"2cb3a559c3312527", x"f6e71f004af198ab", x"0c1bf02d26a19c17", x"5efd023af4466459", x"3f13b254504f8e9e");
            when 21487172 => data <= (x"e02577bfbd41f865", x"cc461a9a7f579fb4", x"cd3a7a91b07596cc", x"9d9f38820a57b4b5", x"4596652014dc69cd", x"ed739e4eb886fc0b", x"823090f1c865b02f", x"c6f34b9c7e101734");
            when 21913729 => data <= (x"8e0aa76c8e9517e2", x"a7dac2d5e01d20a7", x"a11b4a09798334e9", x"cecb1ff2cb377054", x"fb071afbccbd6927", x"4f59d7fb73963c95", x"264359972438a6e2", x"d7b57cff4f75cf81");
            when 21641697 => data <= (x"32598474ae99ab34", x"937fb3afd2a59145", x"3b5a8f8fd054aeaa", x"c0ce7e0fa05236b9", x"1659efa357aebfc6", x"c3a44aba2db40ebb", x"95f9abdfc8b9e071", x"4dc0868f2a83bc09");
            when 32274364 => data <= (x"83d715ffe1c507fa", x"9aa9c2ee2454d977", x"c39e73e0e3565c19", x"69d39eeb5bd18422", x"4dd29990ad5a28e4", x"4a5b7ec0e0ac98ca", x"20961d4da02b156b", x"b62a2c910610d0c2");
            when 10900055 => data <= (x"2f92fda092648bb8", x"254453e7873fbd57", x"ee003a424f0cfea3", x"a4e582bd8c0be429", x"d87b4bc30ba87963", x"68a5618591d1705f", x"8e54e6ea14214373", x"a54452bcbfd05b41");
            when 18972474 => data <= (x"def339c1517a228b", x"0b34e1d55b73227d", x"51692edcdf2d85c0", x"493731dc17ca671f", x"70d2a47cfea54cba", x"8adcc13c1294a497", x"974dd9fd71d4e0b6", x"bd599bd9ad89cba0");
            when 12067750 => data <= (x"c4bc3c1839945671", x"002fbb9ead21bf25", x"0b7991f4d40dff7b", x"bf27abe50faf0a80", x"3d8a0830a2d682f7", x"77368f626ff7e886", x"7c04331673cf1237", x"52ba59886b886c73");
            when 1014322 => data <= (x"bbe1b66f4bb965a5", x"b652d610dcbb8685", x"2b9fa925aa3ab721", x"2ec078bfc11272ad", x"6ad92535991cc079", x"0f31f0b267346015", x"18b40055c85dfcfb", x"2a56552b591a80d9");
            when 18419727 => data <= (x"d69a0c1925c4ad62", x"7f5f101d3801faf2", x"8bba8ca5a4cdee27", x"1ae64a82bf72ea49", x"5fc4b21dcb1917ad", x"4f1f4405864f7193", x"0a550c66e23369ad", x"1c76005aeeef03cc");
            when 21463375 => data <= (x"d0588ec2b7b5ac28", x"c779ceeaf7890fae", x"926e709ea0aa6e06", x"f1f33bc7a1bff7e7", x"24b741b080eba1ca", x"e33c727783aff7d4", x"f34656f653f11c38", x"28ef5a2cd3edb5ab");
            when 8960908 => data <= (x"7192d533ff28ebe8", x"0c262fbdd941e40f", x"630a13d2debf086d", x"4da1b45a11e35b66", x"05994147a0222960", x"6d67d789d87bf123", x"38e0508a7d94ea5a", x"9eb8e3b3ba1dab81");
            when 12572420 => data <= (x"3e6c311ffc047e9d", x"06c9cb260c0ac0c6", x"923c3d92aa535413", x"eda753290fa25002", x"65bf35f19a880701", x"cb74ac773aeb372e", x"0f0b5ff6c96d22f6", x"7d79b75609f54027");
            when 1934181 => data <= (x"96382ba9fe5e3dd4", x"61a385355020dd5a", x"0948d344ca9b7c9a", x"3b9160b297f0f975", x"6de120d55fef44be", x"1b6f27dacfeda3e4", x"cdc11bf2d239d2ee", x"353a72e27d0d2482");
            when 6357166 => data <= (x"5d58d6cb5c09d660", x"545e053291820759", x"c1323f01db118a4d", x"37a27e3af5ef6392", x"3df09b73b6de630d", x"c5948156848fe1dc", x"666fced012682f00", x"2c7e872a035dd406");
            when 24139259 => data <= (x"42dc0c1d949e439b", x"e4ef8da90f7764f8", x"b0f829f2abb98310", x"351e0177e3c176b0", x"1ea08284b0a8ce57", x"f09075bdd13c3eec", x"9d36100ba62799e5", x"ef9374547bd74cf1");
            when 21497415 => data <= (x"48f562724e1d26b4", x"761d2a4e88bbfee3", x"0c82b6e7c1e65ba7", x"43f0e8f5225a222f", x"0c5fd45ac47590c3", x"407f1e19a562ca17", x"afb58d5f18bf9575", x"f4dffa4bcfc84fa4");
            when 9413388 => data <= (x"628c3d59d8627f91", x"8bb0f7b06293cfe8", x"dbc428b45262879f", x"e7010f0e4536691e", x"660a7186bc0cf342", x"07bb21f22b1d7f31", x"174d7231b3d6d4c3", x"3a9dc9f9e00ecc39");
            when 6745245 => data <= (x"537b6bd9e9c7c27a", x"c9f2c087605f1a07", x"3b627e2c0c2d95c2", x"ec82ddb53fad53b6", x"96fea90696842aa8", x"b742a8dfb5e6342a", x"f74891518fa0577c", x"62dab1609a988d44");
            when 1600163 => data <= (x"e2cb7f4566adeaad", x"dbf0c7c6e1909967", x"4895dd8ccd6da76e", x"e5c32ea6fa96cf26", x"7d7f4404c98e8913", x"62aac63b7eabd890", x"297dd665a067766a", x"382a634f3f0023f7");
            when 30571928 => data <= (x"0c95faedec2cf1ee", x"c5a1b9d041dc8e86", x"f8342b3be3579004", x"81b53cb2cbaec2cb", x"5ef517bf762d5491", x"1bdbc55ebec2b94c", x"044e41d46642a31f", x"e463e5880b57c20a");
            when 24331850 => data <= (x"4feac8dcc77402a4", x"2469a621ee56ad54", x"98cd79f763ca06fd", x"5a29ee28e44b53af", x"c95f9223061f727d", x"7f6f544b1e34affe", x"65967ffc05d27571", x"3ab7e3e456645d28");
            when 17885318 => data <= (x"21377ce8948f3799", x"f58f05c91cd9b61f", x"f71541bd8b1dd13d", x"a092dcd0c9363783", x"ba0b54af05047ba1", x"2d186eb980945d94", x"02bd1d12e6beee1f", x"126a653d93640c95");
            when 2919911 => data <= (x"69bbd9ae1571c8b5", x"038efabe5e1c1d93", x"516935794e5b289f", x"17e99d56cd4983f8", x"9b8355332b5060f3", x"dd556d0519718164", x"cd5d157ba6fa580a", x"6379445d8b328f2a");
            when 14154463 => data <= (x"e8bd62961cbd0843", x"512f69e2c7257a94", x"e0641d2af7cec0dd", x"df3ef908759dd90d", x"b128b7a7e321406d", x"ec78053f8f523972", x"8825bdea264bb971", x"303e8eee7aa44572");
            when 16540353 => data <= (x"a43ccc950849ba8b", x"2dd6c5a52f009e7e", x"1cc12719bc3a69dc", x"d4ab55c38f1f6f4f", x"044709f776c4cb39", x"e9f056a46a959f98", x"2b12d3d755dae6af", x"8bd7394deeb9bd2f");
            when 5984083 => data <= (x"082da7c08565791b", x"b360dbaf600e479d", x"e17b9ac3dc3adbc2", x"af5e1f0b9447ec25", x"aea22d78e9fb78df", x"4f05ef0e2a8a4609", x"b4e71c26a3fb4f8b", x"efe2ef5bad2e9252");
            when 18798350 => data <= (x"d6b9c4448d718ae1", x"59c901e8959f847b", x"27d5bb43d51dc60e", x"79e24315affb293b", x"bc458a00268c3526", x"ad36425a9c9f076d", x"60855e9a65597141", x"f45839aa14e4329e");
            when 25712069 => data <= (x"c2240ce91f421491", x"59cba615130b4808", x"193000a654e7475f", x"90f33d0b26eaec76", x"e7f5c4e06d8961ce", x"9a940d8ea54cbabc", x"61d01fd73a91e611", x"41ff2357e2029860");
            when 26593014 => data <= (x"aa2356e3d24734a1", x"5852b7a48293647b", x"78d5bb5e2de56597", x"15b3ec9f1d045c43", x"7ad7cd0c4c9bcded", x"778f492d40040ceb", x"9a02d4406107db06", x"7b48195cd2a4f2e1");
            when 28204175 => data <= (x"329aeb40d59fc95e", x"c8e44fce858b3619", x"8dfa15b36efc358e", x"b3e7dde4231eb6e0", x"5c9a93adfcff83cb", x"60a7b31907ff1cc9", x"dc2fa1b6f2ca00c0", x"c7528b25d858d7a9");
            when 2683214 => data <= (x"ddf5a49b2e554f04", x"e1ea2a5a50352881", x"98dd5381db5bdb14", x"e81093a8e44fdab6", x"0a4be4453b187031", x"95047048537a2164", x"d5abb5a52884aacc", x"d7bd2f2f50bf6826");
            when 17944085 => data <= (x"f57300359d2c2597", x"09370b933e9d710d", x"bdd5dba74b5e95cd", x"dc03fc872bc915a9", x"bb4a6a47a7ea3463", x"f34379142de33e82", x"dfc3eaf5368a6334", x"5a75a48cfb74bc9b");
            when 15595260 => data <= (x"7d64244b36bd4666", x"386d87666b8c8cb5", x"e962007eb6ffdca0", x"2aaa9d59a9c551aa", x"d413f8b21d45dd28", x"17996c454517ce9f", x"609c624845e1bc01", x"fd7859d0aa4d72ae");
            when 4577994 => data <= (x"d608d48c7c369f71", x"669b43d5e34db304", x"f56e45f99c9fb5c6", x"63f445259868e734", x"096e4b7c9ed012f5", x"0ed5801e14eba7a1", x"82888f545f909bef", x"67d7c3db735cf189");
            when 9667508 => data <= (x"4186611aaeb23cb6", x"559c3aa9085e5206", x"355b2ce525f43e7e", x"437ea12cb2812407", x"55f4eac6951255e0", x"00bc1d2d010894b0", x"9a05e6a7845179e2", x"0a4058c44074ff88");
            when 31821830 => data <= (x"e1d28522a2de11a3", x"fb951bda076aa3ce", x"d89b4ff3fc170d79", x"c08ca4b2ada003ca", x"9ea6409598df210a", x"0b467169c747072f", x"5ddf9afdc73841e1", x"e2f7df0cb0e6d762");
            when 17917192 => data <= (x"93932371e1c52632", x"0a68fd28ed211ef2", x"f4e428cbd7d4c299", x"cbf33d5ad5849a69", x"21b2bd0c7729220e", x"79629e831aaf2d47", x"4aa2f4b993772a27", x"956f54020236b492");
            when 6413923 => data <= (x"eced5e8479ab6154", x"9cc72f85974f1601", x"f699a244d469b013", x"1424cbebca5a078b", x"fff15f64fe269b3f", x"00aa003af93e1439", x"59dd3a94c9d151ec", x"022a4be603dd9f36");
            when 18523940 => data <= (x"b8b91640bc4374a3", x"737970a82b6e07d1", x"d5e7d7cd88074341", x"f3d02a519ab85e38", x"84569fcc7cfdb15f", x"59ab4dec50e0e9d1", x"8076d0b1758f83af", x"0fbec043dfc80ed5");
            when 23605380 => data <= (x"05323a8e94237fe5", x"dfc966f19f4d7d1c", x"7058588c60d5163c", x"4cd1ce3eb6a1d19f", x"7af30e6f8d842739", x"9193472d0d113240", x"45643e76e8bcd4ca", x"126a46f42d899b17");
            when 20603546 => data <= (x"cf88cbadccc993f4", x"e9cf778ba129cdd0", x"99ddb3fdba5321a3", x"7914c780d2e43b9c", x"a0487ad4d77c068f", x"fab8b8ec943f276a", x"2342b240fc32ac17", x"960a5fefa97093b5");
            when 27940383 => data <= (x"1afe051cbceb108e", x"2406f8053f3b9c09", x"61005d4e9d8d158d", x"bb008c71d83de09f", x"d97ada6fe7648f1e", x"d85a072e0474028a", x"8536fb0cf26f3efe", x"f894412a28c9b66c");
            when 5581474 => data <= (x"843ef5d64f7ff0d0", x"e9ca0928d3b214aa", x"ce1a1b1deb1e0c25", x"265bb3449ebf030d", x"8f3564507aab0d54", x"dd55af05a4a8863f", x"0af021d8f5d82b7f", x"8fc1c77709903d26");
            when 20537037 => data <= (x"ec69123214c8acdd", x"d42535792996cb5c", x"1373251eaf518a58", x"7708eed241309ab0", x"79e505f267e98746", x"3322bc96b1a298c0", x"f5909b31e09a0ead", x"1bccf72107f70689");
            when 1861573 => data <= (x"e056ca0b443540e2", x"378dcd72613febf9", x"ee54a1e90af0aba9", x"c9f2cf6d69a75649", x"a61e24887cd78657", x"655b4935f8f72942", x"f573ea1f3e19a331", x"a7bd344f191af4a5");
            when 4929161 => data <= (x"6b2875f6ff86036b", x"0e61fd5507d33e62", x"4ed6a77d6259882e", x"bfbc05c0f5d4a2c7", x"b58829d91d0616d8", x"3611485d60b9b2b7", x"2458900395058914", x"4d1756d519d7eb53");
            when 22389026 => data <= (x"d4efd6b2d9a02060", x"33d024ecd72ac50a", x"4316de96c81ce5a4", x"7134449d05efc075", x"a7fa26046fe64e45", x"8e9448ad8914392f", x"962a690ff0c297ee", x"453feec6b091fca0");
            when 26542808 => data <= (x"f1deadf319bbd0eb", x"a25ee5d5b8ba02d9", x"8d834f2c1875b617", x"e6e53799052ddef8", x"91f2477d592368e8", x"75686542ac868571", x"2ce953e17cf6a535", x"5609a5ee4cca868f");
            when 6404966 => data <= (x"518fbfc748e48b18", x"85f14264efad59cb", x"fc85e6635ea2b2cc", x"4aa884c7c3d99bf3", x"67d0d5e24afeab20", x"3f9a254a80e5298c", x"c2eed06d922ec4e5", x"68a5e0de9a77cc39");
            when 3466065 => data <= (x"43a562eba8321461", x"52b87cc782b5d4df", x"c8fba14bfd6e2872", x"899a66f673918e38", x"6e76306037e6e88c", x"451873ce93dc392b", x"4fe1e419584c5a0c", x"5a9d02500cd8fa2f");
            when 8177972 => data <= (x"9b9905560e33d4fd", x"43a8b446221a998b", x"51dc3ef60e1ce4df", x"80c95a78d6ba7bb3", x"c5b552867686e42a", x"1b095b70195bf17c", x"9eda3aef97fae4a4", x"55c5c07f3f844345");
            when 18270287 => data <= (x"a872486df35f2469", x"e577524b14773fe3", x"5afb152ac78729a9", x"3a66c1a9ef72759b", x"4ab8882257d988eb", x"756ca13ecd577363", x"fc6284477b6163cf", x"9163c40ace60ab53");
            when 30780640 => data <= (x"ea974a2db1c592fe", x"a04e5a5b48cc8523", x"b4c315418c92036a", x"190795c86d9e378e", x"935809d811b693ee", x"c0cd8638a9dd831a", x"5bdf2bd0115349cb", x"f7a5b1c5be680323");
            when 2614098 => data <= (x"2e91089f802b5b45", x"c4018536939013b0", x"7ad01f36d90bce65", x"10099224d7acb78f", x"e168451f92468ac5", x"a36896d5cabecdb8", x"f693068f48bd5180", x"8c920080b7325040");
            when 5635717 => data <= (x"20aa0e6c8766718f", x"52a3ab9fb75a16b8", x"0da843e3f0191d24", x"8366b5f791f680de", x"32bc1d087addd573", x"609cfb65de26d55c", x"e097c20dc8176837", x"2a22317711453e01");
            when 15928680 => data <= (x"426fa5fe1fa34d86", x"d24f8fa074144474", x"0ca0496e7726b0dc", x"a2f6117ab3a1f036", x"0278293e1390c8c3", x"c0aabd57e885fd31", x"67810f5dc661f40f", x"684181719b78f276");
            when 28142170 => data <= (x"7d9b1fdab339c67a", x"c7a24ca6f89a2f80", x"5edf0d8f0f9b6be9", x"19cb80621e2e29dc", x"da5c2cf8d4575235", x"ffe3e29f38d08de2", x"2da63c77029cb5cf", x"e8746697ad046825");
            when 12714491 => data <= (x"dab5398072761d36", x"5f9de623fcb8bcbb", x"ae89281e82da94de", x"8dc9dbeefc79e1ce", x"2c130e4293195e8b", x"b4d30a1e6fa15d86", x"ce7a7833332692a4", x"08a0181e7c994ece");
            when 7800987 => data <= (x"b1c9ce46c06d834e", x"01fefa401cc74143", x"6ff7d9bb997c7177", x"e5126e92d04d67b1", x"b5143fdb628b16f1", x"ad9796a94cbce3c1", x"b522661099252798", x"8a70f97a0a47c86c");
            when 20873844 => data <= (x"0a31c7aa450d4722", x"7e658623e1f1184b", x"fca8d25406d8a3d1", x"b7d693dc8813a47e", x"40f1cd61c1a12f5c", x"c3048d9f54d3b5b8", x"c181b323a7dc19ca", x"a6eadd387b064eea");
            when 3111290 => data <= (x"a8d45c43de22532d", x"8f860a43fd06e70a", x"3ee70f4865390916", x"3ae29d3a3936d05d", x"9677b7e705934810", x"34cab6cd64b623e7", x"70129952e9bb9d7c", x"8868fc88779632b7");
            when 3441201 => data <= (x"bbfd012b79f9d71f", x"e79c26590b0a7e9a", x"561c2df28ad647e2", x"d367e71bc889886a", x"04b18c9a50e3988d", x"f3e36163ef49717e", x"631b886d5d2a599f", x"3becfd53ad8448b0");
            when 741144 => data <= (x"5407dbaf225bf8a8", x"c84c038266eb386b", x"0c90eb4ba3782483", x"e40e664beac56f03", x"c1e95f5291969040", x"a5a6305a5a777f75", x"249d4e03fa43ad35", x"cf24ddcac041a595");
            when 27422628 => data <= (x"61c03ac3862cdc6b", x"96e4a4813ee5f0bc", x"f0cb3bc80842e0ec", x"7128436df1240198", x"4981856e788295cf", x"43edb1caebdc5906", x"f080e08a37f71f90", x"45f8fd42a225a4f8");
            when 29707443 => data <= (x"f0bef0b33971afd4", x"41b2ac31c3c4387f", x"f9f5421402de56a7", x"4e951c49392fbb41", x"9c80793c6c708fd0", x"87128537f6ea45fd", x"f1876517517473a0", x"9f9ad7e9bc5c253f");
            when 7191016 => data <= (x"08d5a8856d35d13f", x"e292398c241eeaa9", x"a7636a961d60c776", x"b26fa008aaf749d3", x"3c0eec39fad31c4f", x"32273185d25c8dc2", x"53ef92254aece13e", x"a78ea9fc77235d90");
            when 17564663 => data <= (x"5fb41b46fb01fb49", x"43a2bc926cc82faa", x"d4e48e8d9d2b95e8", x"1ed9cbcc34a2e84c", x"9f5ededdc80cc262", x"77498570cac50105", x"2a11894c0572f0bb", x"34bbdd7c843cd8e6");
            when 30209187 => data <= (x"52dbf1c89bd66e6b", x"df9361acbc28a744", x"55b3b913b2a34b75", x"c0cd7a2995df14af", x"f858efd3493dfd05", x"ebf8ecf77469c03e", x"4ce8c32d230d733e", x"d7de0a54418571dd");
            when 10997132 => data <= (x"2a7c95f8052a8eb6", x"23addf2a29d15f03", x"59121e0d47f83d91", x"a62deec06f3d5d1e", x"22a44e8000271381", x"a88feda6372c62f7", x"8fa3a41800d4b0d2", x"b330e204c3613d25");
            when 2140135 => data <= (x"9eccc78742301dbf", x"6adc8ed3ab70fbed", x"016616fd75672550", x"cd240acea4bfde87", x"647af87b458b09c9", x"2bbfa2593571c902", x"cb0c2916623f0fb0", x"891358d96774b637");
            when 26120854 => data <= (x"7dd72e84af0ad677", x"cabc73b4ea08c31f", x"e9de25522028d2fc", x"efd374dd88d3e657", x"eed27bbf8fc674b2", x"a180d4c2c9f00682", x"fe2f38f9074a60cf", x"566a6f60d3a2e403");
            when 22024864 => data <= (x"74ff01394a3bdc61", x"c3d69a0c94ee2e74", x"5e485687d796b227", x"67860aa4a71502bd", x"836a8a9a8d6abfb8", x"ec4d12998404f6b0", x"75e5069bb83b3dd3", x"f719e9a1dfc9e41b");
            when 28639265 => data <= (x"4690555ef7b075ca", x"53e36d9ee21b33cc", x"d9386562f8b94895", x"4fe2cce0e8170118", x"25dfc0dc96929686", x"fc5741adcffb788e", x"68b9835e1de8250d", x"7e6025bab4280f57");
            when 13185521 => data <= (x"45738c129eaf5a92", x"698832c451bd07d8", x"69e9fe86bd0b668e", x"0286988f693ed766", x"183c366a679d8ca0", x"cae31b9addc1345f", x"975e4e22d24814f6", x"169d21b9749aed7b");
            when 17377595 => data <= (x"ec9936a8b68bbdd8", x"ca3e74cafeff41ef", x"5fb0a58c36cbd6bf", x"d7138507c3ec5a97", x"92861c2fb72f012e", x"045825b48c4bb50d", x"a060327be87963c7", x"f64884f141684acf");
            when 11567775 => data <= (x"30c36c67bf33fb12", x"973aa6dd03647b00", x"9b7a48aaad2e116b", x"e0153c9f614bc576", x"81921ada5aae296d", x"758aa67ea1233318", x"3083d8e7de49a280", x"4f780818ec8d70a7");
            when 19804597 => data <= (x"426612209434c40a", x"6273a6172ce684a0", x"48e6acd133c16794", x"5c85968d97dc0ef5", x"01e0a28e93039c59", x"18b3e3c1cb58a523", x"b008de0d203278d0", x"2497d258a61a1ac6");
            when 14694945 => data <= (x"9d431dfb028d88fc", x"520e48d5a9f5e736", x"9c601f80655b6ea7", x"3ef2f23180451a2e", x"9b40b13e6e9a4f16", x"478a89a9e3ea8025", x"90934895057eb766", x"27661d22f2742715");
            when 14342403 => data <= (x"ad4cd9d88d108ca3", x"6c855b36eb795eef", x"2624ee6ec3d043b5", x"a1522034816db4b0", x"a36dc68d0f59023c", x"f1a84bd8f118cf1f", x"363fc47d8993e16b", x"f8632957e55248d8");
            when 14068534 => data <= (x"1cc68b56b35c61c0", x"5cdbfd1c5be27dae", x"0a6a16403fbaf0fc", x"2c3cd087a42ce0c7", x"3337ab04a3770e50", x"201db67ba69d0622", x"a7e5a994025abb44", x"314b7ded8723e6b1");
            when 19168668 => data <= (x"493cf253468f13b5", x"90220e8de49a4cb6", x"c548ff95c02d00fc", x"6470362f50e2ee4d", x"56a9ab78e5c31cf8", x"d548f3cdee1e4ed0", x"4db7e973bc5227df", x"1c54e58d048329a4");
            when 33187722 => data <= (x"d5b7a5a1a9dba9ff", x"a9ccf8456c48cdf4", x"8253ea02920815dd", x"044321b42e9556f0", x"b4225e86112d9e97", x"82519c0d3a78a4ae", x"b30f88f1bd05822b", x"c46b740774dee9d0");
            when 5644562 => data <= (x"7bb3db321a9723cb", x"2d0e6308919d52ef", x"9394135c4bc44430", x"27b821d7a88c81e3", x"3166b1b6fa632cd1", x"e6309611c2cdd2f7", x"73b5f50d60813e5d", x"e1559d1d54e94ff2");
            when 31319121 => data <= (x"8af46eb240d90508", x"b1982dc11a1ce86c", x"0dcc6ea397e33e16", x"998fe946312583c4", x"9e98c0f0b7d4c162", x"572859907414f7fb", x"1f07fe166c3bb01d", x"efabb59b2a317e12");
            when 1081142 => data <= (x"cd0409b8763ec237", x"9de2b6f04f36740a", x"ddb26dca2c713e48", x"dc820d8d4033f5e6", x"53a197a0568c2b63", x"e8b211e33a63f88f", x"5495ea8b1b9c6bb2", x"5210cc57b6d183b3");
            when 17530337 => data <= (x"eb64c74055abe418", x"deddcc9e848bdd2a", x"09671329e527adf0", x"0382cbc0c18c23c8", x"0bbc9fda5c3349f0", x"d73d2119c42bd46d", x"43ad3e208f20f272", x"f1352a619bcc6aff");
            when 17344644 => data <= (x"7962785aebbcc9a2", x"8d4c5a0a3366c286", x"9ac2269f4c63d678", x"92c7febcbc37f5cf", x"d11341e6c4c54971", x"c6d83047b7f5a5ee", x"59d4f5574ac576e1", x"b919a89bda67c16e");
            when 13528843 => data <= (x"f6e362ca4dc8a562", x"2f1d469e32501c7c", x"b549adcb90d0edd3", x"f2da30034ba806d4", x"b2c9c8f20cddfc20", x"70f4c369228a92e5", x"dd50478d55bf0756", x"3bc9644e6c86d136");
            when 24415003 => data <= (x"c396786c9310642b", x"9613f79dfb21568e", x"62d6071ca2c8944c", x"70751371c79a901e", x"2f2889a6e52cdd09", x"89f7da18929b0b69", x"dc24b70cfd48fa73", x"d30d5afa93f28940");
            when 15930414 => data <= (x"06651a28ee338a4d", x"d6a8e98cbac30e21", x"721da1c7111ad30f", x"4d9d0606688e854e", x"96b245e87eee0c13", x"f2269b48e54d7ea9", x"a7780c981d52e42f", x"7a7b7321543f2fa4");
            when 8778235 => data <= (x"57036f94a66465cd", x"8382bb15371c7eea", x"279b0a4862bdb5e1", x"cecf8b9af82fc6d4", x"41c925720810ccec", x"480a3badec71e2c3", x"5003287f30f2e342", x"dc281eb3a53f0b8b");
            when 28447283 => data <= (x"156014eb03b893cd", x"602d795aeb7a925a", x"6e281e4dabb4b900", x"3b6970fe05366c60", x"e032f354197dd73e", x"2e77537dc9ac5432", x"1e5cad3b4684f286", x"8e76c51855aa1173");
            when 14395640 => data <= (x"30f6e4031e6f4828", x"ca18615057757848", x"c1cfddc04a58ab7a", x"16692b4fb6050586", x"6fd036eacd9c47fc", x"f3509665976d19fb", x"fe4dff2b66efccd1", x"084dccf65fc4ba66");
            when 16239354 => data <= (x"5247495623e299da", x"076a6b4e278db385", x"c8d856920dfe4283", x"3bacfa686e084bdc", x"251060b295eb00f9", x"31fb0aea6ce662ba", x"dc83d19166ed762b", x"f5a7d1673b322cd5");
            when 12343944 => data <= (x"0bebc5f3c1b99f13", x"b7fa363d2b9aeab9", x"e0b9e78614e0503c", x"18863da4d1d74ff8", x"6085ca0835609431", x"e4787da4ab67b660", x"623077ebe852f979", x"df83f9b5c29e3d96");
            when 16963866 => data <= (x"3a3412df03310a95", x"f3b9d879fc9ef866", x"6a438f2bb5d3cb40", x"395715149d275197", x"d89bbae800ec7cf0", x"207eb987975d987c", x"78e6a2f7e962552a", x"7bfb089191926dbb");
            when 15400984 => data <= (x"a876c2cf8ea21b3a", x"8a1967bbe716786b", x"0ba64724d2ce5ca4", x"0b54568a6b06fd75", x"f2dd0f9c043237ed", x"aeaf38fe720cea69", x"bca3e741cb6ac0ca", x"c901d1e4fa476cca");
            when 12905013 => data <= (x"12c2ee363dd2993b", x"fc3fa01ba06dd2c7", x"908b648c7935b07b", x"3ee88449fe897e0f", x"93891d11c072bde9", x"dc2ab7cf8d888a8e", x"f19daa14dd346bbf", x"f3c04d384a170697");
            when 24450625 => data <= (x"98fbb1cbe4edbf39", x"18bc6470471eae0f", x"7e5ce1a328d4357c", x"16fc1ab66fa3052e", x"5cfe9498d9bc0435", x"4c53486b985f85d1", x"db47464ded2c2e9c", x"2caa0b332c9aab20");
            when 5941248 => data <= (x"f221bcb68e5c2a36", x"a9f0a8100e07795e", x"4fe72075ecee1eb7", x"39d7b8c1ba4b0469", x"216baf5653655c0d", x"6f5ed1d42690ffb0", x"3ffebc0a47b15c84", x"3600aad9c89189c2");
            when 1621390 => data <= (x"7ac4defc9e718134", x"0067f71a728233b0", x"74ad9fea610965bb", x"7a0dadbc18365495", x"392cb60a2a966415", x"513c401c0800458a", x"76e3b84f97a3a0a6", x"d3a67b6927cf2e08");
            when 30818254 => data <= (x"a50d7bc877adcf3f", x"686c8b85e456585e", x"4c0ced95932fb605", x"1a9cd567fc1efbbc", x"4cfd3b50c88c2363", x"7bc0ff70eca19bee", x"134735ccae44381a", x"1819d3d11e42cf5b");
            when 27839407 => data <= (x"2190b2b45740172b", x"546de00115990f78", x"b14f80f929aee480", x"a859801679cd3a06", x"3fcd2ca04d11edd2", x"0d43a92cbb368042", x"b882bd05d416608b", x"bf93a7008fe6f057");
            when 17261707 => data <= (x"90b88d93fafebc6c", x"5c8f335b9ac1149c", x"3f1865002ab71fdc", x"024aabec7a32bce7", x"6ef51e1c6b8b4200", x"633013c7d7c44845", x"d3a9a303d8cb7f21", x"cb9ee71bc3907f58");
            when 2754485 => data <= (x"1f424f9623883484", x"1c8f9ebab7d660ba", x"a66cfd63b8435557", x"b8536d3657c3feab", x"466d7e76e78e7d6e", x"eaa1fb90d5aa4131", x"d8cd0b3abb209898", x"a3a699f938a6f76f");
            when 16351100 => data <= (x"ee9dad43c7c0b27a", x"938a444e123df873", x"3848c4518d214cbc", x"d7d8447a4dd5bec5", x"09bf7222c26bb9c4", x"d6893fc751320c23", x"ded32ed7d11e96f9", x"36003f825915d86b");
            when 16371121 => data <= (x"55adc628e9f32cd3", x"7d0934333e410918", x"bab09a2992ae3421", x"4cebd27259394524", x"b8908558e6475a62", x"d66599d4e3aa1bf5", x"566d0fa778240a59", x"10f187ce8e2cb820");
            when 16416333 => data <= (x"4ca0c144f4fe9a84", x"fc51efe8fbb58859", x"332c82e0cacb5f04", x"d6b2962be05994ef", x"83d2b7815c49dea8", x"6e51b20e3c79690a", x"d721b52d579fb876", x"0430d43289da75ae");
            when 1183386 => data <= (x"7811f2b5ff2864d9", x"94f6f707fe886f05", x"5042e13a127bb673", x"459d10a3cd69a071", x"bfe8a63bcae46c43", x"73cc5d2eb19e9f74", x"e8e7c0cdc56af2f2", x"3430b5f289aa793e");
            when 13765118 => data <= (x"efdff0d98e8b5600", x"0520779e2116d51f", x"4b70086e45bfb211", x"ac1ac5682f759725", x"95e6369f214acea8", x"7897345c01c57461", x"906d571276700906", x"734fd5f819236134");
            when 7417728 => data <= (x"51ccc84a3a9b128e", x"8950053271560189", x"c3c7f7ff8c9db2ef", x"c0a81551cf82940e", x"bec6850b2cb1155d", x"7c52cf6e996dc4ab", x"2a90449eb6c24324", x"7724e2f86242e308");
            when 12636136 => data <= (x"198a504a1600a38c", x"b0d9de28ad1b4343", x"ff0dc1dff5fdf6c5", x"d66609ad3b3e5f49", x"b0dc2b69abf04fb5", x"c637784760a13555", x"7c95983accdf0acb", x"2f564d1d8b08df7f");
            when 8268837 => data <= (x"525bcd73ac2e0fdb", x"8634277d7477b8b6", x"33b2692b99ed0a42", x"588c2e970f33abb4", x"6e0c579024321bd8", x"6aacc9d46af2f743", x"d50547fd42af2056", x"a171788f657f90ad");
            when 18657090 => data <= (x"f24ac54923eb5304", x"b40cc8f65cdf906a", x"2bba8208a19edde3", x"218390321092f587", x"790c86f9c9a67dd9", x"ae8762f58a7ee382", x"00eae895c204bcfa", x"edb9c8a1fc442b30");
            when 24033183 => data <= (x"35d4e583bcd4cf6a", x"eb7ca0aab2e1199d", x"1a85251a73ed1ea2", x"6113ed92625075c5", x"7f98d515161e1f9c", x"cfa0ba690dc64941", x"1f6f0ce98a573886", x"bec417f698e49f17");
            when 1529416 => data <= (x"6455292d0c6254d4", x"d044f3f43df30020", x"5b36ed3b4001ac78", x"1cbfaa015d11b711", x"c5525cef6169aae5", x"535d133b4e95c3fc", x"129846fa9faef7a5", x"fd5636435ed23c08");
            when 9487895 => data <= (x"05883858ce39b924", x"57d3a610b1c752ba", x"c9d3a9a3091123f4", x"edcacf486c535076", x"b9b689b1a041191a", x"82598ea8c67e2604", x"e2aa7689c880c348", x"6fcbc04fc4688e61");
            when 24125733 => data <= (x"38e15de417df408e", x"5bd49f5e24a1403f", x"16def45ffdbecbb5", x"c00f941a3afa86ce", x"8fb83cf086fdacd8", x"a440d8c3e2178923", x"51e349df11ca4185", x"5353e116809b6cfa");
            when 9729227 => data <= (x"5fde566478c67b0a", x"e75585c243df29b6", x"64fea98665e8b56e", x"2d4e1a6897e03b51", x"14dd3adbbf2eadf8", x"4c555cf04348aa9c", x"83fbffb90b324fd8", x"4caf622fdd0b7e05");
            when 17401648 => data <= (x"8a41fb7126ab76e0", x"606e86f790e25d56", x"aa9f499fad4471e7", x"2500eaf804a67b33", x"c41222c9cb24cd5f", x"a23a55a5a1afb2f9", x"27dc166fe47f3ab4", x"5f20b481731dba89");
            when 9019162 => data <= (x"bd3f260b7f24e4ef", x"29b9719dde979c8d", x"858b8dacdf9d1a09", x"26730d9606b19f5f", x"0a00febedc90f284", x"80acc2750ba87b63", x"ba472abc25b4b04e", x"af955a33d337eab3");
            when 6573122 => data <= (x"bd4c4d1e005aeaba", x"5e3ba21c0c8e4c5c", x"17a5692e4e1242cd", x"0f78ac3252b5aed7", x"86c5b3a3bb4782fb", x"00ab58e86c5be684", x"7d7cc1dede712971", x"a2541cb863b3deb3");
            when 10812289 => data <= (x"f55598e46f6a0f9a", x"dad330796f1e13ed", x"a9e2d246d472005f", x"aac8173e4c455878", x"5e84ee55c99d44c0", x"f06dd463c00989f8", x"97d841601572ebae", x"942fdf079fb8ccdb");
            when 14192101 => data <= (x"59573419a94965bb", x"e5239e644d6010b3", x"5993008032727a9f", x"de8e71d1b95a1f2c", x"8c9326c0ea7d0120", x"68312ccc1f7e87b4", x"13149b56bd1915bf", x"e95f5501e28b12e2");
            when 28759119 => data <= (x"96ab141e7cc46a19", x"c88d8883b4bf803d", x"8596fa9eda2a5cd0", x"0b353c15ba42f4ef", x"634a3cc66a315335", x"0c59743445dee2e1", x"71bfefc1d98360f0", x"0616c68e27931d10");
            when 2269572 => data <= (x"9932c8c38af528fc", x"947b1e7599732a87", x"3dcfe060eb218d42", x"1571ca812009b0d3", x"a3b50b3582a1425d", x"9afa08fcb76f811c", x"b5ce98cb3e8030ea", x"31c18bac300f273b");
            when 8866164 => data <= (x"44c0ef184faf7e05", x"cb91c5d74f592cd8", x"1b9088be8bd9c925", x"423fa653b262aa44", x"e9564daf078e50d4", x"2333c2a7cc1e8473", x"1f6350a01b672ed2", x"f72c7db5a876d24b");
            when 22455279 => data <= (x"d9b7fc359fef0ebb", x"2f534aed1aa23235", x"997844dc033be1ad", x"fd0ca2c00d1e3953", x"2b6d219bb35e7537", x"14219ff34bda3182", x"d65a3335f4660494", x"44e0839862db3684");
            when 3760767 => data <= (x"e881ee29886504da", x"c811c085eb2864a8", x"881291d4cc7bb86a", x"021879086dcf9d55", x"a577afcedd643765", x"747f285594c7bffc", x"656d969608891cb8", x"41f4731c8148955c");
            when 22023724 => data <= (x"819b29dbd47b3141", x"84ca7c24d9242d6b", x"88824390f6478754", x"e495b24982b837c0", x"8e1415812ab623cf", x"0f598098e64ec00f", x"5153b2dd78280cd9", x"5bb9d210bbcb5c07");
            when 11795046 => data <= (x"a8083d5f963a562d", x"a7072d119abd68c2", x"b89cf3cc40bbb3ba", x"7d968776cc8d2f71", x"705adbf5ebb29fd2", x"552d6a90d98ce474", x"89e05bb916dad2ea", x"380205e66c8ae608");
            when 7176324 => data <= (x"3dcc865fdfdef2ca", x"3c43b56d058c8498", x"7511d5c7e30e155b", x"22083693fc367090", x"b54654e697271513", x"8af9db5be58529f6", x"d584938bf3e9774e", x"0b74d5febafb8f33");
            when 26269237 => data <= (x"1df609c60e139331", x"70834f4a74f218ce", x"675f4c25f4e458d0", x"b26f7aa3628e9d07", x"58eafae49ebe061a", x"40e49bbeffe845c2", x"6cf01f51cf6fcd1d", x"04606b893dc9b79f");
            when 32788422 => data <= (x"7a53065162db87fd", x"8b24f2758ee906eb", x"86ad3782117a6cc3", x"2b25fe05f21b8239", x"4569dcca143b3804", x"d098ebe68a55db74", x"092bc188f0e8539b", x"d407134e8923aa0c");
            when 14469768 => data <= (x"6de3449816abe447", x"c63de826aebad7b0", x"305da4445f0e8562", x"683ba8c1b8f0fda7", x"2b985c2aa09b9b4c", x"8687590babcbf4c3", x"21677bb0730eaec0", x"4ab49ac044715811");
            when 2728519 => data <= (x"1e55f54afc4f226f", x"7c67bc2c12bc817e", x"4330baccd1828b32", x"6847150b73f1ec66", x"2ca132faf5d7c305", x"64fbd16296bafe15", x"159ec713312ef9b0", x"2a9e80f6aeaaaa4e");
            when 26148039 => data <= (x"63eab924909f60de", x"df5b5fbf4d54a3da", x"4685ee4bfde392aa", x"6ec0f55db9081d6e", x"b8d434c91ad91d0b", x"35f6480303002c76", x"93c2ba82d0fd4ead", x"665bc1392f8963fd");
            when 12586160 => data <= (x"24c75032f69224b0", x"654e8b3968b8f8b0", x"086c69335abef22e", x"9463b2cbd3a0bb25", x"581deabad76b75bf", x"848bec01c84af4db", x"80aef7180e92404d", x"e5e75675aa34920e");
            when 32431880 => data <= (x"2f37d1c53c1e2113", x"7c6af8c9f640da53", x"aed2921276d6140b", x"dd79bcbc1ce9afeb", x"bf3c627e4703a40b", x"79344cac86c4747f", x"c30f72a0a9b59d19", x"ddb744a91d1c883d");
            when 9648765 => data <= (x"e2737cce92df3feb", x"07363566968a283a", x"7529aec55680fde2", x"2b06093f8c498e25", x"1bd947d1ec76e7c5", x"e97ea890a4cc89a2", x"e465164118e01058", x"d78d674aad670199");
            when 7669662 => data <= (x"82732f89e365b545", x"2a0cfa965b8dd27f", x"6671cdde7e6f8d93", x"c997ea26b740c2a0", x"1c3f2d7ce46c239f", x"36a4fa6d8cf767df", x"4b05a11b704ee03f", x"c08821ecf479c7ab");
            when 30283821 => data <= (x"28637349a0b21a4c", x"a0087aa05a309ef7", x"899b88aad703060a", x"1cfbb0f84ad24621", x"4aafe6791522c3ef", x"dfa4e2efd94e6086", x"a73da09f990e3b54", x"bb5fd12a1779585f");
            when 18305887 => data <= (x"bb81865726bb5b86", x"043c9f3008b44e51", x"3e60f831acbea2dd", x"720513cf20a26697", x"473eaad7f8bc3de4", x"9a59811f1291a5cc", x"3e65c25af7346cfc", x"ace15b7e7adf507f");
            when 22469418 => data <= (x"f84376950d0dbe4a", x"ba3947002c3c6bd5", x"ad63c281d6ef08fe", x"6a03b3ad558e4ba0", x"cccdc7bb42350085", x"9c6af6644202e79f", x"228bf92dde46881b", x"014852682fcd70d7");
            when 22106438 => data <= (x"577e17cfb3582739", x"a3126487179c77b2", x"91007d56c3b650b6", x"0041e446b6b1bdeb", x"baf1328dcd9fc993", x"226d291cc9c61acc", x"9c858d1a854cd472", x"18e367a86307ecc4");
            when 11882268 => data <= (x"3f2491223b13a5e8", x"b766968a47dbed4d", x"314e6a45265e4ea7", x"5de26e0ae8970e13", x"2a91dc404905268a", x"c005150f1965bfab", x"45e67466036bd77a", x"4074c4c006bc3bde");
            when 22784217 => data <= (x"6be4e136ef99650d", x"346f444ca230f7d1", x"199615b4328e9986", x"0c63743eea489f40", x"10409f890f2aec5a", x"246f0f88ed31cf81", x"65eef82812e35f76", x"f22e5008197b0727");
            when 52161 => data <= (x"d8b28c6172c0c4e4", x"d127b7fe50f9b785", x"54b0a1de0db9c22b", x"711120e746384430", x"87041aa0e23a9725", x"32d8bdc0351cf0ae", x"21ba5d8b4fc348b4", x"c46cd0bd9f2f3402");
            when 4133691 => data <= (x"b4fc22eced723f8f", x"998f5ef584d20340", x"d8df5ba18479ad49", x"3805b4622c3ac90e", x"b426313bba92b727", x"278de2b61984f7ca", x"4eb1691354f751c2", x"d7ef21f65581ca0c");
            when 351438 => data <= (x"72044bb65f83a90f", x"0de674448a163c0f", x"68f10d87fbd567bb", x"ceda0600171204fa", x"3e7d73c0c6b1357d", x"78af7452a35be564", x"63069e5e17c3121d", x"46b61aebbea69e80");
            when 22498494 => data <= (x"94f55bbc6820d501", x"acb2545ccd0ad8ca", x"2c73c00c124dda9a", x"4c89cc9a8519c6b3", x"03156c7c3a987146", x"e2111a8bfc1f129f", x"de6fab7427562362", x"d995171a5606f68c");
            when 27205328 => data <= (x"06656970e71ff70e", x"34a19018cc204c06", x"29b29c9ab5005248", x"2c4ea164f427b9a7", x"7d04d43da7771a14", x"8c026a033558d8df", x"fd1cb9516acb21c6", x"4d677063d9400480");
            when 8805712 => data <= (x"74ab455b41b33518", x"e51c5ed1c3e91a06", x"bacdc09718551b53", x"13d8bf5f906baab5", x"ab3e9db1f0c90768", x"9eec604341cc80cb", x"8ea57df743bc53fc", x"e58bed2c3a0eb2c4");
            when 3203173 => data <= (x"351a3edd3afe5768", x"740bfa023171a6d7", x"062d2e9e57cf19e9", x"385b4f7b4ec39703", x"7d15b6a1fd803ac7", x"0f0148783b92ae93", x"d4f2643fae88d3f3", x"d94171e27c5773fe");
            when 32829206 => data <= (x"fbd4b72d9c0b9a14", x"f81308461d3c9886", x"b9694522626cbb7b", x"6ebe1381dcbb56d6", x"899e286c556de514", x"7515a835b3597bf8", x"6d7a159b088f78fa", x"a6b5d647a7ccb6f8");
            when 2093891 => data <= (x"04b69d64db166875", x"2ad9681d1d26d90a", x"782929b54b757927", x"8a7ded93ffdb470c", x"ea4428ea2457f984", x"9916c25b7babb173", x"a80aef1a90161786", x"bb199189d3fc82dd");
            when 12123594 => data <= (x"9c2c1e0a9b1bd6cc", x"bd1db6eb3dc76a34", x"89ba254a03382f73", x"86f85ba131feb6f7", x"7e5eed434b585293", x"f61f22831651332c", x"af73c7625ae41030", x"60607dbd0e10682e");
            when 23634164 => data <= (x"c14bc83e13a6b88d", x"f6158f8b11363073", x"281397eceb9e3d9b", x"ff3f3beb3cd13dee", x"378649d5061d6a4a", x"8a56f7640fc40b0e", x"2bba2c06875d7c9b", x"047713813ca3ee24");
            when 22951684 => data <= (x"072e92d2f97231d8", x"08c52cac39a8b5bc", x"ce89c531dcae1a02", x"5b8729b34c935459", x"637c81b98eb67e78", x"1ed26d4e20ff362f", x"c271ab257e54bf6e", x"178c05e4ee8a3dc9");
            when 13408610 => data <= (x"36b920731b7c497a", x"7a1155761bb50038", x"116a0be75fadfdc2", x"9dcc04ae1e0d4f51", x"524802c628826c09", x"b93a5953442ee390", x"a4bc2467dacb2f1c", x"e7f616535e432adb");
            when 7440644 => data <= (x"021e5ac4dfc861a6", x"288ffbf0207205cb", x"51c7efd3ced1c33c", x"f8e13ea380369def", x"6832a7e3e4396a7e", x"347f7bad248bcd78", x"b5b7dbcdac5e1023", x"4fc0924f3e458914");
            when 26716531 => data <= (x"52dc6830db5882eb", x"78f330895e32172d", x"025745a484942b1e", x"7f20d85da2cb3a37", x"2aeb10525f8fbda2", x"cdd90e1b5572eeda", x"c12155da794302b4", x"bd678c9da3f3e1b7");
            when 459997 => data <= (x"6ecd0f506ac0aa65", x"985c5d12bd0e0770", x"4925119901f613b2", x"427bfb46835f27fb", x"075dc8d710bba3b6", x"7c73e996007a3bb3", x"1000d910d4200a5f", x"031f4007e8e52e37");
            when 30679890 => data <= (x"848a40eb6d4768c8", x"f86820b7e61d6ccd", x"2807a67d7b318423", x"85eff1e59f67f3e9", x"4df9bc988ee7544c", x"9fcd8688fa2494bf", x"ae5dad8b1c5e8e79", x"b2c0b2512c22355f");
            when 17851564 => data <= (x"d9d2103163778fb3", x"6d4eb22cf38c3920", x"d83816944e5d6fa6", x"0aaaf1ff636b0ae9", x"4640be2926e90a17", x"720a9d9845f3c86e", x"043bbc60c85bd531", x"98d00483b02e83aa");
            when 5840855 => data <= (x"202e9164ead96c55", x"2d76fb6e2f4c5eb4", x"64f9d890395366fd", x"9596f54cd74d1351", x"2824978a0d92633c", x"2bcf7eea782de8bc", x"0791900002f378b9", x"2ba96dad057e3d42");
            when 1230377 => data <= (x"4330ded94b3100e5", x"237fa5cb984a38c4", x"500ff7f69e74fd27", x"89523d0afe8ad878", x"d5141944000e0094", x"547056e91f7b53ab", x"d73e4cec17015adf", x"c1a98fc8a7083a19");
            when 18915106 => data <= (x"2ca720454f6478ea", x"320ace01c2b3a215", x"3b592d5a47be8234", x"7112f5f176fcb9c2", x"284d5d29ebce551c", x"53913e2dc7aadfba", x"dbc118adbd45cb03", x"23b94ac7067a20fe");
            when 22472047 => data <= (x"e9a3f856bd2f5823", x"1ec0c3038f79eae8", x"c8188e274e792c60", x"af1b426038421cc9", x"3ea4926085304426", x"bf3332cf5d5f977c", x"cba19a1f711d3b2b", x"806d3eafac75d68d");
            when 31570698 => data <= (x"3dad83a672b2ef11", x"e780df6e29cad99d", x"c23016e6be95c7ab", x"8a642646b3f85e3d", x"dc9494d414106e2d", x"d0d7e78961354d70", x"91bdd30c59e1809f", x"64150f11b69a396b");
            when 1006506 => data <= (x"7121655a7c1cc5f5", x"8896a31014415dfd", x"8f60ac6b0c3499fd", x"057fab28f9c2b458", x"a9029a55b6a61034", x"a54bc92f32b4ec7d", x"80bffec0fef62a3c", x"fedea328f39dd6f1");
            when 7719222 => data <= (x"5d098dce0e1cd2f4", x"19b5eb59f5df9f2f", x"622724822b88099f", x"0202de12aa3dc7c5", x"9e9368678427ab1a", x"745ba4a4005a0491", x"06e5cb05fd7ce5c5", x"67acf96276189be9");
            when 15310354 => data <= (x"35a091482ae36dd1", x"af38f2efb2ef81a6", x"41af7907336e2c44", x"9f1a76d4083be0ea", x"9ac651eb40c584c1", x"6db61b7ecc4587f7", x"0c0cbe9f132d40ff", x"a1752ede6da6a306");
            when 1375696 => data <= (x"e822aac30c75f1d5", x"f8aa295270e4994a", x"e1c9e4efa24cdd61", x"f5713ccefc626273", x"be18c1a8e871f233", x"633a6c01e22508f2", x"a2e3f7939773c69b", x"31f4f1365a6326ca");
            when 16398093 => data <= (x"2d43e107f823a3cf", x"dd73a63699de24d4", x"f2a1ea96f6dc309b", x"31325fe259b7629c", x"7f0cf073be51c241", x"85aeae2c57cc4140", x"38e3cd89368b7af2", x"611c1d80724e5d79");
            when 7962330 => data <= (x"dd9db2665cbd4288", x"326a12dbe1cc98c0", x"778ef41b3f0c64ce", x"56cda48cf871f490", x"732b0aaf397f2a44", x"a48f4dd11b9426e0", x"e25112078a854ed0", x"56a3bd472580d977");
            when 1308277 => data <= (x"a6b24e77ba8bdadc", x"4507291a053189ba", x"eef1e1eba105c466", x"4dc11cf2fafa995d", x"6c927957b10edf51", x"7e2abeb1439690de", x"cbce25fe32d03c4f", x"28c9923a1a3d954d");
            when 16825763 => data <= (x"30ad28ccdfa41d69", x"6c4de0fc1faaba77", x"e405841ecc808504", x"34a0e6b0a65c3e84", x"c888fcd21843ed19", x"efc19585b37bed30", x"393776bb591d2b56", x"012664b4ca454315");
            when 2468745 => data <= (x"bdcc373848e6daa9", x"7c442cb29e7422a0", x"71c4893670a0a832", x"78e04bb7e34f8fd8", x"851439b16ac5e9fc", x"f67275db5f00c044", x"b20156b5f54246c6", x"5295bbd6db05ecad");
            when 1111316 => data <= (x"ae080ed9010c9533", x"877e22e29b63ffdd", x"b7dc4bf638f44e63", x"ab8d87f8a3901e05", x"738b58f571284d20", x"524bda05ef27dead", x"1259cccd00e8778d", x"f3eeb94270a571bc");
            when 92019 => data <= (x"e707c1c5b45d83bd", x"8ac0c6ea12ccad25", x"9eeda60e8da0ab4d", x"70e540c489661677", x"dce4d499a7a26a9a", x"5aa30ce2d8892636", x"d4a6fd5e4279da67", x"42671cafddc504f1");
            when 11399043 => data <= (x"6018ea6613a613e8", x"78d8c7e68affc8db", x"d6f97f9ad2f4299b", x"8ad320b12a6fde5c", x"666a2b66b2050f63", x"db6a7e81d25158e9", x"9ee41cbe0eea7040", x"9852bedcafc6df32");
            when 13059260 => data <= (x"27ea8fc3e5f8cf8e", x"d55753102731c0a2", x"b89e77aff0076321", x"93b40754078ceae1", x"1ed7ae4c4540be60", x"eb994f65327812ac", x"3de99bffa1a1a4fe", x"473bdd474833eff5");
            when 30648440 => data <= (x"1ad9bc52d2288007", x"31f8e368e6cf781f", x"421b04e81a8ce48a", x"612116a78413ae1e", x"7224764c38d970d7", x"5b3d0c7840c591de", x"7a6f0c4b1b0deda9", x"9ba4f5b10f12de3d");
            when 9435594 => data <= (x"e5feea484315b5c6", x"31ba1f9d57975765", x"0f4e7b17e8e2f52a", x"ce93ec033c4e5f1f", x"4b86365d6fe76be3", x"437fb26b52d3668f", x"db8c7e4b2471bab5", x"738e652a6dc1a60c");
            when 12426693 => data <= (x"eb90f16e2ab1b633", x"8fe3550354dd4c2c", x"4033d24726032bdc", x"e664c35048a260f1", x"984f29e529e9de6e", x"8ff2659aa285f5de", x"a9fa354d9fe241d8", x"44822eba7fa0dadd");
            when 16682510 => data <= (x"ae8ccca02979e289", x"b626890e2ce4730f", x"bc09ddc0325b7668", x"1a178c6da0031ff7", x"ba88779889fd03d5", x"b07c294fdd39630f", x"a6b4d797bcab6479", x"ec4cfcc9ba975820");
            when 17045659 => data <= (x"c80adb6d2fba6458", x"9642f409ad26a8c3", x"00f2b66feb49023b", x"a54a771f109f5702", x"56baaa0430ccbb51", x"fec6a2ea17cf51c2", x"69ae69b26f2d8f48", x"f6265741f279d21d");
            when 6834828 => data <= (x"898fa7426dfcf42b", x"681810dffff38edd", x"f1e94e182c55599b", x"589d84c642497293", x"8ddc77f32e14275a", x"aa3d64660e7a8b8d", x"2b2da6526593d000", x"5075b29095bd0a55");
            when 9116949 => data <= (x"51c11b9a5c40576c", x"a0cda9d988194a7f", x"450a2e36464b2206", x"3dc9613d744ac6d5", x"e2148a8da326ec5e", x"4b3a6c71fea1ffdd", x"89bdb90fe8867d76", x"cca1dbbaba46b0fe");
            when 15264544 => data <= (x"8ebeb88ea6d17dba", x"018e201e8c46515d", x"525e745fd37b4911", x"5158f0ea3bb48f53", x"ca6d4b25fc692c5f", x"a4845b290a26e14f", x"5cbabdf9d0d8a9d8", x"2e819099870c38cf");
            when 26920513 => data <= (x"451fb55921c4e63b", x"a65aebdba2104b66", x"e4033b81549132c7", x"668043ef87e2c1c6", x"c9deb7154a67519c", x"b16784856c03a91b", x"1769736e00dc2d0b", x"4ed71e3b386a0c21");
            when 12588130 => data <= (x"22aba96fc5d12480", x"8d0d0c56d54966b9", x"0a6da49ac2b04f3b", x"5f68c95434f60585", x"f1a54bab0b591f98", x"bcaf40756f7c68e3", x"651c58c0fe0d710d", x"0f2ec8bc2857fd58");
            when 14951794 => data <= (x"b384d1eb8f638426", x"ffb9c6696c1aedbd", x"abc716a184166a05", x"69bb39a9590092e3", x"45ac787736c56a06", x"743788d6a4177007", x"515d2bde4110d736", x"95ce51dd4984ef46");
            when 18558600 => data <= (x"cf2279cc8eea9172", x"ac8a72f6f10bd049", x"1d6ab5e0eb1a7b22", x"6e988f6b051504c6", x"388197924b6b8e0d", x"27cf8caefda0aebe", x"8c758b1a4421529d", x"a1d69fbacfd6e20e");
            when 16496927 => data <= (x"d94d6fa09374cd33", x"f87879daac850106", x"754b7b816fba2270", x"4d8c2b652a2be8b7", x"80deba32baf33d86", x"ae77a3a0377fd6dd", x"bb9266ff651441bc", x"d053c8e835e5424a");
            when 22988697 => data <= (x"bcea4da5dc747247", x"7c229fd3104c01c6", x"21f9b7c052314575", x"9a9a3062d6ca3cef", x"348a67e7b3045c93", x"e319eadc17e83033", x"7ce5c7170d454f65", x"ad5ebd68de82fbdd");
            when 6282169 => data <= (x"9364e4cb86a84c86", x"629526e7e1a35e4d", x"bd48e4bcb546f44e", x"5ef42cc8303fefda", x"6f8d8e15e0d8d01e", x"109875ba7300bbbe", x"66c8a6d51da1e93b", x"0a179c05b1b55504");
            when 13281095 => data <= (x"7d9f6562b39f66e0", x"0511857e373864da", x"211f18020270d36d", x"8660fc3642b7face", x"ea5419353f8a3284", x"1baa37c94055e1c6", x"82a49561d8147b9d", x"2bdf2e1eae43b878");
            when 30981334 => data <= (x"12aa974fbd6e21f6", x"0e64ccfa1fbb7c83", x"9182a9cf61a8e226", x"ce10d088417e82de", x"859c74fca09b3cb2", x"77849fcb11629433", x"a2085119bc923928", x"925673a8d74300b3");
            when 10531604 => data <= (x"218065fa9d327128", x"77fbd751a02c2640", x"89c1d6db5cdd79cf", x"9cbf83e9a90c7909", x"8f5097004eeb9cbd", x"4cf22b5aa966da33", x"1a27ddf8d75f4d75", x"4b017dbc7ed1c412");
            when 6305956 => data <= (x"8a607ed6d77b7bf4", x"b4fb4886c0371ca9", x"c9b16596ff0e77da", x"883ef03a1434c54a", x"dfe0d2e3cac3d5d7", x"c16075dc34ae5c97", x"c64c7c9e1f7ed590", x"606dd13ddda106bc");
            when 13071507 => data <= (x"56a8f11ddc7d5666", x"2167acb23e2091b1", x"b5f88fae2a08a97f", x"4f9c3e30d3449781", x"4c34fa150f0eda1a", x"b07089bd3c5fd82c", x"76c67fa15d71c28c", x"c75da8a45bfb503d");
            when 26285084 => data <= (x"67bd33f294432b2f", x"f82c8558573f6fa1", x"88e516074f0c8a12", x"c76ebce190c10430", x"1478bbc8e8727f8c", x"ce84caa0d7f89e1d", x"8e69a748290d67b8", x"540639a0fa74e666");
            when 32664050 => data <= (x"858d7faff5113ec9", x"b29aab0a23eb8b58", x"b5dc04c944cad6a1", x"ca456c161aa806bb", x"0dc8a4958b8e792a", x"48ff2896749cd64c", x"e377e568bc268b9c", x"ec913b1cf767c6fa");
            when 14846842 => data <= (x"7daad2c58f120d42", x"d59a92a14bafbf78", x"f78fc9f057816201", x"bf6e5235c39f7edb", x"1e2fb3608a1d6c6a", x"bd830fe6bf515c3a", x"29b6e928b3de6f62", x"9e482b6407d36c47");
            when 27111540 => data <= (x"9a9e8013dcd139a8", x"2daea71b62cd3c5f", x"910c84a49ae70b3f", x"4c01f359d621a0c5", x"9a2fd3999cfa2f6e", x"27af74213ec0f317", x"c88c56184970e1de", x"998ed05e98d0c0f8");
            when 13121578 => data <= (x"db4e9bfadadf8354", x"1ac61de54c280344", x"ce5468309f55f75b", x"ef81f513b7e60c36", x"0080010ef802add6", x"4bfcdb0879866a6b", x"8194a7d8e75f8f46", x"b738f728d02ecb3f");
            when 3338185 => data <= (x"e2707b634a0d09f8", x"10226bca1d5a6239", x"0028f60ab035db8f", x"f6105326addb5f2e", x"a8e8c56c40fba9e6", x"45978e847d17707c", x"abe4017c2d734a27", x"9c02c8df0dd2077b");
            when 14949093 => data <= (x"4f588b5fe6baab6b", x"0e443143f6dcf3a6", x"6ee10781d4893462", x"f0ec1a19affe2b47", x"624fad032b8f8f59", x"cb7e1989efc3f490", x"cd5e2dc1d4189c4a", x"fc948a22d9528050");
            when 18785014 => data <= (x"b2ef74c715048d4f", x"70b986ed7a72e822", x"7b2976ca319f1e86", x"cc3feb2370e25d65", x"e84eb5f0179f6a95", x"6dabe108bd3973ac", x"ddefc496d3f2a720", x"8afed58791566111");
            when 8490406 => data <= (x"cb1e53217126e3da", x"e74363b296cda1e8", x"099acff2d7bd12d5", x"a3f245e3c6e6da51", x"12194760e560df7d", x"59f721ff2606153f", x"5e10bf0c80088875", x"83b81d1856250b30");
            when 4593328 => data <= (x"ec5aac0bfbee4a6c", x"51753f84b314a869", x"c9de193902fb351f", x"ac1e9d3adc6d5bf5", x"d25ef8481cc9b978", x"0168351dc854cf19", x"b44b2b42fc2fabc9", x"9b0dee9c26b2d0d8");
            when 29332988 => data <= (x"16083bdd6e0a640e", x"c13c88ac514e325e", x"a133e4e140c7cdf8", x"5af17088d1e566b9", x"22ae717b6f0de49f", x"1c492fb4962087f2", x"686b09cb588d46f7", x"6c128caaee8eca3e");
            when 29565553 => data <= (x"216d16415f48464b", x"8b64d5ab3bb75fa9", x"5aff617e13cee3bd", x"6e5fbb367cfbd38a", x"f006b85e1cb700b3", x"2c6f60fc9c212622", x"06997c6f06f65a24", x"b6aa10f524a896e3");
            when 21469142 => data <= (x"0cebdeb837b2e67b", x"fc350654a4c23014", x"ba240b78df0d4abb", x"63c60235ec26f0b4", x"a9ed0ac91922082a", x"246fc147b446c784", x"888b88b9de747b4f", x"8684b195b5ddbb9e");
            when 16483774 => data <= (x"28caaed4f030a25e", x"b820d7ccf9e8491e", x"4ae82de33657b6a8", x"2b524a05a400f8e2", x"e7b6e89df2287efc", x"349d257d28e51860", x"c10999e032b4bb55", x"da4cb4a1b48d790f");
            when 19055724 => data <= (x"184eb6c8f2d1313c", x"2abdedfbf75d0b41", x"5312df8d58f4aa0b", x"196f7d59339a7ae4", x"93c272c4ab44600b", x"4f5f95fc4871ce5a", x"7d00a9555ccfd000", x"3ddc9f5f5bb8b491");
            when 19627993 => data <= (x"5a5ec22a1f831c90", x"173717a3eb27526f", x"b862e86c487a88bd", x"960ee14f7d089f55", x"b758da41fdc465db", x"fd36a406f625404d", x"75588e84bc9c713e", x"f20e3a2d7b032777");
            when 13981389 => data <= (x"fef9fd2783f25172", x"693fd925a62d3962", x"80153f9d4a32cbe3", x"80073b8d648095cc", x"6a4ccbdfa78536a2", x"ab7a825e120a8893", x"7bc83eca60fe2654", x"094f9175161036e7");
            when 2028728 => data <= (x"580b0a1378bc3621", x"f68f468dcd884a5e", x"c4cea4924e1498e0", x"b77151657e6e623f", x"b3cad0bf549fb700", x"708355d66491c284", x"698f5cb02e304eaf", x"347a763e586a751e");
            when 15710317 => data <= (x"f77ee4b299706a79", x"b639cd6f80fae5a9", x"2b12cf691b0de64a", x"8c25e911e9c13680", x"c12647a96d413fa3", x"9db9b9db4a5f426f", x"25d7eb8c263a5de0", x"24968eaa40b0e80d");
            when 4519099 => data <= (x"e16abb20c608ca6d", x"cba73c12d88c7a4c", x"d50d08f88663d6d6", x"51f3f051ac429e0d", x"0961c0c33e72b6a5", x"c0fc4f829964b9d4", x"0de44fdcf18dbf34", x"c6d973acf557d462");
            when 5828909 => data <= (x"7d35fe673d0bf2e6", x"d478492856959d44", x"1c4cc0a3d229f2bb", x"1d5ad5c7e576f969", x"721724dc33a73441", x"d87c0a04ed09884f", x"15085432b8469841", x"9e768a559c17d246");
            when 23668536 => data <= (x"588be546002eb86c", x"9729df37fa868168", x"54f2af7071f055df", x"8aa5a8d421fc0250", x"b71371f99e35a1d8", x"e0c17029188b15cd", x"c52026ee78868166", x"a408e2802615a9bf");
            when 32193766 => data <= (x"dadf953f02f3544e", x"6ee36c7baf0a2d78", x"e767970d4ae2fe61", x"894db5d4167d124b", x"5a44c9c6196b81b4", x"e41946eda1c0d83f", x"05690f89ee425fb1", x"b9228ae2a4a15384");
            when 8184850 => data <= (x"19a06134c3c60d9f", x"37f9e4fd8276d70c", x"88fb5976b43175a2", x"82b98e713e4ba029", x"c2b64cba2c1892cd", x"3f2b2138a2c341c9", x"2d3d1037451d7e19", x"ecee4fc18df15612");
            when 15454197 => data <= (x"998399a25bb3f44f", x"8af213cd0f3f5514", x"4302ed1d1c28d569", x"d1d96aa18a7ad529", x"299a14316cf9219b", x"ba9a29d7ff524b06", x"328c3f6841133606", x"13536b5aa9c52681");
            when 13391593 => data <= (x"3ac2556b026fa9cb", x"07aa83b0dea666b8", x"db6bf93a9ae252d3", x"8b1d0dffee7a37d7", x"e9a2722e653a5f19", x"de6c8bdbb2770277", x"6392cd739b1087ab", x"0bd058b913a5221a");
            when 33112576 => data <= (x"0360c346702cba4b", x"7d8d6a65048dcbdd", x"0942cb02a5bd40b0", x"d7ec9b4294f89865", x"fe0eb3884dbf8ab7", x"a8e87e830933423a", x"c840976a8e97c2e3", x"1c7a571d5993e538");
            when 9975440 => data <= (x"5828449f563946bf", x"e8a209fa70aa7208", x"90e8ef89ca3cbf93", x"6bb795d21374d6ea", x"16cc386634f27382", x"8b3a6f99ce7aa93d", x"44a00c958cf67425", x"4fa82d3d876491ca");
            when 26106820 => data <= (x"bb5664c840e7e5c7", x"151b4b12bc7f25a0", x"37cf63774d21972c", x"8252bccbfddd5af8", x"93ceec6e8683c9da", x"10501d9c69a955ed", x"3486efd8f2f3da16", x"0e2d10e983910c0a");
            when 10382965 => data <= (x"0c4c4ea869a2f3e6", x"8c16a32517a7d3d9", x"be4558892123b89b", x"a5d215b40b10bad8", x"8fee4d211267fb9f", x"0d78aa3276635c4b", x"685e0e912bce6124", x"7f7f32e78e038133");
            when 10323856 => data <= (x"7636b90e53f356b6", x"e52c7b1a4a42e477", x"7458ca93f019e283", x"dfef6f8f9a685f18", x"89098f20ce2a5e73", x"a1eaf36abdc81405", x"2f2fdd3cb8d19c29", x"24d2b0ec83cdd48a");
            when 29132543 => data <= (x"60814e68f78922cb", x"c76704bc88c81e03", x"19477c1cfbb69064", x"47f7a03b3802cb44", x"33e54a8373e0a403", x"7c633fdde9207d1e", x"7ad3498957319311", x"901a7538b65beca8");
            when 3782025 => data <= (x"6f9afb18e85b80fe", x"2ca897ce51c81b7d", x"b76fca1bc0ed16ae", x"06bf1a96ac13d9ea", x"4520bad333abe9e0", x"4f2c7d7c13efb230", x"cbd5e3507fd2929d", x"d9aacd4410a30926");
            when 9747242 => data <= (x"ffc40b37220681c5", x"bcdaf6f6383b3e24", x"b9a6749c9966cdd9", x"c41bb6a0dd7862d6", x"e789fb31a85a05a7", x"3ecf8748b95f0b6a", x"8018aedb818b7be8", x"a7d4e5ee4d99eeb0");
            when 5526310 => data <= (x"2cf7c400790dbf19", x"d40e1f02b5d49c45", x"58aae824d27d7f56", x"9d6144df5ab67c58", x"dc76b0cdecee771f", x"d7a2af0b81694b77", x"8fc16bbec354a0a8", x"7d3918de8622f190");
            when 25634204 => data <= (x"9788c8d7bd5ebd6a", x"484602a1115d55c2", x"91e70b6637c14f76", x"d8814c63c9269443", x"c616806684f6769d", x"4b498ed431434b59", x"2bc26b414ad8b7d7", x"1a9b59902ad7d537");
            when 12665659 => data <= (x"029011dd7f14af5a", x"a2ffeb6ce38f98b0", x"837e4ef703a09bf6", x"2c2fc48462cbe617", x"faba430d2672528a", x"deb75a88d6d16d3c", x"88da9c31f1979684", x"bbbdb40040eb9371");
            when 30080198 => data <= (x"e668c26a62ca32a0", x"f66c857016d7a6d0", x"4865abf0b1c5dfd7", x"debd854ee000ef93", x"6efe298415348bc6", x"fe70d83f5b42a2a2", x"0f31b14f32a96021", x"c2b7a85535bcacf6");
            when 21394576 => data <= (x"7e30d94c776ff1d3", x"3ab847e2f879ab86", x"4d7aae001773d1b7", x"57563d688d2be69b", x"9dc3b43eda48a826", x"d26f3299a10c78cf", x"9aeccee5d22f8517", x"04aea0bb3a3eee6f");
            when 22160454 => data <= (x"9f4e75ad81127301", x"ca8d97d1203ed0fd", x"690b258c768de1b5", x"4addbb4309c5bc38", x"9c1b34c49fef9dce", x"d41bea22489b0f01", x"c94c4c0dbc62dc6e", x"98857d48f5b72dc9");
            when 27580763 => data <= (x"8c023cf59a4e54c1", x"4967d84d26a29439", x"e645a4afd3150016", x"3c512963cfe24304", x"13eafc189b8b61e7", x"ea61891a41df5567", x"3af20a0f7689a202", x"188dd7a09feecd14");
            when 32441320 => data <= (x"cdd83807ea091fec", x"ce1600bbec821afc", x"e9af990c2cbfad59", x"1416fc68ae4bda0b", x"509eec6beb935bc3", x"33f11d3ead6acb50", x"138bde5d54a3f68c", x"e71c5d2b57291498");
            when 5959138 => data <= (x"cb7529fdaf39d746", x"d8819ae0cfe7aeb9", x"db1b4ec15f8615c0", x"f3109cf6008765b0", x"63b4100aad6c8530", x"940d4685496c5932", x"3b9511d6c42d4ec0", x"8b3a309425f0db5a");
            when 13773595 => data <= (x"294a760bc9654b03", x"9d179f87e1f8daec", x"cc3e68535a08006e", x"075ec695c9e724e8", x"2d1318888710af5f", x"a1871cbf158b3554", x"c258b0da2b56d43a", x"0b9fdadf5221d76b");
            when 17995848 => data <= (x"4430c9961adebfc4", x"6e944e6d640cb8b9", x"6c070bd8dd95bd33", x"5e396dc29e1cea9d", x"1ff580bad82d6c43", x"37e9005ac3266ebf", x"8904761cd2ddd070", x"abe3add7d7519a51");
            when 29578198 => data <= (x"0b36927657269fd9", x"26bb34e210b3b220", x"c323cf0bedc0cde0", x"7c13ba078134b65a", x"b6e418ec1311657c", x"a12df52bd73c74e1", x"a5e300a73e35a7c2", x"cb99ab14d3c4b098");
            when 3161998 => data <= (x"4fecddb33a78b12a", x"5e1b280d68c74543", x"d2ab1f768e6f399d", x"2637c98cd4ea3932", x"2a96d2bcf41b7ef6", x"a46f5997262ec73c", x"af726c8ff5207430", x"419fdb334a4072b1");
            when 5521540 => data <= (x"7ed45b131ea24c27", x"8b51ed18aaf99e28", x"55f50822bfa02f3e", x"efb654424dbbd8f9", x"b7d4ed2f30cdca39", x"5c0ced8d99c86d0d", x"e85aff1575872665", x"3ba482e21ef59ea8");
            when 17829057 => data <= (x"a3a1bdb0f6749ed3", x"8c92cbf71dde07b3", x"3b7fdfc35906526b", x"0a51928b0477a4d6", x"0746dd9d4f75bb6e", x"2d9ed7a395736d03", x"4dd237759c7b6d91", x"39e7ee80c10075cf");
            when 10106457 => data <= (x"836a85e571458bc1", x"fe3ab817f032853d", x"df1758336a71a8c9", x"06bb3ac847385024", x"f5397e0410b2bc5c", x"936c343ec88fa3ab", x"d3b91270b6d6b7ed", x"e888a14b338054b2");
            when 14297789 => data <= (x"bca580458364f71b", x"c2f3d2595fe13222", x"50e543c85e91eb7d", x"e003d7e3f7bedf2b", x"d3deb383eed3f80e", x"bf1caacea3e6a4b0", x"c610225cb74b8fbe", x"e2fbfbbb4b07b4b5");
            when 27679176 => data <= (x"967f2cc85af2f63c", x"e161de66ab786b49", x"d417fc7425c74cfe", x"a770ca77f0113091", x"b48ff4eea1b23c33", x"fd82aae404021762", x"411b87375c0e1216", x"078dc99b833e22cc");
            when 17278073 => data <= (x"1457da35d60f27d0", x"6e63dcae04479dcd", x"a363a07684118cda", x"ce64ba8de317c2e7", x"abeaa002f1fc7088", x"76917462f65d0e83", x"d88ecd2ff8dc33c4", x"79678d1fd47cb2ae");
            when 28082963 => data <= (x"fe091c1e1d92ebbe", x"f91d429175bc8856", x"43ca1967ce6387bd", x"735e3dfe3dcf8b85", x"3c6b280c97593b31", x"5e8592ede6e0adbe", x"5c433e84a6789d16", x"d2f5ea1a89dc1fcc");
            when 7969769 => data <= (x"18fabe75cbe4599c", x"9b0c476ec729da6c", x"eee623df865f51c2", x"16e44acb308633c6", x"9e6967de4a49c36d", x"1584c57a3436bcac", x"b0f43468c490c699", x"46d98957d2b1d941");
            when 4829618 => data <= (x"a384a4502ef53fdf", x"f6e793672659d55f", x"4edc2f8f5eb5b782", x"e87bec090e8c7940", x"43cf877b64ff3c26", x"09f287135feaa28a", x"4f4aa1160ed1f91f", x"f2aafdcd437545a0");
            when 4748445 => data <= (x"ef9776d94407a74a", x"6cf1616508dac441", x"c87015c539777b10", x"b4b6a750d282894a", x"4e16b959e3638ac5", x"380e8e616838a459", x"385c75c6e94b381e", x"0f3824adddd7e83c");
            when 12786072 => data <= (x"45b33254b96d2b47", x"c982d601f95d3cd5", x"29941fc4c5d48925", x"f0615b633f24e6f9", x"a232697a9f3b722c", x"f301343c9abbc8e2", x"9653231d6afc1f03", x"122626fc0134bab4");
            when 31796330 => data <= (x"b4b8dc2c2e428af0", x"e0971bbccf2dc2a4", x"8538fef11d568611", x"6ddb68077b6dcc0b", x"43e52a7acd34e404", x"1365eb2816171e11", x"329de0516e9458d7", x"270e1391e99ebc83");
            when 14950015 => data <= (x"abb2acd0017b9e4a", x"f1525cf32e9bdeb0", x"5dcb5ce807eeb68d", x"a93770be2b15e6fa", x"8b62842f84a2ae6f", x"a5804b4169bf4dcf", x"9584fc4f6ffe196c", x"7a4a6d21f0e4ad7b");
            when 10152415 => data <= (x"29e089f037d58f80", x"e5acc701f1221096", x"55f9cee5a61ae638", x"2c8aca24f4343362", x"58864899286b4320", x"c4e45121059b162b", x"6ef1c5f539545730", x"23f6b860b1e01278");
            when 9695765 => data <= (x"6f5e4b186795764f", x"ba043aeab8b58201", x"3b2226f87e32c6ed", x"e271c00ade737ef7", x"9934a4a0202d853c", x"17c398122eaf62e4", x"d0f424824adb8e29", x"42a09eefe9c965b3");
            when 19717032 => data <= (x"b58059ecc28acb94", x"70f626206bd5fe05", x"8dda1bf4c27adbf6", x"00accb74daa1be22", x"163bb11e58591357", x"6df73bca2a15440b", x"7926f9a6b2365117", x"6ab88a182091d91d");
            when 473573 => data <= (x"a848b455087db8f4", x"a27eb5f17f7608f2", x"dde650b20ec8b330", x"b1cdda38402a75ba", x"d89176ad199f5135", x"84b042c7cf22b832", x"96ebd818073f5aec", x"d5c80862670528a5");
            when 19892481 => data <= (x"b0ee46670ae6e41c", x"b54cec6787d8ac8c", x"59b011c32fc16a12", x"29becfb653a5cdca", x"73e597c2bcf2759b", x"b34fab699e425e56", x"6ec36e0bd02a904c", x"0441061a3eb5c116");
            when 6968125 => data <= (x"9b9286af3fcf3276", x"bf9fd36655c4fb63", x"96eba802707d1261", x"e50f40a48174ede6", x"432f4d378eb3ae32", x"a6eab3be22b2c493", x"712f5aa847845cdd", x"573f5937f2771bd4");
            when 11892972 => data <= (x"4619369dc8dccdd8", x"96c2b988d0d61b37", x"0719b21504618056", x"96107b06a8901548", x"8c3d019bafa214a5", x"38782e6e48c796ab", x"73d1960c7b9aab72", x"a625fbbf38158c4e");
            when 16507365 => data <= (x"1ab6d85394738f42", x"fb145807a2385653", x"c24b4ce115a26e3a", x"aee88369c8cc080e", x"ecff8b6622047184", x"ab6b53f5863f7e26", x"23dd2b9770a560de", x"4c37c0e8279e151d");
            when 26749242 => data <= (x"c6711bcf07ae63dc", x"a76d4e9311759d80", x"40f735890dd22cfc", x"c1921758f18ab483", x"8f1ca08d45528488", x"0ed96bed59415c00", x"efd0b1c8fa27685a", x"566a91c99dc3aca6");
            when 8410541 => data <= (x"d099524475d5d41a", x"6c8fd8ec9334a7dc", x"c67ea7cf6f7d6498", x"934b3324f3b7bacd", x"c745af056c5c0ae8", x"1590ad36a2bd459f", x"dfa8496164563e86", x"ca1d671e88d9d048");
            when 11212414 => data <= (x"31c21bdead83b3e5", x"33c36ee78dc4184a", x"2deef2fa3c8e4d55", x"9aba81c5a444ed25", x"25fc4adedf51e35f", x"39cbead284471daf", x"066f6e8ac0554e4e", x"0e4553ed835b6164");
            when 12030313 => data <= (x"eba00ee484c503d8", x"f5d3b218f70fe1b3", x"c5098358f76fcca8", x"fc82f41be2bd905c", x"2f198fe7e27717c3", x"b4522f1b523ae2af", x"4d61e52ca074611b", x"32b2bfadb1cc9cd7");
            when 2430537 => data <= (x"77c4dfb944ea2095", x"5682c8f23956b8f2", x"b911d96530e4c78e", x"7ff74d4d34bbef8d", x"7d778b05f91fc215", x"05d94336e9ea282b", x"5120402237044e17", x"85593d2ba870d225");
            when 20718215 => data <= (x"4ea476b17b2b52e0", x"a4169fb92febe447", x"ff536052d10871c6", x"698d6ecf0cd920aa", x"63ae87a50b28b8d9", x"dce27ba1d71ee57e", x"e3b3dfbee36a2ba8", x"13bd85df15e2963d");
            when 1940350 => data <= (x"a7664cc6a69b4956", x"60ab7dee6db9ebf6", x"62ac49fec93c5b9b", x"fa7e42aa9fa551d4", x"663b52b8750d08f4", x"5e3ca3da819fc2df", x"d2625ed7adc148a8", x"650fe33e8593f3c7");
            when 32157643 => data <= (x"252ad5b9eae2652d", x"573ea41229dc7590", x"2b4f73b2bed90790", x"70303cf961d16daf", x"0e301db7de8a5f72", x"94c0c8569f91d6a3", x"cfc64514e0fa0c67", x"7f3d9d64accacecd");
            when 26989983 => data <= (x"eac33464efa6f329", x"8c85e65862900402", x"6c8100ed7b00fb38", x"612f8c6468004cdb", x"3efc78a5d27414a6", x"ff50a6dae4fcecef", x"0cefac51af720f60", x"aa4dcf8e81526de3");
            when 4358829 => data <= (x"e28c56c413233794", x"daefbe1bb71f4197", x"7942d0a80278d14b", x"0f5a7a235dc92362", x"0a369551d2b9f962", x"43fef06d0d0754f1", x"b77fe2260aeea52a", x"708536bf0ba44929");
            when 13906758 => data <= (x"ffe2f6858c2a91f2", x"4a220485b315b6c3", x"60e535cecf6b7849", x"70297509e7cc8964", x"8cf7b8622e388b98", x"7e57b49134da943a", x"e160b298cf9b4a08", x"ef4a599b2e6d21db");
            when 1144088 => data <= (x"d5c4582dee373980", x"4c21358e957b84b7", x"d864afbeba7259c7", x"ff55959744521ee9", x"76d4631cc6c99dbe", x"b6be7853028e629c", x"0cca893b3a7ec4c9", x"98ea80e5cbcd7dcc");
            when 15506210 => data <= (x"2f82902d7385dc86", x"d967826feb5dead8", x"10b0e5069403e290", x"2ab58e016e30be2c", x"fe401c19fab12a8c", x"de69b3bcc84aca3c", x"4d81053db2451bd7", x"913deceddcbb7c6a");
            when 29194911 => data <= (x"953a214e3add29d1", x"974803d0eb56cb4a", x"b52431dba6f937de", x"07600cfc618ef3c8", x"7bfc4400ad934da6", x"fad45814495ab261", x"acd35763764b78c9", x"0d6d161a66a8d2ef");
            when 14784998 => data <= (x"02ddbcb953db1a18", x"bed4c86214830fb1", x"0a100d8263b29ef4", x"d8ffba60ac214e30", x"74e9d2244fcbac2a", x"617308149f0d1bc3", x"85e988fd67ff01a1", x"5fa33fa0f39ef385");
            when 26878787 => data <= (x"919c9c942c643516", x"b492a8c2a63a73b3", x"07ff5873cfdcfaa4", x"cb7c2475d8e984a9", x"04b99a3fdcfcfc85", x"a3683abe10ff11ef", x"1b00ccdce7d22887", x"ae260658343d6b72");
            when 19234658 => data <= (x"b4acc7fb736c30a2", x"2ea083731cb1012c", x"1bd511f628ab77f1", x"f246c2951e4835fb", x"201b9704ee1ddfe2", x"e9ecb49bdcc31a55", x"45e5820de8fcd526", x"1b57f2749f4e200f");
            when 33105476 => data <= (x"e3813d64af072232", x"b7fa92f5393753bc", x"a707d638fd4a4833", x"9641f0714e8c24ed", x"2b12f2bf4bf1264b", x"530b75f131b912b3", x"808ed9266d54b3b8", x"1808b7dca4150c42");
            when 16736324 => data <= (x"c59383a7d5c644c0", x"51083c28e2dc789a", x"90957d364ce10b1f", x"bd1f46803a0d9549", x"71150dcc5dbd4c5f", x"c9044c583502cd2f", x"ea330e8571c6b073", x"0d7898b5e4155173");
            when 13532247 => data <= (x"7833fc3ec959e77f", x"11768501348e81ee", x"961d4df61e7208ec", x"a7c1771616bc0396", x"36f241d8c3ed677c", x"e5df6e6057d45d77", x"373915ba7908fe0e", x"eac5496054c8ef6a");
            when 26369777 => data <= (x"d97797986f6e5ab2", x"cee3b2dfe21ff984", x"8f6fc20eab0c57c6", x"7b0f013f72adf124", x"5fe6c3107af655bd", x"456066d1a10c586d", x"5ecaea5d2a82fd93", x"af87d022de3a5d2a");
            when 3827324 => data <= (x"c3e8136037638d51", x"44d81ab4e87502c7", x"f764603b0851e9a5", x"cff93289d4f06c1e", x"d92ab3f9a03db1dc", x"f979a0a24b8f1290", x"9151da5c51e9768f", x"3bdea899bc78ebd2");
            when 2701194 => data <= (x"08cd03f340244a39", x"b579ba6c14083778", x"d54389c142217ec3", x"ac983f6076e01b91", x"06857c78a9dde249", x"1ca4f33301896c7a", x"7d5cd72d86f39fef", x"52d2b40329ba9c24");
            when 17371671 => data <= (x"213499c277daa0dd", x"af876c7cf269e6f6", x"2f3ee4c83f40729f", x"9d1a01be9edd3b86", x"b003a67c9c83ea3c", x"c1728348e355c8dd", x"16d57f9f01e69bfe", x"3095b71cd69eb98d");
            when 23707210 => data <= (x"9118c870beef1d43", x"29bc1de55d4bb641", x"2336186483a0cafa", x"0e5944a76dd93c7c", x"1799da208208933f", x"94e10aa68fec4534", x"cd4548724367ee9a", x"727ee51fe7f571d9");
            when 16473146 => data <= (x"d0fcfc71f1c0ddf1", x"6f75b5b561207a18", x"6066586d6e517c03", x"8bf3407f18ee3acc", x"743bd81f3c70f173", x"f06a70aa4d247232", x"b84ef7323b148e62", x"f4310d7f3f740914");
            when 10356556 => data <= (x"3fbec914a23bebe1", x"49f9ffbe700ea96b", x"7fed13d5368e4553", x"95e4641e189e4b6f", x"7d42c65697fee554", x"90216e27251d6056", x"2640986561770c9c", x"cb3a80c8a5b8c528");
            when 300790 => data <= (x"8918e29f2d365482", x"ff151e364865ef7f", x"e2f7cda91992f65c", x"158b6b15bc86193c", x"a50deb39ec02c05d", x"670d8cc9033b4e8c", x"c016fc4a558d4ca3", x"837bd5850f9bb092");
            when 26392891 => data <= (x"a0c1eec3e4a57acc", x"b7327e7c26702f6c", x"d974abeae484fc49", x"e5043986eefc366e", x"7aa9ac82398ae12f", x"c71eca41575fa98f", x"af700035324fc75f", x"db6681cdbec39966");
            when 6313291 => data <= (x"4d04bb37bd18a58b", x"d606c3f0b4b18959", x"76ad8292cd8f7b6b", x"97f2d680df45191f", x"260c018624432842", x"4dc9b75b7ea84fee", x"819f0a45c14a6783", x"070ff3a7a97583e0");
            when 5821784 => data <= (x"8726ef1dc5c81f7f", x"9acfdc4eb550a47c", x"09989fd1aa3f0365", x"35be1fba859d6ec5", x"597349eb0b185d99", x"3d73918edeba6523", x"b8b570bf1c198ad4", x"a2920a4c364592e9");
            when 31704737 => data <= (x"df43074226f23469", x"ff3571ca0e097e08", x"cce3959fa1a4c971", x"d3655a3e3353cda3", x"cb629636e0d12c42", x"6c1c90f56e798a8b", x"fe1f676867f3f66c", x"998221a02a7420f5");
            when 1340418 => data <= (x"39378d9e5fbe948c", x"5c6d39651528d741", x"78b3128e535515b1", x"ba618c4cd72b9b12", x"80ef3a40dc4023bb", x"c34e01018486a24f", x"b1457c6111f7302a", x"239073d33eb43728");
            when 24053048 => data <= (x"5fa29cb91c28a733", x"1c7271d07dbd25b8", x"118b9c1b86f229ff", x"965577dd7bbdf168", x"8f0c6610851fd76b", x"7ca3d5a1074e785e", x"ed07282bdd186b4e", x"4d922c9c827fa1c6");
            when 29102051 => data <= (x"3647c50802780f1f", x"ed38a9fe3a5fdb3e", x"00c81b549314c54d", x"b876fcd3f025ba03", x"69ee807c5f3bec1b", x"88e22894d5bca9f2", x"924d05e2128c3de0", x"4fd8612b8bcb42d3");
            when 7298306 => data <= (x"b3a303c629046562", x"690bd22a5f086fc0", x"e203d4de966565a0", x"417d96db9626d43b", x"f632f07e5ed5b58a", x"bbefb2c8fcfb219d", x"546cdffd1961f9a4", x"11a189eb713e4dd0");
            when 14098594 => data <= (x"c5d6efc9a911ab20", x"ebdc464a62101db4", x"7fa8959d75e9448d", x"8cb62cf05524653c", x"2ee8c0332ff95569", x"895dbb4af26ffe1f", x"92c15de073157a2d", x"3dc6f6c0367fef21");
            when 8618097 => data <= (x"5e19a20c77e1ac99", x"16cb927450916e49", x"645d866ccd1ce859", x"87888d4c82960bf7", x"c0f08c0768a353ba", x"94689209f7fd7475", x"7a4be695ceb39e97", x"668359c3cb7e5e53");
            when 10767859 => data <= (x"293a838d42ba6897", x"2f37d73848a25555", x"04307b8bd4158148", x"49112d93b382a69d", x"bfccdd3b0c9034f9", x"04798454b36ab493", x"8e1bd830bfc0dcbc", x"83f6e6559f648554");
            when 3037982 => data <= (x"290ff9616d9edd4f", x"cb93d9a8a6218f8f", x"06f5087e8276753c", x"6f81a12c245d01fb", x"9acb31fa2ea7ef2e", x"f5ff7ecbcd66994e", x"79424a1878e58edb", x"bef9a78e5ca1c035");
            when 33380941 => data <= (x"a5ae293db5a59621", x"39793ef4425f6032", x"ad33ff064bc339cf", x"8bdff88807215948", x"6b08b18666fc6a02", x"9f24082dcc586bf7", x"a0045f28c5f98196", x"2e7d52d87898ec48");
            when 10070925 => data <= (x"c7edbd71c6ab50a7", x"d8ffb57b0f4e9cb1", x"ec0a53010953b75f", x"c844486a8ea0a25b", x"13baf12ef9de90c2", x"58c210fc7462f1fe", x"e0f0c8a8f1fed43b", x"27d64ba0d4c04121");
            when 4378282 => data <= (x"fdcbae3eaa1e3a3c", x"af352e4ee8ba7b7d", x"f20133f3d1747bf7", x"f22b07b961446f82", x"b707c3d048d9ea47", x"cc84099305391064", x"c94158fd32beadc6", x"aa6f826e6e0166c5");
            when 13084774 => data <= (x"56f45e8639ae1b97", x"50df9ff6e5a037a8", x"14ff95d79b2f9744", x"714cc4cb4398f5f0", x"b8e59c4ffda207e4", x"f8916ad936586bd6", x"03777fdc533766b2", x"08cdb43e7b52aae6");
            when 16445044 => data <= (x"385f5778d00a7cf6", x"84ec21301e957c36", x"edfdac95e3e0862e", x"6cdcafe66b8b1640", x"352f25f7874225c8", x"05f2271cd84b8b14", x"9e82b104356ff82e", x"bba03dd1009b299e");
            when 9238218 => data <= (x"73469a9fc4b77e7c", x"2baf9a980ef4f246", x"7c1ea7f857af7ec1", x"80ed15a9ca4dce2a", x"8aae5176b92f6f30", x"1e8e72e673d34cbe", x"59f4057170b3e53e", x"0a6b32c1c6772b12");
            when 31469667 => data <= (x"970ed6bfe3430373", x"75c8b488e945af91", x"b1c45cd91e06dd66", x"1d83ad3fe3ada0fd", x"8d8a2f1bbdd11523", x"6f638564f72f6ec1", x"da06db7323ce1dac", x"7206663734790d7c");
            when 3621477 => data <= (x"091871d2a3d71aee", x"be86ca81639814d4", x"de06f3619a81a20a", x"0335e2d81c1aa106", x"3412de95c6f04bc1", x"52e0a0caa44faccf", x"bdd89a4551809ec5", x"04a24daa648961f7");
            when 25373501 => data <= (x"93422e109e9c3d74", x"a6088b5178d8c28d", x"973f65a1bad9ef5d", x"d08628fa58078e42", x"219cea395123787a", x"9e0676ea7ca594b4", x"41d0a262465a6fd8", x"62851b37a61f8247");
            when 19615307 => data <= (x"b69eefad73b821e6", x"a2b894a3d22c0698", x"95dc577a2d11b69b", x"9a5fe03a3cbf3535", x"a7b518dc00b17bde", x"b7ab7edc007f1945", x"b091f5a3a8b870bd", x"60916d2f2510ad53");
            when 26314597 => data <= (x"e28c51e8051a2d60", x"87d254a90ddef257", x"8eaf0f626492a997", x"fa089cdc9c03c07c", x"c899aa08cbb6a70a", x"05dbc82bb0291090", x"cdd8c594893f2d51", x"d6b53d73d97955fb");
            when 31427724 => data <= (x"12ac48219ab78205", x"bfbb3cf73f6a2197", x"7004f874c4d85ca2", x"74e05cbd1b5c95d4", x"e89f11e6ed2c0a14", x"a87bb3c76caed331", x"4518fa4cc5ab8fe2", x"8c355aa7cb583439");
            when 22570096 => data <= (x"69f6d1d751086170", x"26d8df5a6430482f", x"84b75984f71859bf", x"c13eca1032b4f870", x"7f326ae20dd52e57", x"b6b4b4ade5660791", x"6a9af47752a0a3a6", x"752513e7a3b3ecf2");
            when 18179654 => data <= (x"a8c7653d5049bca1", x"ff75812e69e5795c", x"e14da678bc198baf", x"7f4066b39f9d2de7", x"ea7caeb8b3d1c4e3", x"fa8e820febfa6def", x"440346dcd74a93b3", x"7161997b12265933");
            when 15543584 => data <= (x"436cc75e97194bdc", x"590b7e50d093df9a", x"cf3bff922826bb29", x"1da486af928f099b", x"06e0e666cba6c50e", x"3fa2ffceb19b6316", x"927e3b3fb974264c", x"2b8e8945b8de1268");
            when 31532699 => data <= (x"aaa3cf34bfa5a9d3", x"019f3fd81131f880", x"8345fb2cf9210bb8", x"6b70e1b3691e8dff", x"b16800993e372b3d", x"648bc9eb13de9272", x"0e2b7c40c3bfdc1a", x"65650419d4dd285a");
            when 4796779 => data <= (x"d66c55304cde275f", x"e92b08824b678604", x"26c08c1cd0d889a0", x"0b40f1c0fdf782c5", x"471926c3fc16ae79", x"f3c0729ec48e7904", x"df38f4f835a6d446", x"24002f26966204fb");
            when 13387786 => data <= (x"de6dedec123c6c82", x"82f75e4796383b26", x"cceb01da963472d2", x"c51ee4b8dc64bbc9", x"82975723f2fdf939", x"f2ba23adc1d3edfb", x"662f1d2be520b95a", x"61141f3c8330d3b5");
            when 14534787 => data <= (x"c2c6ab3324236168", x"8c77906062449ce0", x"167cf460d36ff375", x"ce3fb6e3d651e88e", x"c232aa7f7fb72a6b", x"0c142c90f6f201aa", x"ece766f5bfb08e5e", x"c0c79322bef20c2f");
            when 13089184 => data <= (x"c324ffcafd6de19c", x"23181f431c014055", x"124c566b0c61ed57", x"7e19df94ec16bf4a", x"2415da9a44906dc3", x"eb9dd7ddee251342", x"1e7063475dfc2146", x"2ac7b73a521b5ff9");
            when 15309301 => data <= (x"4cf379e2bff97d05", x"29ea45dbe3836258", x"88e7d671aaa80382", x"a2af3c5f50ec7286", x"92dda1c1cb4ab46d", x"28c1d3396792be4c", x"9eab53bbeb60dad9", x"b74693f7f2a39f9c");
            when 15151355 => data <= (x"f93f7e0342dabc18", x"97f9fe1721dfaeb5", x"afec6d622d3a29e8", x"06fd14ab4727da60", x"6e49422b900b71d9", x"e6e81b826a22ff4c", x"711253c82a8228e0", x"206aaf8aa3d1e8ee");
            when 1388897 => data <= (x"018c5d61f1bc4c82", x"1cf0b194aeedbc4e", x"f55a3c0de1893ba0", x"25122027e14ec6b0", x"b52a0d5e18cf7c33", x"34079f70c7118e02", x"f4ae5909bc2b5f9a", x"735218669cb5cd9f");
            when 18186304 => data <= (x"2e8c93a86a15d291", x"04760dbef3f9a620", x"d9d283caa1aa9a3c", x"595cd4d2687c1fa4", x"3daac379d41016e6", x"57d2a6e6ebf5d015", x"a5c9552392579312", x"3a7fa230b69026f3");
            when 28646330 => data <= (x"f0371803ec8cf979", x"5b2ea614cc14560e", x"2ad0cf0fb8aad849", x"3aada9054ece3a95", x"cc828bb84c19f87c", x"5da0f0fa6a15528d", x"d695625767992b4e", x"5950d53e1477b2a7");
            when 945745 => data <= (x"4e16fe662ebe8d3f", x"4ebc8e290a9ac810", x"b011b8abfa6c6827", x"d337467b0ed1fe55", x"f2f51970a1559eca", x"e9a26fa3f0e30c83", x"3f3fd7fb0accac53", x"da59f86b4c01dfbb");
            when 7982842 => data <= (x"5de2fcfc7f589324", x"71fa5e6f3b18dbc9", x"59d9101f92e0d7d9", x"deb53879ecafe824", x"77f432181547f365", x"fecee1c1605250fb", x"0467ac74a1e23e8d", x"7d64432d91b88722");
            when 6526098 => data <= (x"7f001642cc65e47c", x"a7a284be7ce9d177", x"1f3e75a96537658f", x"fce55138448c67fa", x"4729495fe6d12cb8", x"ebd236c9bc92031b", x"af533c25636aea60", x"69df93ae8c7e01d6");
            when 32184770 => data <= (x"6430e869aa68b083", x"f113ebfe8d34f233", x"afe74d324c57ea8a", x"d10651a983c4930e", x"0c1ee1e619db9a9f", x"47233bea7c4f10f8", x"7afa2209692b69a8", x"b9d25c176ea6e512");
            when 1980597 => data <= (x"4b427e4478b5b88b", x"4c931c7902e00f66", x"147859b96d55f35e", x"aac46859569e0df8", x"f9d6cbd47ebe855c", x"932d22c0f5f97277", x"4b6723ae4aa8c048", x"52d40c5958b18609");
            when 8548147 => data <= (x"3be7e71a1e3c877c", x"de6bb6d0e7fc718c", x"a95db60d9acba33d", x"6472d3e2531f382a", x"01f7df74da634e53", x"d2bdf32c9c2ee325", x"f04271d3dd90da8b", x"bfc9884e79f69524");
            when 2252101 => data <= (x"585a76a43d24deda", x"9090b489e5ea516b", x"cc741123c4ed1911", x"f27aa2837ca6a1ec", x"3535818fea28eb01", x"00022fe00d417818", x"65140612af73a918", x"f3bcda40a357ba28");
            when 595597 => data <= (x"499cfa819bb25210", x"bf95f718ecd73d2e", x"5c016e83e0e8d825", x"8bded801e0901fde", x"6be905acf3c5ddb3", x"a9c460df3d7af426", x"4147c2333ee1ab88", x"bf60bab9af9b7aac");
            when 14500831 => data <= (x"1f7413b4b9743285", x"0b738b4178741f33", x"1ad52173d38aee13", x"61e0a27621ea33ea", x"9c9b4a2e569f1a8a", x"399ad63bf07b298a", x"55a3b37562f6679e", x"925b0df885fd4adf");
            when 7298586 => data <= (x"70714b0e334cc402", x"22198c8d23f094cf", x"4b2901d2f526b385", x"d8cda68207685d64", x"cbadb8484b26957e", x"2129867efe9506df", x"01c54e34c6c27682", x"2a9693b954ddf2ed");
            when 15444685 => data <= (x"59c919cd75fbfc6b", x"98ca345576c21938", x"a9602c0247abaedf", x"f8b9c0d5fe641346", x"b346f8297cf32799", x"a8b4a9f485b2f6bf", x"a6db8fb32aec555a", x"91fc7d69bc3b3cf7");
            when 12303834 => data <= (x"10576f60840de36e", x"401c63c0ac14cae7", x"273044985eaed992", x"77e4ed690646530a", x"b62d2aa28c5eb482", x"34d301e5bff68d34", x"bc3d2fe9dbf44bfe", x"180bb04a627b537d");
            when 15826317 => data <= (x"cf58d7da45c632a9", x"8ae616b297444727", x"5d755617b07c5e19", x"a6108ce9f63b1f5b", x"898ce30379ac4350", x"0fba1fc6947174b5", x"d0a9b2cb22c5e922", x"440f6b2ec05643df");
            when 4323388 => data <= (x"d310195819147a25", x"c8770100342e536f", x"ac86e32675feb164", x"65d48c2d4b5151b6", x"06d0cc2afe39d6a6", x"e0b2ca090a36a697", x"2bacf8d64f52e1de", x"c202d5ee149c5ee8");
            when 19310865 => data <= (x"8e885cfa15da6741", x"e633b5ff6b11e551", x"939e0e513acec73c", x"43c9a25ab8be6728", x"4a13bd2cca08cbae", x"ace398d4eaacd924", x"ae298dbd3e4a2ebc", x"3a15c56210bb5455");
            when 29904544 => data <= (x"ad47443e701bacc8", x"404221fa8be08ab5", x"017d3403ee318df5", x"389ed781e9a811ee", x"f3d6a1eee983a662", x"68d3c2434a78e568", x"2055265e4ab2024a", x"e944729c2c8fa00c");
            when 18103147 => data <= (x"c195fb1c4a94d7df", x"5da943473f1ed768", x"f6323e7ef83c73ad", x"392023022c2fc3e0", x"75b12cc144ec5dd0", x"4094144a47869afb", x"c50022074a705609", x"3f8170f4c3b7b5e2");
            when 26909164 => data <= (x"90edb8a2d89b1e3e", x"2186f79c2251a059", x"db0e59d366a701ff", x"3898ef7f1de9c53a", x"b916223c580eac4b", x"d0d6c8851a81c753", x"918ac21460180cbd", x"54c1f6ed741fc1ea");
            when 20515598 => data <= (x"efd43aa961081e54", x"3998a94e794c16bc", x"b4b0dc67322fe4ec", x"802f75c383bb978e", x"1093fa0e86ccad46", x"94322d9ae317657b", x"a6177ce0fe9fe3d7", x"30803f3200a14f6d");
            when 493861 => data <= (x"1dfb51ad4213d1fb", x"00be331f4948dbfe", x"ab40d42395188500", x"dc2b59086fde15f4", x"1198268d334f777f", x"c5bb63fc2197180d", x"facc102c8160ca12", x"c96894d686f13f9d");
            when 3114372 => data <= (x"2ca80d1327227e36", x"6a38cbbe23aea5b7", x"fa6edaebb9b1b2c1", x"3a9abe73e8876597", x"387c6538f7e12c91", x"f8f5e6d46f22c2d1", x"67a4d9a237c5db71", x"64e99c29def95047");
            when 31259728 => data <= (x"897d8b02fc215ead", x"7ca82682d1560b0d", x"e3aee212ca307da7", x"999cbac76a6f4eaf", x"ffac9167c08dc4bc", x"0bf397aff0a5a855", x"c08c1284f4bc506e", x"69744d5e26ad41ee");
            when 15918775 => data <= (x"528d76737a923a30", x"ac393c755787df2a", x"05310a5cfaef012d", x"10a49e9bbf2f9090", x"86ebccfa20332e89", x"f9f0d97fcaad0faf", x"00aa2ff44c0d4106", x"d33822a4ba69147f");
            when 535811 => data <= (x"3909697f14efef8b", x"8231d297370c6e4f", x"84f80d87970fd694", x"c8570bf8cd78bbfb", x"306679d7537ac568", x"f450d2c38d7903f1", x"d963aaa3b1ed03d6", x"583c01a678922f2e");
            when 26704533 => data <= (x"f414fd59f8b01d2c", x"5291566d079a655f", x"c805b5090e4ea289", x"20827f373589d9e1", x"5e29241ff12f2bde", x"6f24e025c425aaa9", x"36b949b17ccd9f5c", x"e00065ccbb4d7f4e");
            when 2558360 => data <= (x"572d91f1b3252f81", x"06a81b271164a240", x"bfc85b71edd690ff", x"f3bff34c5fca1257", x"256eab441f9dca30", x"8686308496d9affd", x"af894fdcfb4405a8", x"05dce6dd0468d33e");
            when 12007284 => data <= (x"a1fc1a73eba7c4f1", x"68ef4f398f9ed3f1", x"bad8ae89c6bc9852", x"5927fdee02db5c0b", x"5b50cf5c5eb56de0", x"43cb5ba492ccd0c0", x"8303f0d1f4812f3d", x"a1f04c1091bc7979");
            when 10026878 => data <= (x"ac5b5912fdd7fca3", x"186dbdacea2698dd", x"9fafd9b697ed6817", x"b0e13778a017b4a9", x"755ddf82dc78c565", x"7f0a1075e7cf5a26", x"f8a29a27fc49462e", x"6934224597f52433");
            when 3338878 => data <= (x"28219c189ec54050", x"1d805373ccf07ae3", x"8586869bf9c72f01", x"d2439d2a6780cf7b", x"5a7fcd9ace34c36e", x"8d3a798480f66cfe", x"4ad793a37b08d671", x"be29d70070a32310");
            when 24998050 => data <= (x"0df37158f822a5ba", x"f199e47dd36044ef", x"3ad3dc8af23ec142", x"93de7642d7e41481", x"1eb4d9ed3a280709", x"86d8a091faca5f22", x"cf6985fb2affae60", x"b0f78f6507cbfeaf");
            when 6145472 => data <= (x"c53133de44e107b7", x"636b75df03bcd889", x"3da6472b747b7b71", x"c75e8f5dd0c49aad", x"9d1098da845e3630", x"a1cf8279bff8478d", x"d5037ea47264c3fd", x"08e1a0aef175e49b");
            when 11932902 => data <= (x"8bc0593576415cc8", x"5ee422f2c8718b9f", x"a7f976bae45b5801", x"1043b5a2d5e5f1a9", x"f855274c947f3e28", x"e30595fa42d6da67", x"f1eac87a128774bd", x"8eaefa22b88e33b9");
            when 24613991 => data <= (x"8ebcfcc1afc77a56", x"93793a439ac699a3", x"c57b3f4a4c3c8a9f", x"ddf2434a0bab59fc", x"2fe3aef4b236eecd", x"9842448e46aaa7ce", x"a5fad1b7c2db7ba4", x"94b94bb73c533fed");
            when 29053676 => data <= (x"133fb7a2a1486452", x"6ab79e24883ebc51", x"073980f7b992106c", x"e851c7150eabcedb", x"e2169776ecbf4637", x"75cbdb081ec34ea8", x"e397aefb67a3b1d6", x"4d078e0ae40ef582");
            when 25550569 => data <= (x"1283f46ff0d3b2e4", x"c0c39cc32c3f33f3", x"2f25f155613a0815", x"837665bf12f5069f", x"171549e6459d4c7e", x"1b210d29e6be5d58", x"12cd4ccd334c08bc", x"a64e44a41244ae0f");
            when 9725688 => data <= (x"125e1941b205152e", x"86848e87f8a83c90", x"3ced25b33ae35848", x"9b254af640797b31", x"9fe3cb65c0290434", x"48faab241c87d195", x"8df262307d9c30bc", x"2ed1b48ee4d0d3d8");
            when 29226336 => data <= (x"a379d7394423b62c", x"84d4db7cc62346ee", x"8898301b19f36577", x"67b681c6d58eb90b", x"53c06af6d0d7447f", x"52d804cfa3dc408c", x"a066a96941105c41", x"9543c6e22f7793f2");
            when 17862882 => data <= (x"1d24ae1751718caf", x"06fea0bb12a22638", x"8e25ea3023083e2e", x"83779b133df856ca", x"9c48e3587ba6d34a", x"0e76d4020a2aa5bc", x"fbc836ef51d09873", x"a94e952afda549b9");
            when 30949390 => data <= (x"b161804487d18282", x"b135346a7ce3e7b9", x"e13a72fb10593889", x"b6776953dada134c", x"d63c4aa3dbda8106", x"2d64761aeba1fa31", x"8f7a4f4f8d46fbaf", x"eab03a2aeae9e1c6");
            when 21299708 => data <= (x"77e6adbab99fe279", x"a4c1fc20f0a90134", x"fc32780e479a0c26", x"a907e6f09b99593b", x"1dd22b3945534c71", x"b88fbbb3bb4dd5c9", x"24c948414c66b9a8", x"06514c53cadfef38");
            when 30110317 => data <= (x"4f3db700a20c5e41", x"102c9fe061e9cc73", x"fc942c7fc9a6fae0", x"fccd15703e31bd7c", x"c8964648bd8bd8e5", x"e53cc29e6b33a604", x"e13af1a9ebca5a0d", x"7388699a2f508939");
            when 8135687 => data <= (x"0a84a90a06b243fb", x"abe887c614bf2c3f", x"66286e2a2b296747", x"ef2930a1bc9a3043", x"57ed35044f83bd92", x"c8e76db9348f6f6c", x"2baf9c9204746e55", x"60c2d34f7baa3a95");
            when 1613135 => data <= (x"57835cac08f754e3", x"564b4f450ef01ba2", x"2d4997db3e0bfced", x"cd9edce374c81e09", x"9d829bb5f96e12ea", x"3a94514b432885d5", x"d9f95f1e7e2a500c", x"8918bdcf3a1a12f4");
            when 7821487 => data <= (x"82f5b630f34b59f6", x"2e463e1b1e77e8e3", x"a30af8832748a5e9", x"d8b37bf674a19ce9", x"d0a7285462d03c56", x"7c3218afe5f5f5d4", x"c1de4b2ae2495687", x"725c4629d2106b43");
            when 3649300 => data <= (x"8084a871f39b992e", x"bb7ee293a18dc3e4", x"5308bef3ea4c8a3c", x"d9799fe13485fc64", x"e80fc7122365466a", x"e0dba388316ecba2", x"c593f566b72c8d0a", x"8cd849b52fb7111f");
            when 9741151 => data <= (x"00f6da7ed603ce70", x"0513d8e148f03f8d", x"6a65dbc42fdd5fbd", x"9034257900bb3901", x"0b63b836802e7f85", x"7731fdfe21786dfe", x"10b77ff232499473", x"609e7798792a39df");
            when 2501023 => data <= (x"511462e154b1566b", x"18da41ea21f6e291", x"20e8c4850f72cf54", x"4c03774fda3f9303", x"e38b55f3e93818f4", x"32219a49378d1236", x"a6f2dd2edbd0c7ce", x"c4f71b9e694fd1f6");
            when 19543191 => data <= (x"490f9be4a283c0f0", x"d415ad4da98b0265", x"a77815b0742b0465", x"442473596cc4d256", x"8f70d894a49be30d", x"b96face0e53f222d", x"ee205af61a05b9db", x"0bcfae88d3dc4ef4");
            when 1104473 => data <= (x"691af9e102f84dcb", x"1cf09681f07c3818", x"f48420c99c8d6213", x"0b11f9484c6c116d", x"8df873074e753101", x"a595955215d8c6d5", x"89fc04ebc1ca9d73", x"83c998265b31e2c2");
            when 4936789 => data <= (x"dedc6334e7167754", x"393576a77d9f10de", x"37eb7ac1f54c18f3", x"16c15dca9b3ccc25", x"7e06d17682234df9", x"e691441ca5bd5253", x"fdac9f303cf5dfbe", x"38a4d2e4df345d3c");
            when 5771230 => data <= (x"d6b1f7fff234059d", x"924830ee96ed78f1", x"c07711f7491580bd", x"7a36597f42867fa4", x"06a5e476aa03efeb", x"d0eee10af2684212", x"363483bf6855bb1d", x"eec7d2da1253c25f");
            when 31205568 => data <= (x"0c485445c880e1cd", x"8b117f054e5f1af9", x"c8b6f99a77dcf5fd", x"ecb3dab45bc7c650", x"bba93944df6f6fe6", x"f868376f6f70eb28", x"475426e687598137", x"9b890e554c5fd9eb");
            when 4462252 => data <= (x"83efac7b5bacccdb", x"b465d3ae418ecd60", x"84721d7730fcc9b1", x"ed7068030e00225a", x"bd5096ef0c416903", x"48d87549e7cc951b", x"d76c81179ad12b03", x"d4b6c328ed591d75");
            when 15693802 => data <= (x"e9ac49bee9c0b461", x"fa8bb9eb03659faa", x"596c71fd4496a757", x"6f426f617d4f86dd", x"608601466c422e03", x"2d1c04600d1817b7", x"92b3676367fe0012", x"769786419f90d4d5");
            when 6981884 => data <= (x"5c261a8a57bf4ef3", x"895fa03813b4aaee", x"deabccef1a699382", x"65cf2817a70ae346", x"77dd4cd1314b1280", x"e34c6e536464446e", x"fe839b569be11bc2", x"354862eb6f385882");
            when 22223949 => data <= (x"ebd5a16622c33686", x"616f0360573e027c", x"febcc3054bd6847c", x"1ad0e2588ef02d8c", x"8378eb1ac65b48bf", x"c2883055aa5f05e9", x"43511cea73f65f40", x"1c79176069907442");
            when 28510995 => data <= (x"f254b45f34fb52cb", x"811c8ad672b083ea", x"3f9271f4be4b9fcd", x"b58f7f914fadb0ce", x"404604a2f4d929f8", x"660d57dcfcfb33d4", x"57f13c503e27c60f", x"b3d6eca8e3620267");
            when 14296302 => data <= (x"5c584a987b6202e9", x"1dcc1a283a1928b3", x"ef3acca6519f3b88", x"aad68da1a45dcd0e", x"3a81125fbaca125f", x"5fefcfeacf739585", x"f0edcae6edbfc557", x"a988254c6f286604");
            when 10759183 => data <= (x"3dcd08cb957cb205", x"f1b823c9e7a309a9", x"e71dc5914ecf0000", x"5a481c619d344fa7", x"35ab118bf3104f4f", x"f4da1ee8677432e7", x"0631c8469dddcd34", x"c8bc2b1a0ae2f325");
            when 9475092 => data <= (x"a135ef50be023691", x"a30ba665945d66bb", x"03111f485a9349b0", x"7b412dfc8e7eee89", x"af490678644d2546", x"c39f7862afc9b63f", x"9d81271aef420c2f", x"7a6d88f0de323531");
            when 3680312 => data <= (x"73692a56bbb8d62c", x"0b70f39ce7121e1f", x"1f0d53ab130b6857", x"6109dbdd2e4737c4", x"dcd912beb3660cb9", x"d76ddfeba68c9615", x"46cef020d527176e", x"0023be45963d0494");
            when 6918807 => data <= (x"97c88b06d947598b", x"708f2c682f08418d", x"b016f7fad7eb5f83", x"e1c662101bc8d79b", x"d59e82674f1d7633", x"77bcb6ee090e4c4c", x"4e9a1e8ea7377709", x"2db9c418e28f7779");
            when 29810506 => data <= (x"a027a224368c06ff", x"7f787beb7f1a6162", x"9ffaeec032ad4756", x"356f1b799927c7d4", x"da87394fc6ca57d6", x"7f6646f5d2df7418", x"d6d94785d97e4a3d", x"4a71a300761daddb");
            when 17824575 => data <= (x"5959d21e96c451a7", x"d087096bdf93219e", x"d4341eba59d9f79d", x"dafe7134d181c263", x"0a6a94fbc7df3dc6", x"3acabffafa88c783", x"a44d803d369fdd04", x"3a6d44aa364cc7d9");
            when 25808473 => data <= (x"59e4443cbf5e8fc7", x"6abe5089feee3282", x"abc34cdb943cf400", x"d19ed226811c116d", x"43c1803a67957213", x"de1a55515f457159", x"3095340b7717f2c0", x"650ac848e96e82b2");
            when 21833286 => data <= (x"566a0555f16c6c87", x"125f5ac35477cac5", x"160b68fb54744a35", x"0bef1e0df22a18b6", x"4c0bca5fceb3ad6d", x"d4a54573eb348859", x"30479800f68fa674", x"ed3e68cb983be827");
            when 29251509 => data <= (x"d43d2879c5781712", x"1e1df57f9cc3cc86", x"7c5fa178da309d21", x"5a8c126db34860ab", x"a8118ffd1aa33d0b", x"9cc5dbb193a2d3ab", x"221238f035d9b4be", x"64777376afd0c931");
            when 2581977 => data <= (x"f69f147614b6bb04", x"e5088a69ff602339", x"23a950844ccef475", x"81b0f1ace11b9ca9", x"b04c5ebab6a39413", x"9cc4fcb9401d325b", x"0e3ef786b9ff1f4e", x"df4336bfa250c97b");
            when 6460330 => data <= (x"e8241f04779aa7fa", x"c8df51f07aa86229", x"aa105975bc228269", x"6108a3134fb824ab", x"3ab4ac3c16c4865a", x"e4977b81b017c67e", x"36f5bafa3c9f6c97", x"99c3b7eb1c5146c2");
            when 23230895 => data <= (x"3aa338880eb20d07", x"a34c197696641037", x"86342a001d52c0b0", x"3838f66a2a4a0580", x"3479de6492061790", x"483f444c244b6e82", x"181505a093c98c78", x"0a41b7be4aa6a397");
            when 24200891 => data <= (x"f249b230fc6aca79", x"d8b7b770eabdff06", x"d4a98a75f75bef7d", x"8f3e12271d8e6415", x"e41bc618dc961570", x"d65d93f0cdbeef28", x"ea940214c35994a6", x"4d85245a2978741f");
            when 31595131 => data <= (x"dd3266dd500edc43", x"77500f9ea7351dfd", x"82bc5d97ff4322de", x"a34e5b2c53d280ed", x"126f98513637694e", x"2b3653f968456aa2", x"c530c505cfc1c2b5", x"6b3c6ee3e402bddb");
            when 12185239 => data <= (x"700e8fd49d8c562e", x"04800feb1e7d0e69", x"532094e21636684e", x"d97e17ff019e7676", x"9e1bc3ef224bc46f", x"2d1ac031bbc6ecb2", x"ca30ab1d880c5001", x"0f720fd51a5a8bb5");
            when 32370661 => data <= (x"99888b2688fe3484", x"61b794314278ce5c", x"93647660ab5c128a", x"8c4da4d182728803", x"ab81dd9684a6eff5", x"dd1a20c7336a34b4", x"6b8b6f4e1185d2a3", x"af563a326de7ae3a");
            when 27057855 => data <= (x"2671b05ce2ccb5fe", x"6acc70a7a90dd0fc", x"d89df112991b78b8", x"e7efad67e16be238", x"a60d1db4442b6633", x"fbc444432f43deaf", x"865675db5da90460", x"17e449e019cbadf4");
            when 5235940 => data <= (x"c2d5fbe68f0d79c7", x"73a0810fb7cb9261", x"7337fec167b0579f", x"457694e97367fc2a", x"25587dfda850e1a7", x"6fb316b33a6ea142", x"d552b8ce7e78bd80", x"599dad9d7306e8b6");
            when 30655451 => data <= (x"0607aa6e6a3b10b9", x"6e63a0c8eafc4a4d", x"fe9bff39ecc9321b", x"f50a05823e229b49", x"212576038014795a", x"fed28dccb7efeb1a", x"3fe38735f0cf3b31", x"eaabb54bc322bb25");
            when 8282396 => data <= (x"c16ae44e19bbf464", x"9081ff5900318677", x"33cb34d01446011e", x"c8701eeaa69dec60", x"c8d5e229435aa1e6", x"296c5c9b1f51e778", x"2867677858da3132", x"f714249f8054c862");
            when 27425157 => data <= (x"65f323053b7844bf", x"08e5ac9e3fb03a9c", x"473c3dc4ab624281", x"e74877225c9e197a", x"056ed215ef7ee894", x"71492c7610febfd2", x"b67abaabdaaa2c52", x"d61fd82e4f98515e");
            when 19270497 => data <= (x"0752a2e11de85b2d", x"13e134b3a6a5d1f6", x"5aa54369fe1545f4", x"94a46bcd60238bda", x"f4f4fd930d05f477", x"ad3b109a014c92d3", x"ef34c47a0aa8570d", x"b12c099d330002b1");
            when 17290987 => data <= (x"cb64faf6facaf1a2", x"5ee7c6af98dc3233", x"0bd690a506d5c351", x"b018034befe434a5", x"b961ddc366fc4896", x"5a7ba7ec52d90a4b", x"ec0d8587a4fa9df5", x"a148a938dacc13cf");
            when 12126970 => data <= (x"98f9adc113ac938a", x"6bcac5e090838ba4", x"702e43e7d2794320", x"ec5f2c125bc77b3f", x"d16cebbdcca4ce91", x"3cc4cf2c90feabb2", x"52731979c565ada5", x"58b5b39ca64efd5c");
            when 3670157 => data <= (x"df4cc0ba911c7c30", x"ee7fd23c4abe2338", x"7297f1bbeae30047", x"100dd1deb492ed78", x"d6df9a1531b0697d", x"172463cb1a097269", x"70bc50679e6ef5c8", x"b4ddc8cfa9139137");
            when 31599804 => data <= (x"c8c084444d5d00f5", x"8b40b12111a54aa6", x"4e5022c67d3ddf7b", x"aaccd9424208222b", x"ca6b15b8a5d8a52f", x"963b162a413cfcdf", x"934e9322e283b925", x"c551f0bca465dc16");
            when 23666660 => data <= (x"4664cb7689f2b065", x"e5a914e2e7d4b918", x"f89a3d39bf4adc49", x"82f296f5b6ae248a", x"4317b7219f378540", x"7c124cb34e505260", x"9e82e7c23719e904", x"75624535b8afa853");
            when 10001248 => data <= (x"34fff3326c502415", x"36007eb2b77e787e", x"b81809a82c4b820f", x"8b4ed6b367e8f7de", x"cdeb5f9150498a6f", x"7c78bce22342c8d6", x"ac9c3fab5f336939", x"9e18f71298642d61");
            when 20437212 => data <= (x"4929c53a433370a5", x"59a3a2ff6824ce41", x"a9e0e287aee12cb5", x"cee8d4aab1bf8875", x"03a7c109f211c4ac", x"5f992b0cae731479", x"4f9f6918ae172cdd", x"78bcdc76e3e50197");
            when 9279365 => data <= (x"903c7ccf57363119", x"4740625eba95f79c", x"739d71f778dcc060", x"6583271fb168ccd6", x"c35436c126985dc6", x"ca343d12fd9e92c5", x"711a32c5740e2b4b", x"344c6fd1549dcdc1");
            when 7920649 => data <= (x"0b9cdcaac606d105", x"60a5bc8760866b3b", x"61b7bc686c72a065", x"43d747fb7aeb8281", x"6f1aad87e6a7899e", x"8a4ef83e0eeb070d", x"8da609de0b8893d3", x"5b8aceee9ac04910");
            when 10401068 => data <= (x"9be692d0294ad956", x"7cb7c4c3091de148", x"dfa5ff967d468a9e", x"85f7c4f9170cd2e2", x"eb404591105b341d", x"49bb8b4173739a06", x"8aac074ce0281326", x"cc4abdae046c8534");
            when 27881878 => data <= (x"55de16e60ffe094c", x"0bcb542b655ec3a2", x"884b868a9ec27449", x"70b146b57593813e", x"f02251359c88ac48", x"9afb023d3175b85b", x"0815897ad15a4cb6", x"339d54e124fb5a0c");
            when 17659757 => data <= (x"8f56f77116cbe6cc", x"64585943f0fe5d13", x"622ffad948e4a39a", x"d9a04fac11d3bd1f", x"1f7ca8935441d113", x"cdbeedc1a5b3701b", x"dd5eb59431a17d99", x"5461eae051e42130");
            when 21436689 => data <= (x"ab9a026357d7411d", x"e9f16e9cc6e8790a", x"486ed43f8d6bd72d", x"3111b428b0d62782", x"73956b4605fb4b33", x"54cc15033cc7f14a", x"7c145ee7d1487b50", x"013c4f789488177d");
            when 28285767 => data <= (x"4d46f8f2bbb223ad", x"382f90dfe955e301", x"94324eda03d59971", x"fe03cff361ccf831", x"da9b2f0efb6d6d4d", x"e7a85f3d2f4bb002", x"9a4a68dd1745ae8e", x"ed01a79ceabe2a36");
            when 9997419 => data <= (x"9bc731392d67c765", x"4f063dec289d6379", x"04f0a83031cdc700", x"fbcf4668edf5528d", x"cfb7d818bb6d5e71", x"72e67a492ce21200", x"09585eaf7de9dfb7", x"2696dc739a25e18d");
            when 31857649 => data <= (x"a9a5d608af37e5b7", x"60d9503e4874cf19", x"bb2263a6f55bc55d", x"aafd97dfd97de8cd", x"93ea9e054a809e65", x"7c36200daa75ffab", x"d15cc971dc12045d", x"9edb1a4a0c841191");
            when 12923554 => data <= (x"b29111d49cc7e8af", x"cb12c73aa7c478b5", x"11cb09beaf859b65", x"ec630b4313660405", x"4ee4064e773dbf48", x"b769257124f314ed", x"db545a8086a190b0", x"fc2644a459cabcf0");
            when 2386505 => data <= (x"fc305a2f11d0e230", x"1d7a4e319b676b19", x"a6e9ca4c4ab2e4ae", x"7974b816adbf093d", x"1912153111ca335c", x"953419174c356945", x"eef025f27719dfe2", x"720aae8ac766ceed");
            when 27388677 => data <= (x"f96687a476b8b477", x"bda38b9852c8a53a", x"31c7ae32975c8c4e", x"e703ef5e88752afe", x"d62d9120ddbb3ddd", x"3854edbd3dd9c9fe", x"fb14ea33362f823b", x"62b6b561d5dc8a06");
            when 20740549 => data <= (x"50001de02181afc3", x"c2df681cd97da604", x"361275a2142009fa", x"4cc40b0db2efced4", x"da1e8cc0bfb122aa", x"080d6d6aa159410c", x"fd8440d3e0c599cc", x"84793b36625db413");
            when 30043688 => data <= (x"cdfcd8948c9def71", x"791774ee159db2a2", x"34e21cb624b151aa", x"06dff91498fc4fd7", x"64d819746a012041", x"0859e0e822502dff", x"06e85a6040cc4b7e", x"31fba18702b75fa4");
            when 7346231 => data <= (x"d4f62f2748801889", x"dde5b130d3c416cf", x"07f646f7c3e7b888", x"bbe6f0486d050ed4", x"d4474b3ad0ff09c8", x"6efdc66410efba4e", x"3f60155be2450488", x"6c179dcc33dd87e8");
            when 3508148 => data <= (x"ef3783aab5a251f7", x"d30d812735c0e9ae", x"804d7d20dadf5d13", x"f26a1a08b7eb40dc", x"fd2b303b099f2450", x"8682a2d0e2e13601", x"7baa29fce296e4b4", x"73a2181a3a637420");
            when 25776793 => data <= (x"5e442a868778d1b2", x"4b3fd444f21ad83d", x"863a80aa90a786f2", x"3319ca4d799f59e9", x"3dd90d1b77e31ff2", x"2c768228c4248725", x"0698ad0529294b5b", x"cf4678b500630ddf");
            when 25243473 => data <= (x"d0f41f015675544a", x"bd538ec7b61fbf98", x"161c6932441008a5", x"1ed14065da31e8fc", x"7b2cf91aa7f8068a", x"274d4dde3f83d597", x"8e3fa156388f5e5f", x"3232c7089b3063c1");
            when 24103930 => data <= (x"fd6157ca285315fe", x"5e53a88fc80a00f1", x"558aaba99598bf35", x"9f7b83893946e18b", x"7e94881623dd6dee", x"b729ed7f47391104", x"2e6ee9d4d3defe54", x"45c36184b76316c9");
            when 24573591 => data <= (x"24f7a851b182ce77", x"4ef70612bfaf07db", x"e00fefce7353aeb0", x"b53a630e6b380859", x"94ee5fdedd2fc646", x"7d3ec6d2f049610e", x"086ebe28869f6570", x"08fb33d1a641c6eb");
            when 1411727 => data <= (x"12b68f53ded1e70c", x"3a4d2d80c36253bd", x"d14aabda378b3d03", x"a3037cc22c80964a", x"242cf39c87844c63", x"42d5cee6882065fb", x"e1e2de039ef38f94", x"4960d6c78eb3eecf");
            when 13495290 => data <= (x"e83bc45dca3e2a23", x"9a2c95e5a6a9df21", x"b62cbc4bca8986e4", x"5e70504b0fba6f6d", x"4d1e9fa9dec827fc", x"bd70c389c61e8f63", x"4af36b95bc81b565", x"9612cd55ca76da68");
            when 10068250 => data <= (x"53d921fe27b28272", x"9f38b68eb6b7007b", x"4e8969f4471e04f2", x"1934e31012f064fb", x"79f4c32fd508467a", x"cdb2b9e503d93fdb", x"a895e6ce14bc21d0", x"a928261863026a0c");
            when 18507156 => data <= (x"c8c7d2bba7863ed2", x"6990a95f504ca9f3", x"98030a67f7442b3d", x"6dfe4f916f176767", x"8966233823be7fe2", x"0903c0136439a031", x"a7a5210f1b60f808", x"3d5381c48cb1c1c8");
            when 9626514 => data <= (x"34e918d4fa7f79e1", x"aefc228e82f08d5c", x"543110dd83dbdd94", x"bd8b9daf31489d82", x"2d1730788ebfe642", x"193d7655d96b6c7c", x"b7938abdf47010f7", x"1292f734a5017f83");
            when 8412297 => data <= (x"bd3f6e61996f0745", x"349653f09584602e", x"edd40cc20d48d249", x"225006b9e9be29f5", x"6e9af5a49e189d5a", x"28626a6ef4b74a46", x"9bc3f53811d8a7e2", x"f053a8cc5278fa2e");
            when 13412671 => data <= (x"eb2c6449b926232c", x"34d1458ce1f74a05", x"7e9d84cb2a1bff51", x"f915389fb5d246ab", x"c95792992b43ff16", x"9bc4f965be5822e1", x"986b1659ccd663c4", x"5d43c9194c207b2c");
            when 24134937 => data <= (x"96122cbeaaeee83b", x"c27b262d3fa160f1", x"4b8c20fbaabb7a70", x"d5cd5206ecd2a5fe", x"0e06b0766613dfed", x"749b07fafb92fe13", x"57c88f74dfa4f7c7", x"49176cae5adf021c");
            when 7360604 => data <= (x"2edd6be7b12d9f3e", x"20a51263f3165ee2", x"a27bfd0c522b5f2b", x"1795a374097451fd", x"95101480f2e218ff", x"0962f2a8e8eb79a4", x"b112d3e81822283f", x"cf620ef44165372c");
            when 27930342 => data <= (x"8316434d16a3ca0b", x"453d71f37e526977", x"9f049d0f2d275768", x"b7301e0ecee8b8e2", x"ccbc8890f6d357c4", x"4585041e0becaa9e", x"3f70943b824a75f5", x"b03b7dbb53362f75");
            when 210146 => data <= (x"a98b77c29b0f10fb", x"9480a55ad82b1472", x"319d7a67c1223207", x"07923370ca8829c0", x"bbcd5a38938ab9f2", x"353999913ab71390", x"9ab20fd9dc2963d6", x"0f818c95f8de2cf5");
            when 2397593 => data <= (x"db0b4290dd56c099", x"6498d51fdd5f765c", x"8f9bfb952c8dc43c", x"47535f0e393eb63f", x"f91b52ef76f975cf", x"d3fa1cef7c32475a", x"8e05ddff0f7e67de", x"8165eebc868dbd16");
            when 21094975 => data <= (x"6e6560a0bb5e0df2", x"a48a79a35124deec", x"5d0e9eae3c674ba4", x"f61b8c9984edd63c", x"910ca2a08f9859f0", x"eafcd31c5a9a9acb", x"14f57eba8c428858", x"43268ecbd5e748ce");
            when 21651094 => data <= (x"6d2343a391e9b2e0", x"70f8bb55daf195dc", x"1d939a2245560568", x"5e246c38c195881b", x"d33680ca51bdb4ff", x"34ca187bbf1ff3cc", x"79b93ef4ad3b1def", x"de3204d38fbe8f64");
            when 15060198 => data <= (x"7de828fc42bbb4f1", x"83b5ebaf7b9b40c0", x"6251a9b588acb407", x"06f8a6a28341c808", x"ffe6d72895a698e5", x"522b38ca4d6a66c7", x"3edd2fa1ac23ec3a", x"3cf6cedc5b831195");
            when 9054730 => data <= (x"ebf0e2dc20560469", x"937459412189dd1f", x"6de708baabd52387", x"4bc9ea7f95a2511b", x"d4d8bff23d3ae989", x"e31de8e6bea9dba4", x"d41ccc3f7b74854a", x"e8abc48d694d33d5");
            when 17869343 => data <= (x"22445cfd00c87535", x"a18bb976f373c5c0", x"a772995dd7e446f9", x"d8b9404eb274b1c3", x"c9d9e72ab57d9ad8", x"438beea43ab61b80", x"39d1ec20485e0e74", x"29c860ac5ab17ad9");
            when 15071707 => data <= (x"63bc4cbb744c7db6", x"50284c24080e089c", x"0675758a01bea36f", x"6d395397f0f98c5c", x"e2d78b9716941acd", x"00122f07533d3cc0", x"a2ab18509cfa6c37", x"1707cc38f8529938");
            when 12309965 => data <= (x"cf5dbb45a1a24f90", x"8f4c7ac078ac99fd", x"098d9077ae5cc3f4", x"13a4e0ce2873d1f7", x"acbe184e0c44a60e", x"c24aa0216e2bfbf6", x"f90792e69759749f", x"342a0bffcd4850d1");
            when 8397381 => data <= (x"33d7e9d631010ba8", x"ac97f613fa95fbd3", x"479f1c8dffdfd02c", x"33a3174b00df1c98", x"b230cf344b7fa8af", x"afa5e8df4ed56628", x"bd749f6c759de8d9", x"d9b5cfa0c5f345bf");
            when 11737832 => data <= (x"3502faa3c086835c", x"e964dc92bf5460bf", x"e6e296b7546a997c", x"f685958cad66b490", x"2848fb9f2c239873", x"5866d34d8b7bea85", x"172db1741e498d6f", x"8fcaaa53d06b8736");
            when 32778933 => data <= (x"c4a5cbb0cd74b468", x"c900fe6bce9acce3", x"c553bf8d8702048e", x"35277d1195a574fe", x"235c781a68dc2224", x"88ae1a0dd7a49a77", x"e95e6e6c84351e58", x"0efcac4e6b4b1928");
            when 21479761 => data <= (x"936237889d2d50ab", x"bf8a26a7eaf3d6b3", x"e851182f3adfacbb", x"bcfb1bd125649e8d", x"a160061803fa1898", x"d1111d07deadec35", x"322c724378978c25", x"db4e5d752fc5b29a");
            when 32685682 => data <= (x"00b4de6fd7a8cf82", x"44001060315d5703", x"30de532a1c4c4014", x"44bd586ec72721a4", x"8e64fca8e4d8ea36", x"44340216a4f85ec4", x"6b9fc615d1b8f695", x"aaadeeaf3ef96278");
            when 31503972 => data <= (x"9cfda073ef152490", x"a5e1ed3c2e54dfb5", x"380f032faa94dea8", x"e4fd552ba097260c", x"87b6c58521bf7d97", x"bd8d96bb3bbf5238", x"f99807082841a47e", x"a9ec744546cebedc");
            when 11478822 => data <= (x"cb7698a28ee4734c", x"3b440b91f6d26034", x"b1ee6a5dc76c6720", x"ce115340ad064173", x"f082b88951b91108", x"694218d901a3538f", x"5ae69c1342764ceb", x"5790756fde0b8778");
            when 28314853 => data <= (x"4e35747d07d6357f", x"04ec784edaa1d363", x"f85ae18195e7be27", x"6d70df423b373b98", x"2839f8adfa15af41", x"9e9c15693b505e75", x"a9e3b7458eecdc87", x"fdac7fd986fb98b3");
            when 12354941 => data <= (x"39e97b4d907f7055", x"cb710df2bb2c2e16", x"d540253727c94ff4", x"7515fef5613204a2", x"a3087401ec6d8499", x"44933f4e39bbe369", x"3582c218531945c2", x"23b449e5fc3d17c0");
            when 26465242 => data <= (x"68b3346c2f89b0df", x"a17f95e7d134e803", x"3a3fbb2d0db290a1", x"3dcaa2ed36d2cff1", x"d363617f8ba873e4", x"6ff1f48e46cbec8e", x"b0e58e1dfc4284e1", x"395aa6fd97d48728");
            when 2760274 => data <= (x"4bae3e9a0ec12c40", x"dad44aad06840975", x"e4dfe3074b08aa40", x"9b772ee94fe8765d", x"a25fb58e4a759a65", x"489971eff77635cc", x"fc55d67d0d59885a", x"874b079622c2f8a1");
            when 3269120 => data <= (x"647cd981eaf84b46", x"ac590fd65872a01e", x"f4da7311cf91da02", x"60050521d73b7271", x"d2d9c871deb06201", x"1c4c5431752c86c8", x"602ff1124c15c0ce", x"2735a6d7992c1c3f");
            when 20643557 => data <= (x"28e0d85555fdddee", x"66cc02952e7d4949", x"6a39f11fc373a7db", x"713b6da4ccdef829", x"0b1591d48997d9bb", x"25dd98d5c7a54f36", x"17f630286edfb3e9", x"9eba963a8875e88f");
            when 8729106 => data <= (x"18b0a512f470c6d8", x"7017bbdbabc8dc3f", x"893e125a5a17761a", x"ad0b961658a4530c", x"cf15256e5d47a385", x"0feeba59ccb4ff54", x"6d737f8e55a43e74", x"4ea9bfe1a00c51ba");
            when 5682088 => data <= (x"9400d07be84a8c8c", x"c536cac5e974c3f6", x"a6b2abfe3910465f", x"77aae69b185cd394", x"5d17b59ec23e60fe", x"be07b37bb4e55c95", x"954ef5c96b898acf", x"2ad84a4aeefbad82");
            when 3254416 => data <= (x"ae203b948c3613cc", x"2bef06dbaea6f2ad", x"71ccd9944edbddb9", x"54793e3a861f76fe", x"d485f5fe62c6da0a", x"0a9bbb60dc56b71e", x"5621bfc4c7bfafdc", x"2ceed4edf545dd35");
            when 20428185 => data <= (x"cbd32bf0badcd4ec", x"80fcfb537cbaad19", x"e131c00d691a09d0", x"b9eca5e58f940e07", x"35b97fc8083d9c32", x"4742c7d252e9ad13", x"3c3575ead9a79856", x"254f1af5c73ebeb7");
            when 26799438 => data <= (x"ab90e0964cd5de98", x"1350872c35b062fd", x"05fddbe2c9058cff", x"7b8862e9119d7884", x"831cfb2be1c3a9f1", x"b67b5a3076b88b42", x"4f26398387200ce9", x"d81cf66a4964ad2a");
            when 813967 => data <= (x"32bdca0dcab8b436", x"230c088c8c883e0a", x"a2492f6d71a7486f", x"b2ce3ac51e26abf0", x"4beca158fe28819e", x"63b3bcec84acce27", x"5035e20297d564a9", x"24d093bc2a4df3ae");
            when 32236547 => data <= (x"10a40064bbf16634", x"e79c42238fc01531", x"40522a1577e1e90d", x"a18cff55fc202979", x"3e492c7d65210274", x"349124dc60d8d86d", x"57bdce30f6dc1caf", x"ccfc764c13e6de00");
            when 19703908 => data <= (x"c63afb72ff59eca4", x"084251b3ce8cb175", x"a1c3081a9d32c445", x"cebd6bb52e6f6ccf", x"b3f1e2555db571bd", x"9c9b7bb6ce5211ef", x"90f1db2d153a1dcc", x"00a1f555d738ecff");
            when 15536677 => data <= (x"99d648b045a64f84", x"648e35d3f0c08211", x"34e8f5dfd6f0fc2e", x"210628b46c31f470", x"b3db9e0e7e04216e", x"5816134761c9def3", x"6a134ce6afa4a6c3", x"8a89fa321ee70db4");
            when 30280656 => data <= (x"37911565df3c29a5", x"47c10f0603947517", x"b34e357bb7cb93db", x"9b55422aec750d1e", x"947c63645e1ab459", x"50d393b316e28e01", x"c050455c3dd40b3b", x"1f142a09dc610948");
            when 31523270 => data <= (x"ae7755d709acdba2", x"79f4448e23859a26", x"efeb61404d437e22", x"9a6e7546c3d49c12", x"c7b2c567bbe747cd", x"3485bfa7ba986004", x"f4e6097d1cec9149", x"64ba740bed15014a");
            when 33259786 => data <= (x"671cb59da2e26ba9", x"d4c2abbc5b87f1fd", x"8f7cd6aa4c6a14fa", x"bcb26ff400d46d83", x"4b4fe82da3b4121d", x"15f36d4aaba0937f", x"96873e9843856e01", x"73a7b258f904f735");
            when 24151068 => data <= (x"7d264cc983e6ece1", x"be91e695cf8b201a", x"b0bfca3cd99bf420", x"857b2549591af740", x"3e4da2f77a7c2ff8", x"4ca9ad6e07cb2626", x"dba4f8a0b752337c", x"cdf31ac31ffcf580");
            when 2767952 => data <= (x"c71ead2c90fb495b", x"c1d4ec3bd0d0bfe0", x"807be6602b950c5e", x"43c07d1fb116b875", x"2f455397fb2e42f5", x"5ad72b91a775db5f", x"89a174c1bad4bc99", x"fd280e8231fe47d6");
            when 12517291 => data <= (x"604b387d21d72e17", x"9081d34cce7367ac", x"3afed6a9b1d4e255", x"23b980d07e0efa78", x"e03af883c365326f", x"639ce07e636f8c3b", x"027c046b6f8cf0f3", x"b97e3947b4626ddc");
            when 31548312 => data <= (x"ba22b30f24e3ba27", x"def53b423219a387", x"02c773396cef86c3", x"ae9dda723231ff0b", x"9d3e29b4ab37c263", x"2dc4f0d6208cc1d0", x"a959d418e0f4bec6", x"e34567de523b2bb7");
            when 18114560 => data <= (x"29a70444c8884107", x"bc41dd56196c1b8e", x"9f88800be6352ab8", x"0de3ed56f5061f62", x"e66f3d76396bf7b0", x"f6fe17fcbb95f774", x"97635164e3e610e9", x"cec576196f55568d");
            when 947440 => data <= (x"4a2e3f6166b034f1", x"c0dfdce019f52896", x"86249c6b3772f608", x"b8b31ce62b7ab97b", x"ed322eeffa1e4566", x"0a0146cdd6425e8d", x"86491d36fd744e33", x"c40d65257f791a4e");
            when 15198191 => data <= (x"2cbaecadb183ec2e", x"dee4e27da35e7f95", x"8d2ef5138716afef", x"7fe2e1b479015e37", x"dd592d11a00d1ddd", x"da5de18eb328f849", x"15a08b00efd28534", x"7878138dc845f89e");
            when 26866127 => data <= (x"1bb0510251922323", x"7b6c690e389ad2a1", x"23b43a52e57f18bd", x"de5323a51f370e60", x"ced712b9aa025bab", x"3d3e39730bb482fd", x"c8b7c4437c0e6548", x"1123f52ecdd43b13");
            when 13068964 => data <= (x"6db1934594735777", x"e58e8560b3d638d9", x"da0d9a5c5c77c170", x"526fa947a1cf8322", x"90e5ca12da125624", x"f278444dd4c51c9d", x"f92073100e403ae8", x"62e1b78e041bf9b8");
            when 12803822 => data <= (x"808ec236f92af5c8", x"c247c2deac6e8b2e", x"49d08afc68e27330", x"9b45ff0f09b78f51", x"373d531bd5b4579d", x"72f0a4229735faf1", x"33db869aa8d7de59", x"9ef0147927a4882a");
            when 8188626 => data <= (x"b75e1fec101eff07", x"0d409ced8589f656", x"033717d380f28d62", x"efd244269f2ea07b", x"954641695383fe03", x"3fe12fa28ad36004", x"22b77a256771dc1e", x"b4b268695ada7961");
            when 17511513 => data <= (x"72cb2525ae967a1f", x"231301aa6688129a", x"d3250b3aa6c10aa0", x"7c07928140cf8a9b", x"478737aa79f2c76b", x"6bd3203a88d32805", x"553b68a1ac0f6733", x"5f0168b08011f7cf");
            when 24712531 => data <= (x"ddc92be1780ea528", x"583420bcf477c012", x"0f46148bfbfc274c", x"487be2303531e505", x"150363a8196bcf70", x"c06639af47438682", x"f39a5ad5e72916ea", x"26c3b4574985567a");
            when 1819980 => data <= (x"4b53c10a48a1f71d", x"f3896eab4897e26e", x"958109f9ffcbee8f", x"9129e6e6e25a0460", x"f68a6a046583ac9c", x"8872ee3f324eeba0", x"2c8fe8fd272ea34b", x"fe1fbee63bdd0e32");
            when 14898745 => data <= (x"1d6bc1caa86a3f81", x"732f0c9ac8959357", x"491ab9fd39d53766", x"e52fb8f1741607f1", x"a0d3f3e0de8c8468", x"a4fb050ffa6cbd49", x"d591643b1168a049", x"0baedd622c53d4d7");
            when 29888298 => data <= (x"52d801a1792ac7ab", x"036b0be5584b3919", x"e82ad90320e70ebb", x"47dce8c06e76b934", x"3de43640e0f1d8da", x"044c887533d64916", x"ba54528ac4da2474", x"4817dffc6f13a8eb");
            when 26671166 => data <= (x"999b482bd80d90d5", x"a91610545a8cf94c", x"43376e3107954819", x"0a9d74883637b44d", x"6e863c01225d7fa5", x"58730ddaf5619ab0", x"7ad8151872be375f", x"e123395efdec54bb");
            when 25352307 => data <= (x"d631b24e0f40fc82", x"caccc744f55c98af", x"09858ca884af3b75", x"ec276878f7375f48", x"daad9da05f723e29", x"99788d478806de7e", x"d2072ad169a4bdf6", x"8a8f660584bb14b0");
            when 21189590 => data <= (x"3910178b39fffba6", x"31e8ff5cc41313e6", x"9e474594a91f7dbd", x"7ef1b2bcb670ba03", x"1304ab8488f761c4", x"325a6660dbfb331f", x"ad2288ff9045302a", x"1d064a4e86128df4");
            when 16320817 => data <= (x"8d30ac7c67295cb0", x"50ff6f464fe2d61b", x"9c198cf42287a533", x"e2850100812e9f61", x"7c393f3252e18e04", x"06993cdaaaafd3b7", x"d0b3c3268979a036", x"b3ceb9c2d90fe1b0");
            when 26033708 => data <= (x"fa7de07cb879f9a3", x"e717636c22246e14", x"7b740adcd2fe22e4", x"db17b4e9ebbeefec", x"632595ad1b2167a8", x"33ccc336a87c3b61", x"4350467aa108c0ee", x"75e1309e4164e8b8");
            when 11017737 => data <= (x"ec7f320396d48fd1", x"9fa27251c859b37c", x"a1591f85361d3796", x"d9a54dc1da6c077b", x"77f411da6a923bea", x"3a38b5df1d06c118", x"e7084e4d2f7f69d2", x"9cd4a70d7193666e");
            when 26175416 => data <= (x"2b5611f625bba8f5", x"e14cd499cbd7aa8c", x"09bec20e27bc1eb6", x"cd9dd81ce2818825", x"e5e55eb2e9d6e2dc", x"eb49c673a7d8fabe", x"4ac16b3c6de16e1d", x"b8f87b1c707575b5");
            when 15912303 => data <= (x"e2766c8b6fc5b759", x"a3601d8c0e6bca3c", x"c4b426c59473b3b0", x"5233316647325166", x"36e1b8da2af68fb6", x"277a9880f467bd8c", x"7e16871a6c9399d7", x"07469d8e796915aa");
            when 17537513 => data <= (x"853900e14b5c67c6", x"5f94e656025adff3", x"39a0fb0ff4385a0c", x"d21fa86a601e8546", x"37067236e7b6faa5", x"afcf2bc89d6ef1a0", x"5f3cfec54c502f57", x"3627c91c87087ed5");
            when 29968089 => data <= (x"b1ba06c537b99a08", x"e5e71e7275e224e6", x"b1f15b8c19938688", x"55198030bc2652df", x"cc11c97c17a3492b", x"c7752872fa64ce14", x"ed20e6d6a042e1db", x"75d503fde78a20a0");
            when 10391035 => data <= (x"ad973d91b08ff261", x"891a7cd3f59d989f", x"b5bc3928081b77de", x"9516f08395aaf8bd", x"a0e9a954ecffc6b8", x"466db354ea92b70c", x"2a4548bd58d77be7", x"face273092b7308a");
            when 29542294 => data <= (x"84f231f3a0bf50a7", x"154465ea8c73e6d8", x"f3054116a468a20c", x"bba13cd8c2218b57", x"77be33653a882770", x"974cd5523d5deffe", x"d5de94a9d45c3514", x"e5812115f7bfac86");
            when 18495470 => data <= (x"a0b3d7e9d6c0392a", x"f59599d10f18460f", x"fe3fefcc13d26776", x"384ea8da7c63cab8", x"7d4a6c5c15cf13b4", x"e7a41a9d58a65a41", x"c32fd34e87bacad2", x"d10223df50d714b4");
            when 3945852 => data <= (x"f627ecc2dcd21e06", x"f59175fe9f41f555", x"bd775e0b75484c9f", x"e7b745e9dc017269", x"a51804d9a772aa07", x"455c0cc8e6f515db", x"08b13c47d675a070", x"76a2126782303cb4");
            when 24276181 => data <= (x"bacdbddef0583913", x"a43474ede95e4e6c", x"9d9d2716e1b398da", x"d09bf05697c8b455", x"681c42518674ba6f", x"3f92badbcd34cb42", x"39e939d269bc3e80", x"7be52b30f1065e55");
            when 31891835 => data <= (x"45e1ff85a4e1be0c", x"7f8341063d833e4c", x"ee04b84e7f39287d", x"76020cfec1d003ad", x"27ccb88eccd4c23a", x"ed2b631b971b9018", x"933c14ebb63ad24d", x"930f218ac216ed2c");
            when 27153947 => data <= (x"3bf4a15e61e0da6f", x"607246c942190d4a", x"309d1c9055b8adc1", x"602803634f99ecce", x"daffba38b9d5805c", x"67ead2366018b4af", x"28a47a399f7b9e5c", x"02759bf7b0837b81");
            when 8032974 => data <= (x"e96b81ed1c558950", x"fc61112330f03516", x"9bf71bd80050d611", x"76bd70afea43d79b", x"20f70c86796117dd", x"f93063fe3769c7a5", x"43dcd9799e799608", x"7d93034559d5be5a");
            when 17971432 => data <= (x"634729d83f526ee0", x"8ea0d43f62e148dc", x"2982de6c727cf820", x"16e544d92e3997f6", x"29a0ef470e06dede", x"c2774dd4794d5b03", x"b86d48c8a76ff5bd", x"f9b4468a5472dc89");
            when 20460655 => data <= (x"84fb44ac813f4eee", x"2cb776eaff6dad84", x"06bed75f10b5c70b", x"f916abb749e64564", x"a9654df93fa5bad5", x"54b48799a620cde6", x"72d59be6d884adab", x"7cca31badd6e7ae0");
            when 16277774 => data <= (x"c53ff9591be82ff5", x"8cd9171dc765a7e9", x"95c966c17cf26185", x"b97229d6525c0743", x"10268ca6d58bad84", x"de4289a4f9a274b1", x"b84941cc45ea559e", x"22e06cf0605c33e6");
            when 22963652 => data <= (x"a406d04502aea804", x"3d4a566faabf4825", x"fd44b9976f8d03ac", x"943347f16b049ab7", x"77b4c546b3030cc9", x"e669c2eebae83891", x"39f6d1edfce64ea9", x"7d87d0bd5a0227ca");
            when 18218880 => data <= (x"2ae036bbc9998d68", x"78f88da1e18351c3", x"aa1e0da2d427e3de", x"c1e88a6071cf35b7", x"c67bfebaaa572ae1", x"caf0e02c8a01b25d", x"581e588ee37b3765", x"a1d4ce1cd1b29eac");
            when 26941260 => data <= (x"5de4692e8246d346", x"f8f702bd69ee3e18", x"a909e04647354c4f", x"f5c5e9672817d3c4", x"708129a64bdd7880", x"81b2cd0af5252904", x"4fb1a455e1253db8", x"7887aaea161bb798");
            when 21483802 => data <= (x"2e0c4b4ea1945f2f", x"3c11e023e7d8f176", x"b4d26f0992adc363", x"b7d30783237ae1ca", x"92075fe6c9b62f45", x"792d1a3b20aa4e64", x"2c0f07c01eeb741c", x"e8dec56085848951");
            when 26069528 => data <= (x"bea9af8847dd1659", x"50561e65c0f22a21", x"2217391414856af2", x"93079bf0e641e5e1", x"4759f78a62b5fca5", x"274be35fa0821d23", x"78251f4d001a8f55", x"8448a36b02e43819");
            when 16882013 => data <= (x"84eccfed374adc43", x"684268f2979498b0", x"062ae9040cf23f4e", x"a695be6ff9643900", x"57e0941e6a6b2476", x"669b94e033b354cc", x"a3d9e25e2fe0db1f", x"c751a7f29ae64b1a");
            when 12150571 => data <= (x"78445de42e9ba5e9", x"922e85943c86c360", x"5ead1200329c212e", x"652e1bd539b5191a", x"dbf7d39a42e58dce", x"b321861623dacda8", x"63ca53385c2cc861", x"bccf16e942823d1a");
            when 15928448 => data <= (x"427cc85044b5dc38", x"2eb5f96483ff846c", x"51975e737f91b8a8", x"06071b60c064c1b4", x"4e7967f9b6d1935d", x"8032c7b7088e55e2", x"207fe302f3686880", x"8dfbb708ba06d461");
            when 3993324 => data <= (x"b74f83a9bd8bd742", x"6d192d079994a5de", x"2b5cebc5cc1377ac", x"606fd12f6d3663e4", x"796a3eb5dfe821d7", x"087abfc0419c3a25", x"f17f1b081f3820f2", x"abc0e413682c2b08");
            when 11628609 => data <= (x"0dfcc3165925a5b6", x"1401d336c2c2bb9e", x"8cfe01597a2ef5a2", x"9aa4b14f6015813d", x"72cd77991ce41b2a", x"64620e01c287d32f", x"01dce363db34be0f", x"1ea8d32a39b2849b");
            when 2570372 => data <= (x"1a2a5da1907eb785", x"2e088a35c297ae6f", x"d263e8b673535264", x"f736002db67fa877", x"deaf1df9e9258ce8", x"9701bccd86c3f5ea", x"520b4c81a0b8c6ff", x"fb175800610dc8bb");
            when 11089200 => data <= (x"7b4bcc5723c1484e", x"2a70cb9a0cbe1b2b", x"a00005cdab8384f5", x"2dcf95847efebf36", x"29e7a02cba8aa550", x"8e7ccf3e8a719a34", x"e1d1bdfdb72982a1", x"205489a41d4358e3");
            when 20747297 => data <= (x"475fc8a1b48cb7e2", x"5e21d7ee887c8ff8", x"a9a08bc634e45587", x"97e6421fe3e90773", x"ca25fc3d7e163617", x"d973d93b57c91bc9", x"cff08190ada764c8", x"6ede24758c8610a0");
            when 14155428 => data <= (x"7de5f90b65e2a1de", x"869dcc0e94f78eb9", x"e78451652db89707", x"993db0d3c75353c0", x"b4eb0491e91a2e99", x"a02ccefde110d052", x"c951248a314e7114", x"42d00e49e0bc6f63");
            when 7318856 => data <= (x"42480e09292cd596", x"5a86be2e7cd15562", x"6cf0b426f2346af6", x"27656f5ded19bac0", x"8f30dc6a08961e6c", x"5a8b5e99d441d791", x"167f59df136f962f", x"c440bc1b4e9c38ba");
            when 4092604 => data <= (x"d8ebddde2167f1af", x"d06487ca01b3fdf8", x"d8bcf626b29a6bee", x"adb6929c0bfdf1a4", x"5257ca943344a958", x"5fd011a5958b2ecf", x"7b410660f86f6a1d", x"50c2819f864693ed");
            when 27019383 => data <= (x"1f5dc492e0655c51", x"498c2205022b0c05", x"fb72edeeb29c5037", x"6a22ca28f190407e", x"e6119b8dd3f48883", x"5bd13317ab1698de", x"8bff24f6468b0d80", x"4df72b1e0bbcc99f");
            when 556028 => data <= (x"f13c115563172c14", x"c5ff937f6ea5c14a", x"efc8948887912c3f", x"e174b61c67967a15", x"1013435df12cd535", x"eac7288352820111", x"cf521c45a9523cc5", x"043baf107a7ec61b");
            when 24547304 => data <= (x"d85434451924392b", x"0654e87f1f53c378", x"d928a195c438f75b", x"6d26b8b5b29d416b", x"0c98c317122dba29", x"e0459118c38aa721", x"03fda901afc5a135", x"79724254929b8b64");
            when 6004111 => data <= (x"eded612f981d6dde", x"faee13f087899770", x"6a022c6f7d1fbab6", x"4dfdb6e3879f33c0", x"c2c6a05ffe7636c1", x"efbc08b42c9fda07", x"46e796f139009414", x"82d3ab6e414e780c");
            when 18259598 => data <= (x"972ca8d737f21979", x"f72c07eb70a54f09", x"dd58e497eb53307b", x"b9c4111983f85291", x"f9a1054d912d19c4", x"d8bd65ae5ae6c4ce", x"839a0d665369cc4a", x"7782a6a7839dbe36");
            when 5250465 => data <= (x"dca0e01a8295264c", x"0ad521b1846dab40", x"ad9e29864bbdb51d", x"98d59e0095846c42", x"4d4e7c1f1bd3195c", x"7a7b13fc4e2462d7", x"96af4aa0dc5c40fb", x"5798dd0470d63aec");
            when 21275037 => data <= (x"a104b2e271f3e755", x"dad47e8aa32d4ef3", x"bf173ae4afdfa3e5", x"cac5f977053b8567", x"a4f280644861df3f", x"f8b5a7f068affd7d", x"4b047a3e81f26f93", x"559f90fb2181ad36");
            when 28521923 => data <= (x"f847b5938fe26e9d", x"24a1e905d38fa666", x"658f0d9c4cc496bd", x"54cc7445c8210d8b", x"e65f63735c17691d", x"d495552968398711", x"e86c8c64a1f42f00", x"3eefbdf2f1c3a6a9");
            when 3975092 => data <= (x"fdd8f1809c36f109", x"b440f2557437b191", x"8f509df62ec99f90", x"973a0e625483323f", x"3fdaa0b73c4367bf", x"089d60ab8fda0d73", x"10cf4fcaacc18338", x"224183a5db22ca8c");
            when 19620267 => data <= (x"e2822d88bea98c6c", x"0e580d8ff8a53f3f", x"4b0c18aa073ff3f5", x"20f8b159bdc6c07c", x"dae51c002710c25b", x"23e3cdfdc3e22a02", x"3eff3b5f51c4288a", x"f6fe04920b1b576c");
            when 26658421 => data <= (x"657fab9eb955e949", x"b12c6557f5b78cc7", x"3374c45fc3c56e6f", x"5d3022e9a45400bb", x"42df63167e5c2333", x"4c9d7e1f9f54ffbb", x"da19cc9c5a860c71", x"777a0f90f3203e17");
            when 12918273 => data <= (x"f7c88bdbff765e8f", x"411b29a217140136", x"483f91a4355a7779", x"6dffd16d88b7872b", x"1ed555e9d328d8e1", x"43f157d67358e3fb", x"23d8f04612c0cfb5", x"901edfe272947bdf");
            when 17953647 => data <= (x"8dbe5a758a12c2aa", x"e4a7714f1544c5f0", x"862a9b80d2a4ac4e", x"2743b88d7c370c5c", x"d7fcd5e1b76be7c6", x"b88b016751160667", x"d28ae45ecdb2dee6", x"0b98af4ce58c499a");
            when 4298637 => data <= (x"6135bf793f850be8", x"33b9be71765d2c28", x"90260681cd604311", x"29a468b776210e14", x"7bfe4bd348f36f36", x"4a759264ba4cc85d", x"afac5f86539cac72", x"3d29e2b5ffcccb45");
            when 2455929 => data <= (x"5da1ae592f32e0ac", x"0e4f9f794c0dd4e2", x"01d6fe712532b055", x"e8f513a64ab6d822", x"08fb7147e81ef92c", x"e16dbee8621cd45d", x"d0e1095888816d3f", x"0782033e1e053912");
            when 15159420 => data <= (x"1b07f60a4138b064", x"da6b586fbb32b6c6", x"94e61d2dc20a384b", x"bcfeb43e2fdf3955", x"6f5a5912c32854a1", x"987a62c74b2651aa", x"7f36462e7ce17525", x"9a0b09f2bbd58d74");
            when 7126143 => data <= (x"a0297a7c2525848b", x"6d5a45cd299b047b", x"46c5003415c56471", x"52715f54fddf9b33", x"3a8c1030d8f198d3", x"46d2a7e4c42d2a15", x"ebe2b51fb48329f9", x"908995decad48f84");
            when 11136229 => data <= (x"fdac9a24cc2c3b9a", x"766d358eaed723cc", x"d9743e45a0e4d9c3", x"9335676fac2fb016", x"131f8f415eb51f6e", x"aa3aa3fe887fd7fa", x"adb86d41d5ee39cd", x"699a4cc37ae07a09");
            when 10334087 => data <= (x"baadd45654bb46f9", x"caabe5e1be7fe56f", x"b785a7454826ea9a", x"a05351edb3014d9a", x"1ba03b96b4f0e710", x"4a5a55c9dfbef7cc", x"d1518e500c1f168f", x"7348862008f3b651");
            when 3058364 => data <= (x"2dba8e5be85fdd97", x"a7cb20a17a7f808d", x"d7427d5434f85286", x"8b0c15810ea88da1", x"7789f90530b76ad1", x"65ef2a8c7e270fde", x"1693515f4730cdcd", x"ceea8b4f9b23e8f0");
            when 23876264 => data <= (x"33de5f7a72e74a79", x"eb67d8bfbb7b90f6", x"fec0186c6902b083", x"38c4920da3c6014f", x"7742feb3ccb9bd9a", x"c3b91a126623eb70", x"6cf5e78d3acd3bc0", x"5ef48c6c6eb874d5");
            when 27816632 => data <= (x"69dfff3fe1e8dfb9", x"6745a7a17fc69573", x"65e78a345f163690", x"db51ca4d6083477b", x"6465caef0055143c", x"28d0109f790427f9", x"3a4ee35e8c5132d9", x"17cec3e39faa7a04");
            when 3163212 => data <= (x"cd484f1e8dda43ef", x"d2742c77ebe44b84", x"f413ac8a91c09541", x"3dca802b44890d66", x"6351978736d36761", x"7bb8dacbeaf9eb22", x"b2002563aa61792d", x"eab80163b2c8ece6");
            when 20554940 => data <= (x"4550a15752d6a01c", x"0950827e2952b0c1", x"7af0e765066a939d", x"4800240e58141e1f", x"660e44b2bdcdb6ea", x"f875b12d8a4c3399", x"e2cc584eec3a9d84", x"c2d9cbd679377fe4");
            when 23729132 => data <= (x"aad7dfda93da8ab9", x"87dbd762a17b0ce6", x"8e4ee0fb98593559", x"0b437cadb63c2f19", x"f53c0a78598ac0df", x"403c89c0b6449403", x"d41393b8cfaf86d0", x"7921c4190bd67d6b");
            when 25963842 => data <= (x"fea2cc83da417e86", x"418a11fbc60f1890", x"b5f11c1ee4f11114", x"b51a8561ea12999d", x"9cdabe90dc529e84", x"6c9c0b9d22ed142a", x"a7e4925d4ba64b74", x"942f8133e0567f61");
            when 20481282 => data <= (x"f76e84d6ef84d26d", x"eee8ca84346f3ae0", x"a89487a0ce26de07", x"95d1edc6cb4334eb", x"aa7aa463927c6d42", x"65dcdb8c3747e33f", x"1db586f75b5e9da5", x"f0a6dd017a17f75c");
            when 30631237 => data <= (x"060636f0ca2527ba", x"b6f933e71a42771f", x"2182a5ed1d7b4f1a", x"2fc938b769d1f7f7", x"c5890197369c91a3", x"c2a6e9ef19c9b044", x"d03bc64531cc7ddb", x"25fb3865e969fbfb");
            when 11645752 => data <= (x"709b8dbbbf45ef9b", x"d52d4c8314f36087", x"09c3252eb587fba4", x"139b448c5e777d30", x"775e58c1185a61cd", x"778dc6013de6b214", x"97ac42c3e02f1431", x"6e41aa1e5543aead");
            when 26600810 => data <= (x"73e4c969b93f1a5e", x"028242abbd27b8f4", x"fe0fd76fc3e7d98f", x"8662dde33addf295", x"a1b15d04556358fb", x"d22b73d6193dec02", x"3db9882d2a10ef98", x"bb24525a4bf6914f");
            when 15175342 => data <= (x"1af78156378df35a", x"3ccb73c52dc36044", x"e26650e9c510fcc9", x"d6b8d4f3af823261", x"60f110f98657f8f1", x"8b7adbaab8a8fb40", x"b3e03bfd21446d3b", x"15272570f51e40f7");
            when 23717401 => data <= (x"16c8cda1f65d67de", x"321ac9fc8b541186", x"86648e188f59f8e6", x"083241f1183bb4b7", x"5e4472cac91ee3c8", x"8a4cdcc0ef3f4fbb", x"75a3437c346dfd8f", x"88ad200a449353ac");
            when 5872950 => data <= (x"c5a7db2ea2b13536", x"9dc7b6a3ce6cc758", x"ce0f449a0bca6757", x"3ea8db37b0a746c1", x"89a3ca99abfc31ed", x"19198aa61b9327a1", x"4525c868ddd4120a", x"348bf068efb06515");
            when 27101750 => data <= (x"5a7d26caaecba659", x"1a35cdf35ec7482f", x"652c042f4dc7f742", x"0f520c8537c81fb5", x"c7a81251c9a8f411", x"492d0eb0223b3595", x"0c3750cce4c2b72c", x"519afe84cc6dad1b");
            when 27500064 => data <= (x"3a33505a56f5059c", x"cc9bd2a238e2089d", x"6cf3f78e33483324", x"6b95db1b424874a0", x"c117071c862445ef", x"8560ed073a39e8a0", x"44395b8d434df427", x"1fd24dc4e9f937be");
            when 25506970 => data <= (x"a53a2c717bf1cc97", x"501c3dc92819de87", x"d63b7488a3e3d0be", x"deac3cda8d31d20f", x"32ad07c6603424a7", x"09907902442caa6e", x"929828c7cb6cdb89", x"cb4ce7aa236a729a");
            when 20652045 => data <= (x"265e536e90533d0c", x"d477607653ee9ebe", x"52acaa57e36945b6", x"2c28d8aeb2939f67", x"d0f3ded366fa46fb", x"c565955c848f88ae", x"b04f9723cfa5158c", x"d1f627ec410983ba");
            when 21943280 => data <= (x"5ed6fc6b9435d3e0", x"6b2d82132646ae0d", x"a585531f887dd7a8", x"88af6203fb1574ba", x"9347b6534f2e7900", x"208572518f825134", x"eff0efe8c32b13d4", x"c8aaeb02cb45fe76");
            when 9879864 => data <= (x"6a6fb73991231c0c", x"89fa7f8ec2fedc2b", x"bbd85ba79d132b20", x"3c08d77cd1aef92b", x"809ce86d548c866e", x"137781427fb6d3e7", x"4509233170f9a6ef", x"8e5ebc679c28820d");
            when 1084655 => data <= (x"7544475a7520d214", x"4708098cac1ead74", x"2dd1dfdf3110e32e", x"2915bd5b7530d498", x"b36bce51de5e7843", x"def05c0537db3b3f", x"643d1823e0b1dd9d", x"683afb8c791e3b8f");
            when 28607104 => data <= (x"619400ac7c255f43", x"9f8b88eba1a42360", x"87472dec3fb91f11", x"10ba2b300be11eca", x"179e6432b43d09ba", x"217f34de164e6234", x"953183a542856787", x"22e90be0f3903d37");
            when 11867839 => data <= (x"87b4580832b7ee47", x"3239ac737cb39e59", x"9cd8dfa33ba80c10", x"1381085574689aac", x"2ca9705f48f12b79", x"bf0fa075b395662b", x"57f966a8c88bcea8", x"7b567eb9089e3231");
            when 27971183 => data <= (x"9c6380de5a6577fe", x"38454dcdd3d71892", x"098d11e8545bf072", x"de7803901c803879", x"90fa86f44421567c", x"b696fa320aa47047", x"e2c64593df7e5e87", x"ea960198a3bef2f7");
            when 25947580 => data <= (x"827474b74b22f07f", x"076b806fd50729fd", x"7a246db0d6790dd2", x"fdbab9b94f042319", x"15da5a2dd3cf57b3", x"b8b24d2eaf3951d8", x"7f6b225f28dda5b7", x"2624f2cfb6b9ef80");
            when 31068615 => data <= (x"93b36e76b21317ef", x"c70387cd9bf3eca1", x"0ee26737612e821d", x"0c562428a4d2a55a", x"df1815c162a83cff", x"eae10bb35e2c3600", x"81d0a85da464a7ae", x"7c66bee5ae699270");
            when 11909367 => data <= (x"2a938105b8414ce0", x"0b0c1c29753208e1", x"7ff43d2489b4d7ef", x"2a292622c5c83ccd", x"fe84ab7fd05d838f", x"ff98f9d4cb8aa441", x"6a15fb36bb1ce00f", x"c1ce5618a65f4e80");
            when 31809534 => data <= (x"fb24a2d4863c6a1e", x"1f2f1df85d43f1a1", x"cf4a21f3d995cefc", x"a60f7297e72e9b3f", x"af096db0705627b7", x"3ecc9dea5c89849a", x"0829fe9d1687d35c", x"a611c0935b8d0b6f");
            when 33071422 => data <= (x"26b48e84e322f0c0", x"b6e4ef0a90c2b45f", x"451ac1033ddc709d", x"8230bacd272d2a8f", x"b96c59e35a2f9df7", x"886efa363d610fb1", x"58a29c63046b9900", x"eb1f40f10d51a918");
            when 22332479 => data <= (x"dd5d0b33e19f9a1a", x"568d7ddf5720d5b2", x"de789fca68d32d6c", x"4fea27487ddf3a3a", x"a66f291597efbbe5", x"a4b58fa7bf5e603b", x"102d0506f68d809b", x"c53cc525903855e2");
            when 19855509 => data <= (x"d7caaf89c5a97708", x"c1988e862049cb01", x"b91f85182eaba4e3", x"0d4b50165a582907", x"b370cff7e04fa7f6", x"4ac3d2486ea602eb", x"18bd8ac1ef15a4f2", x"618bd15f859f4911");
            when 23639524 => data <= (x"ead855592e0e2176", x"4ea4b489a6bd3759", x"b3fa1d12938b974d", x"2c95d9c008354804", x"e11905992df7861a", x"645c5fc9fa10e5a7", x"3f13e8d53ac7136a", x"ba38f3ac1eaff2cc");
            when 11200351 => data <= (x"f6f7e04adf2cd5d4", x"36efe58f3d2e9006", x"673caf267501de58", x"c70a55c06fea06ce", x"1aa0006f9a819dbf", x"d4e82e4d067c4f34", x"7ccede67062b8644", x"cf4a82200fd38cd8");
            when 19046451 => data <= (x"764875784f531809", x"c14bec737228a16f", x"b78bb9ed2f692b2b", x"91a03e88722da76f", x"e7f6e5bb76c923dc", x"387f928f29134043", x"81a9688c78900001", x"535a1c75cc5e1b64");
            when 5299849 => data <= (x"650cd8872c27f344", x"70fe050e8dd61082", x"3f8126b4785bfd35", x"7770af2508e9776b", x"a8efd1b457e4af25", x"6afcd661c5261e82", x"1d75870941dc4496", x"dd4298357616a703");
            when 33843498 => data <= (x"5ab34db4a8631591", x"b12d4f2890fbfebe", x"3740b2f398f18a55", x"4d8b8379eaddded5", x"e37df60018b2ca5f", x"9850eb69c230e75a", x"16b419b474d9cee7", x"ba7a1c9aa1497170");
            when 465979 => data <= (x"37962980ff8f14d6", x"c665c1ca948457fb", x"f14650bec1236228", x"a78ce5967a8e8e79", x"98be7165cb1dfe55", x"6f9869e65e7b1038", x"7f69297f3f871ad2", x"5164359c620d95f0");
            when 15812026 => data <= (x"d026b30c8ba479d3", x"8a809b2b62e293c7", x"0f3ac9c53fbb6ff9", x"7a61b9852c7435d5", x"f8bee2e544a36e3e", x"60ad9cb67b1d4cd2", x"fbeb2d5b6c9e8f98", x"0d5ce7363bbeba9e");
            when 20876626 => data <= (x"09f8bb8fa72defbe", x"3e38ad3b5b4e52f8", x"4f71d7ef65002289", x"918420bf700062c4", x"3475a03211abef28", x"cb744917a3d1a26c", x"b2c19eaebe4c79f3", x"62d420fb38fea013");
            when 25306771 => data <= (x"a054f57e0938d639", x"ef887d7406e83617", x"c617bcb49fbd0b86", x"1b06eda0a379a3af", x"105551caa1d52361", x"21a1fd88ca2f72a8", x"d4752cbbd9b85dcf", x"382233e225d1c4fb");
            when 29492089 => data <= (x"ce578b9f764d8ce0", x"9383aafd74aef033", x"b8ef5512202f4bae", x"0de4dd52f6fc490a", x"e2edc831db200435", x"fa842a1af174685c", x"e0d4d96e809f8d5e", x"97ebd9f39cc977c3");
            when 17771923 => data <= (x"5d1aa375d87d08bc", x"f79387ad976c8e29", x"0b234116e91ad998", x"8988bc233adab917", x"58dd0db8d874587d", x"f4c6e2a72f38aba1", x"7a368992b5aec69b", x"9046071d46ac7bb6");
            when 28693865 => data <= (x"4ec8e658b8641370", x"ace4ad9de666e33f", x"9fe0c3ddb19ec066", x"7d7c5290d9c9a3e7", x"77c0f5c89847e906", x"77144d91db287b39", x"fb342cc130ce56b8", x"e1dc5c194b684329");
            when 4011408 => data <= (x"3117967fae595f03", x"3954e7ef7f43eb90", x"2966ff3bb9a6c1e0", x"2d1a99d814a37149", x"f7865d13d6508dcc", x"84b94cd5ce28e81e", x"fa56a981a446de8f", x"a6ef118e61d7a8b2");
            when 1272728 => data <= (x"3cc5a3e7033dd3db", x"15429397eb270bfd", x"f00c26f3aeb7a79c", x"4722efc4109c9709", x"96dd4072493328f6", x"5a6338362672b844", x"7f8d163bb0cfe8b4", x"d4d279ad9000f6ed");
            when 17391982 => data <= (x"907eb0463e3aa8b2", x"e067f8cdb6661a23", x"f177fb58f514c2c7", x"ce81534c99e987b2", x"24503fb0da4328c7", x"5d03f8797c7603ed", x"79e4df75b63e5ffb", x"3fba1d5ffe58354f");
            when 18655624 => data <= (x"93c38d20be5bc256", x"e6b8af157a461bfc", x"2e7e5c47b9020e58", x"f1b6fa5d593d1812", x"46806127930fa6d4", x"b398096bd330b876", x"d307c63593a8789e", x"c31bed45f3947f85");
            when 21999754 => data <= (x"5eeccaad21f27bc5", x"7755f7fdd4c916b7", x"a5acabb37a27b2f5", x"bb66dedf70501467", x"c259294752b1d3b2", x"563f79f1bb573d24", x"19318748284872df", x"0f43bc7569f9b62c");
            when 25785429 => data <= (x"a70b3fc9ee9b5151", x"5a64ace6fe44668e", x"2f07020bac6a961f", x"a61298812728dc6c", x"7a1a326d86f89014", x"bb312c73e40c1131", x"d857102ea51bdf69", x"2c7146a6a6473dcf");
            when 31817585 => data <= (x"d39da954c86a7e72", x"40975abedc99950c", x"771065d9c629b8b3", x"de4d114f5aad941f", x"d9ebaa6b88fe2eeb", x"1860efe892aa256a", x"6f5a4648a98f4a0b", x"b99260dbd444a27c");
            when 16571653 => data <= (x"551cbf0ab959e432", x"7b404d3c26a8efe6", x"0757de0cf6161e9c", x"a6c7e137d3d6a678", x"fe0952042f8b1257", x"a0eb7d7e06048358", x"4a26d2af60eddd15", x"6ab4ea73d8d703af");
            when 7219487 => data <= (x"0874bd8c71d86415", x"58147654fced1fb1", x"b2612d9a0054bfbb", x"62a81e62af2acc26", x"62a85f8105b5cc3a", x"ed05af0f85818608", x"dcac73fae39652b6", x"d9e19ba24d455055");
            when 14970808 => data <= (x"feeebe1f98adc073", x"d3e900828ba70618", x"c2a464fd1498f62a", x"5abb1d34594e3a9b", x"df99b9cff624dc96", x"d2760fae2432dba6", x"2e73d989ff8ad81a", x"fd1bad889adfc20b");
            when 13219456 => data <= (x"6d8ee5a54b3df315", x"5d6f034f75eb5eb8", x"8d5c13329bf3d4c3", x"71b801bcd980110d", x"45976eac1285327a", x"90506f93e071ad14", x"9baeb054261c9ba5", x"2af210e44dff0e75");
            when 2197461 => data <= (x"43c7ce47c501e59d", x"c0657f57c76b0b20", x"adc7d0cc43d3703d", x"bda8590d8130cb4a", x"6aca8c0ea7c7dbde", x"4bef9a0c01ca15c8", x"2735f80a4dfda505", x"4a48b0b5b75dc9cd");
            when 9808674 => data <= (x"46700b1377c1d8b2", x"64efce5489aa6e44", x"94b2c451768342da", x"f03768d80069602b", x"7daa53bd675b13cf", x"a7a31564760824e8", x"87d01c0eab4855f3", x"39c211849f90d60a");
            when 8005011 => data <= (x"f0c83156d17a9fac", x"dbe32a8cbeda4183", x"06eb7698cbf70d63", x"e9bd51d5321467a4", x"4c16fd4f17a2c15a", x"46c1a06b5ff91dcc", x"1ead0e6938c93429", x"1f5fa9e423cde2d9");
            when 30550043 => data <= (x"e7ffa9c34cca1b78", x"cc9ef1471762161c", x"35365c138ee65378", x"a73bc82d769c2612", x"328078e81ad21ded", x"d1093656b47f34ef", x"5e55168307c49bff", x"625809d642f9028f");
            when 10203845 => data <= (x"6d144ccda1d286ec", x"3aae17eef282ab28", x"663ed9f232084428", x"a6081d77f04cdeb5", x"5f2da98bc63c7be3", x"0eceb6d5f460f2e6", x"c0eed253128b0c24", x"a30a5767e70b1bd2");
            when 8791226 => data <= (x"0a4048a87e1759ca", x"9e0e859e85f7694e", x"bf6df457968ec72b", x"86fd49307266d55f", x"03410ac770419f15", x"94e6e6fcc64e9efd", x"b87ae76e30a3adfb", x"1855278126c46d46");
            when 7101858 => data <= (x"67902d7b53b7f175", x"6eb95d6c7caa26a3", x"dd930a8aba355a20", x"53ae1629b07c547b", x"f3422588137e9528", x"61c5fad4ccdec937", x"9159d485c4d61ffd", x"cca9697ca632198e");
            when 9656381 => data <= (x"5f8bcb3e2af6f5d0", x"84dc53b74f2b4735", x"c5f4f4d8b0049a38", x"273449c3e65200b4", x"d7142766ae7668da", x"12caf1d718450743", x"ec4980d2f0d4bb9b", x"72450e5c4fa7dcb1");
            when 20469778 => data <= (x"9eabd36518861843", x"83ba205dda1f5119", x"b6f499b95d8dc5b3", x"badc19650697db60", x"1f129e6fc13c4c82", x"08a2415e92453c41", x"92cd6832f5c7e0fc", x"b7a2db93406668fc");
            when 31004467 => data <= (x"77004db43a054b8c", x"293504e54087657a", x"09e84f2bb18dc2fe", x"c4e76c63cde1f9dc", x"0f9750ed59d87771", x"cb723b81899acd94", x"20822cd05b67f101", x"faeb57bfb798e6cf");
            when 23247307 => data <= (x"195500833300713a", x"67d51c87fe4d83e0", x"c79486b7b1e1e9c0", x"f534e761e84c785f", x"84892885320b4019", x"7e6db8cafe1416fd", x"386d05b01afc0aa3", x"b1a809d28a10aa24");
            when 33519179 => data <= (x"46731eb0c1deaa03", x"3d38848cc07e868a", x"752075a553fc9146", x"837621b5e291df2d", x"01e1ee8f644895c3", x"3ad16af9f9b8c1aa", x"1cebad986a455523", x"d3306711e97532ce");
            when 17973571 => data <= (x"b47ae765d99ee17f", x"2ee3fd2318b35487", x"7acff62312aa86f4", x"25d71b01478f6adc", x"938262f5c8d14a25", x"d2aa3e97d8128542", x"cbdbdbbcc3e9e545", x"9a34c351584d8334");
            when 14750173 => data <= (x"014317b82ea70740", x"dd078d478a396574", x"9f92812c4bfb00a3", x"ec46811b53370e12", x"4b29d68327cde6ea", x"b544bc14e224bd74", x"98107965409b31c4", x"56e6688a2564cf12");
            when 3942417 => data <= (x"4703e49c6ff724c1", x"fa4e1edcce8c9ed6", x"7b12471d7774a252", x"9830b93400e9aff2", x"5be93d9bab07011f", x"fbc019d951f9c440", x"a20b41d88d746823", x"0ec6b3a4478962b6");
            when 19135127 => data <= (x"b7288df4a11dd31b", x"ba890c6b6f211fc7", x"ff6047824fddccca", x"7a84efbae95f7799", x"f51e5dee1515f07f", x"fd8a217991684e8f", x"1392053bfd63aa3c", x"9b05b60a72d982c5");
            when 8194992 => data <= (x"43bb5042001ba6ad", x"ded8f5f2a288d709", x"1559f56004524561", x"5889f06b65aa0f91", x"8e2ba193a6410a00", x"e39285e0418b5602", x"312bcdea9c7adfee", x"03f8c6f290e97149");
            when 30297921 => data <= (x"eeeeb89406311844", x"0c6d87a3daed276e", x"d1e8dfc1a5cfbc7a", x"19f64a9022df0785", x"75024f364bd58378", x"9a4006e88f282d37", x"eebdb89b1ac122be", x"e4f7ce6ffb913b98");
            when 1180530 => data <= (x"114787d444171711", x"0a7535d90e23a22a", x"7fdc29c30291a75a", x"a0b2b1a40447a2ee", x"c5e29c772ee42ecf", x"72c8e39e0a79715d", x"025156f61ac1b8ff", x"e00eeb8d94aed86b");
            when 10475451 => data <= (x"ecea98008903fb34", x"b1545dd7fa648910", x"a93415a8d452bc76", x"4a660c09acd9022b", x"5560ddb358699805", x"43e8848bab1d2f15", x"d1a74e02da64b699", x"44011c3a606d70d0");
            when 22399556 => data <= (x"23e9f90e4d38c049", x"7189d776e5e2df86", x"08f0323ad5d50385", x"c4767430340767fd", x"65e18d8863a153e0", x"8afa5dafe3633bdf", x"6354a7145d6840e3", x"145d359de5e02022");
            when 30322503 => data <= (x"dae9871c993ba807", x"8db450b5f57fd1dc", x"5edee57df5c4b155", x"8b0571f32e085ef8", x"09d96bde25e7993f", x"08d8e1c4f8b56fe2", x"d8367af5dc159b34", x"427b76e2b4c2d665");
            when 11598979 => data <= (x"129410fbef14ff5c", x"b3ea1d0cbbd14136", x"8296c8c73e0079b6", x"889e1b2fbed9ca9a", x"3630d5ea93d450b6", x"33e0d0eda64d8681", x"fa2a89215b27aec5", x"c898e5348724086e");
            when 9587616 => data <= (x"d2c84fb33c4b4b2b", x"f78fd3dc859b45ca", x"6f5674a83c95bbc7", x"689b8ca1292ad027", x"d8178cd24295ba96", x"3d08263f1c449515", x"8475ad8b39cd2db8", x"e696215fad8fbb89");
            when 11532132 => data <= (x"e62120920a7c5819", x"06a279d208610f5d", x"ca48e7f8e0dc4507", x"156b595066afecdc", x"a7e880c2cafa4cd6", x"1d7d34992f1a6a0e", x"e83b713e0e125fdb", x"80e3af66c9a789dc");
            when 18551296 => data <= (x"cdad78bcaba1a7a8", x"52572135f755d049", x"929d7fb2f6cedad2", x"da5e98defef169b7", x"33d78fd8a18d3701", x"65bd1eafc92eebe7", x"cf90bd809d67e83d", x"013b928517aa45e9");
            when 10973352 => data <= (x"d94064a176279e60", x"1bed63afc0871d67", x"4a3434416a92b90d", x"956b3ff73b4bdc82", x"d860efb781f61fb6", x"30bea7db81c1d822", x"b2b547688bf040ee", x"46fa03be400d132e");
            when 5603282 => data <= (x"33f55c095e2973de", x"1140a9c744f00fd2", x"a0bbffa07944b0c2", x"fff90c254f7b6832", x"317b1aef7222cb87", x"573c90003ebf110a", x"e7d20f16f59b8c59", x"f2e34199bb81fc66");
            when 25875304 => data <= (x"24f338e67594468b", x"5b026c6e759d4b56", x"1f08c21995238bd2", x"8ce7ae8becb0fad3", x"0e274de3ac39439d", x"130347e7e81f72dd", x"76d682628dd705cd", x"9afc519abee3082e");
            when 27290825 => data <= (x"f1475c99bdcaa289", x"8617f2c7b7791625", x"379d7b70717aac6f", x"2cc076b242eea3d7", x"a98dc73f650cf36b", x"fb8d2c95840fc8aa", x"4c793e565681aad0", x"a0042521f791149b");
            when 33850043 => data <= (x"13d5d0acc891f224", x"813bfb029f08e93a", x"7edc9cd3628ffc6e", x"455d278048107008", x"31095c69f1024374", x"72ff2f42330d4b6d", x"98612dccc5e7eca1", x"8512855e48721a02");
            when 2940276 => data <= (x"ef168fce7a8f8d30", x"8660b940bb4a52e1", x"d9c660102d4909e3", x"6624d917d70576c9", x"6918bb41979d1409", x"da6ff7b59d79c071", x"d4c704cb7be418d2", x"20cd332d2f88d894");
            when 895919 => data <= (x"8b672251a75495fb", x"69740c4b6961fc46", x"12c51cb2a271dfa8", x"cc0630465ce70e67", x"1e299d781f30a5b6", x"38f7ada6dc6b020e", x"d1f44537666d9ea7", x"b1ef87e141088d9b");
            when 32220948 => data <= (x"0c93f0580c297366", x"7f2fd761865fadac", x"e56de83ba93fa171", x"dbaa58db51dcd48c", x"257add2f52a0e2ce", x"4f790f02851236db", x"d3d25d9c89580202", x"2f0a6fd8e8ed497f");
            when 27068594 => data <= (x"d2e725f9391630d2", x"aac7fd15fd2d4eee", x"21f13cadb3da27cf", x"96fd1fce9a63a962", x"a2a8e8dd6361ffde", x"116d469d317ae9d8", x"46c883c54280af95", x"6d28d579e2ec7d3b");
            when 1163948 => data <= (x"1f561e7558d03421", x"81cefd2840883701", x"33fa8f972861632a", x"dcfbf422688fc9ca", x"6cfb620542b2c615", x"ffb825f13452cdf7", x"067533cb38b2b805", x"07d2c3f7f5cc20ad");
            when 5372394 => data <= (x"a844a6ae85a63643", x"a84c71407412e46b", x"9176fc8bcc514176", x"9d7827840ac9e660", x"483f49c5ec725447", x"05f34b7c6b9697b5", x"9625bf6a2b38d0a0", x"e4a5f04b06e6512d");
            when 27484113 => data <= (x"b9f0bb1d51b4589e", x"ca5ea822129217e3", x"2dc1c64fa506df2f", x"fe80798751cf5817", x"8718a4a58177bfa1", x"33a73ee4137e1f6e", x"f437b64ec9b3ba1f", x"5778ee5cc5afea8e");
            when 15842095 => data <= (x"8ff4d2db8345f43a", x"f1c7bcf4f9dead8f", x"1e8405ef58421170", x"889f788ef5d1b00f", x"08186f11aad5a981", x"2517edd35ea1736f", x"c9bfa0daa351459f", x"ff0c42cc96a22619");
            when 25296395 => data <= (x"48567a643e9106a6", x"54d7200f045836b0", x"f3ddcaa11408033c", x"97f19848bc5cdec9", x"9e5a41bdbbddd59a", x"c46861cae74e5cc5", x"49134354c9295e82", x"5ad9b3ddde26113f");
            when 25577384 => data <= (x"45d7de3689d55420", x"5fcd8b381fb9f146", x"5b2770cf7244aa65", x"faa621146e7c58b6", x"69a554808c35b71e", x"5b53cbfbfabf256d", x"c04c25579c59acf4", x"184ff623ef96ef51");
            when 29124210 => data <= (x"158dbaed2d52ecaa", x"e7e95eb2ac7a8b64", x"a4b8648d2bbb85f6", x"8c6c60066991be0e", x"1e99f489a022e173", x"dee0785d76f128fc", x"f30eaa001a5df927", x"54c35089e46e7aa6");
            when 10625646 => data <= (x"6d52846c03da0efe", x"8eb243b3a462c32e", x"46b046670557e0b8", x"2105c66500af893e", x"58e2fe8ae367414e", x"6fb1a17f7279d037", x"24bb174a6f68ba00", x"d2c1d96c2f417555");
            when 16328585 => data <= (x"7812e1575a192113", x"3cd248fe0f279311", x"81a566b7e42689ee", x"3dc4f3daf289c956", x"839a0cd7171ce865", x"c1443de69d04b8fc", x"02a229c775ee3edd", x"6c9f1c8571f4274b");
            when 31199596 => data <= (x"91e9d4980adf1b91", x"8483136f39356d28", x"440abc885c846c72", x"7cfdabf9e56c28df", x"9848de460921532b", x"0f94558055f97986", x"259c681b8708374e", x"a5e86f713b99f408");
            when 391545 => data <= (x"ec4a3044cdd00c2f", x"5f20fdc230d47b81", x"ba0fec9f4a8b0d86", x"d10abf383ce6a603", x"efb3fa59383dbc0e", x"2ce98739da28a7a0", x"6cab145dac52b537", x"27978c963145a0cb");
            when 19813695 => data <= (x"1acfa6f86815c3da", x"2eeff7f246a5bfe7", x"bf6d360c4e07aac8", x"81c7eb9e7c741c6f", x"10f7d496f1eeb283", x"7d1aef4aa2b903f6", x"0b936b25081de8ad", x"4d258549b2b49dd1");
            when 14683660 => data <= (x"00905a859bbcc1a8", x"247d5ad516672b16", x"57901fdd3d56a940", x"65bde19c3598623b", x"07708a46264de834", x"6388be3c7c14ef72", x"9bf69e8506171adf", x"55cd8039a0944419");
            when 31509227 => data <= (x"ba8f34ace1bb3728", x"bddbe4185e4b58d8", x"98d3f2f5878fe98a", x"471403bbc711efbe", x"0028dc75b479cd8e", x"612f46dc71838351", x"61fb0cc0a4fb0f40", x"c129ef09a5e91f0c");
            when 14607214 => data <= (x"3bfd0991269cf574", x"06b91c5a3dc60d80", x"96f5ae9e39ad4495", x"8f5980c554847ed0", x"ef30c1fa1701101b", x"3d9f797bb6d191c5", x"033a0e919c910176", x"172bb0fbf4154bda");
            when 21615577 => data <= (x"9aaa57e08b16ee7d", x"81e4ea8cc188de10", x"de8bd14e5a6ae72c", x"8e94ef156f33002b", x"212c3ff3b70a177a", x"9cdd38b06cae5e73", x"5f3959602530d76d", x"77c36c5c98f30bc2");
            when 33416122 => data <= (x"219d5d605ab4069f", x"9e934cd2f5700fbb", x"9b7170bb3799c1c9", x"8e140c23732b63a0", x"204479f4de560243", x"bb7392134f63d702", x"b05684ea4de807ba", x"706494c9d5559282");
            when 2549225 => data <= (x"da32b35f5a70f4cb", x"714967450597bf08", x"974131f360c4b216", x"4ec52606c81b59b9", x"96037f9e6b8476d7", x"398ac6deb59bf9fd", x"fdc44034483fcc77", x"46ce629e48496d3c");
            when 2695532 => data <= (x"08536e45ae3ce074", x"686e5beec21ae9c4", x"4dbdf9d1ceb903db", x"a4107b5ced15e79a", x"3201f233b05d9f56", x"1028ab1b7bd93976", x"1e2b8252e528d46a", x"2dad167a402af8b9");
            when 2377353 => data <= (x"6a0dfb6bff279da9", x"31e58c2c2c02a9a3", x"b0251d415eb6cee3", x"16c43cabeeba9319", x"79291e196a30ad6f", x"70eaa6ab78a81d3c", x"6194541439a16619", x"dba5dc15bfdf6765");
            when 3672807 => data <= (x"f2e7644bf4658d7c", x"bf9b120aa873a274", x"1632f2a000868af1", x"df7dacce87f55281", x"e98f60a1107816c7", x"4015a2bff99b6442", x"091599bc3cbf4eb3", x"ffc7ebd150549151");
            when 23791291 => data <= (x"5b2b91a4236a2026", x"af0e400388beca14", x"16824216e8c8dd0f", x"686932b8039c1e8b", x"03b5b3da3a411ceb", x"02cb81da7d1ee85f", x"a4d86f465b211eae", x"8df63eac9d5e708a");
            when 22849850 => data <= (x"be4571e4906ecdd4", x"5d62c76b99f72dac", x"645bb3d4fdd8cad6", x"30c20aad44250817", x"2aebd775e9cb43d6", x"37e6701d210b0259", x"90138f2047e5cb01", x"a371d78bd8ca2486");
            when 26513226 => data <= (x"c447b5a6505f3d42", x"a84ff3380664572b", x"d30996573b56e843", x"0100c4ef7e67965f", x"5b3f50353a6138b3", x"ac98f095efe25cbe", x"b4f866c0d2824429", x"84371222edf70994");
            when 12727473 => data <= (x"24242901cdcc1d24", x"183816f2085e6da2", x"e1a28e68bc22440d", x"3aefcd3ab6a31f19", x"03af66dc9d4da6cd", x"da9d9a3002918bb0", x"079deb5f5ac33cb8", x"eeb18c186bab1b50");
            when 13377606 => data <= (x"ab27e350d378a127", x"36c3ec7b21233a60", x"578372fed7a704e2", x"661a6e7f0c3d4d33", x"891be162613e98d2", x"182a8196fe721a91", x"e6443d911b3dd29b", x"520eb3c1e6979bba");
            when 19115805 => data <= (x"5766d47dbfe60ed3", x"ad2a9be79d339e80", x"3c545ef2379da579", x"a1c5839945bd138a", x"182422819334510a", x"4aba5b958372968a", x"c9c3d53afde19841", x"f61deb5bc6d3a336");
            when 10179156 => data <= (x"5dc267edcce4c87c", x"906cc5f83d9a6110", x"1e1a758522baed6f", x"5bdb18b6c4365ee9", x"85bd5438ca0dbfa5", x"8b0bef75fc222d75", x"904418d9973f8db7", x"cfc66da0b6572307");
            when 30522652 => data <= (x"6b22eafb85fbe3ad", x"dbae038d2334d0c0", x"485311f616734f44", x"f30bc515ff9b3db0", x"9e43d8dce1917678", x"00b80abc1231d27d", x"6e97c867394c4477", x"a3361d9357ceff43");
            when 5365100 => data <= (x"65bad0e31d155031", x"88a00832d01c7939", x"0f5437cb05e4713f", x"eb5ae4bfd1165cd9", x"347cc4d5dcbb7e25", x"ac54965817ff46b0", x"0a3aa1edbb2c3ce1", x"0d8eb48a1a3dd12a");
            when 23083339 => data <= (x"07255daf722a3743", x"db13e2cf7357ad39", x"2f6801965e2ff67a", x"edd741d3ca77dc7e", x"d9650f27b7a96837", x"223d8b8030810aa3", x"730e15e1fc0aa04d", x"460804a432bb0bf9");
            when 8613252 => data <= (x"7e5b59e819e8435f", x"ab199788bde96977", x"50b96f2dc4b3230a", x"b6cfbfd94341c8d1", x"7ec1914be57589ca", x"61f40f53c8aa8730", x"ab941313f9af4bc7", x"73a15b8052fa94b4");
            when 898761 => data <= (x"4d48ab70c93342be", x"a1ad7b540c8099a3", x"d429cae5557752de", x"3fef645291105ac5", x"dc4f8763b8f786ac", x"b2ddb761c4ddf045", x"5c60cd9170c5ab34", x"938b1ad7ca8f2c88");
            when 17853775 => data <= (x"e9e69043473595a7", x"3cbc1a1882d0f546", x"b8ae4f06344d11e6", x"28a74ebb497c24a2", x"44ade83977105da6", x"60787e8b085cbadf", x"6ba2d973768b0526", x"3e5dbd29081260d5");
            when 33804826 => data <= (x"1b53493dea95ffcf", x"5acc1816d6c790c1", x"32b99c3db0ea7a98", x"d2c352b12e186cd1", x"5c0469a9f66f8b2a", x"3ea87bab497eacff", x"8c442fb30107240e", x"b8a3fc06d4d93817");
            when 24080537 => data <= (x"989d5f0c17e2e865", x"cd0d501c69440b21", x"1458a71b88364e70", x"582375c40dbb43a9", x"7bf43c57726781ee", x"ca3ba406165684c9", x"59794dfb0b6d1af9", x"7044d3ce279a6bb2");
            when 23109642 => data <= (x"46948e57f39f198d", x"bf6b3585f15d8975", x"2a02772c92e23d4c", x"4bedcd7f2b216830", x"af7dfa4862b4b26d", x"0c5b3296035dad92", x"b4525029d6aabb24", x"99e4b7659499f252");
            when 16683167 => data <= (x"5acdbf3ab2dac5bd", x"72121752b85da5be", x"1adfd7d52c23a0c2", x"18ffe607719bbc21", x"6e73b4334c5f3d2a", x"26f2ef501f2c9f69", x"f722768b70d45a12", x"5c9507f7d071408e");
            when 27700103 => data <= (x"e89d4d0e81ec63e4", x"d32f30e0f703955c", x"0981a49a016a790b", x"9f38bbed1cff9aa5", x"43a95187a7d1626b", x"ee9b35bc4d3cd366", x"c9cf129530ae5588", x"0f58a88c5b4d2afd");
            when 24383637 => data <= (x"6389b3d2e080f902", x"b9a394e482cd696a", x"b9e87ee8fbed042e", x"4ff2027f3ec9a1cc", x"46d6ab590e9ee9a6", x"04e70bacc5fd70e7", x"374e69a85b2088cc", x"ea0d0d6d9227b797");
            when 9563406 => data <= (x"38d69d91eed30dd3", x"cb81a3034ed9aa36", x"1f53fcd5c7517f84", x"3b18b631300eccfe", x"2ce0f41a34bb6734", x"126d12eb849fc30b", x"f8dd1b7e7cce6575", x"10a0b254e5609460");
            when 966024 => data <= (x"ca8286275f0dc2f1", x"53ae7a2554823dcd", x"b95b40afe9f75f06", x"bbff46567e987e28", x"23c1576478a32e25", x"31f86eb034110594", x"250940d8a6a6deb7", x"1de81c5ba0466a68");
            when 23701445 => data <= (x"fa610f72e4002fcd", x"9e54930f03664453", x"b82e6acad6759871", x"9249870e24478264", x"a608c880fb310787", x"d7651f0d2c25ce0a", x"5b6484dde47402cf", x"7f59b35d3fb9df9c");
            when 30489733 => data <= (x"15feb1729d58a642", x"fbb443b2b07ff583", x"727c290c6ce6260e", x"378471e14a2057f3", x"e22f46df3535d32d", x"d76fc5e1f2b26cf8", x"ef89d01bb6f9b755", x"c97d8594eb925b85");
            when 2550985 => data <= (x"3abd1a4a9ce1f8bb", x"523395e8db42be35", x"35277fcee6e5dde9", x"180d05ec152debaf", x"7b3d6466c5c2110b", x"06c415b978aa505f", x"607ecc136394c0f6", x"fa5011d6bd567ef2");
            when 23273675 => data <= (x"57cfd55e3866d85a", x"8296f9a6e2fe136b", x"68fdcb13087d3a27", x"dd15d9a7a255f184", x"8c3a6a2a674dac19", x"52d2a3c255bdaf06", x"be54babb8b5ad0cd", x"2f8d1156ff014f1a");
            when 4654624 => data <= (x"8509e1eace5bc3ff", x"57181454c5c313d2", x"c9dd3a659048f82c", x"4288bb86e7e31b9a", x"b79cad62fd06c6ba", x"000666d12917e850", x"8d75414d379e4f4b", x"086aac200b75c776");
            when 30477969 => data <= (x"bad8acd3208de375", x"b398f898199b62b3", x"143a399134dc2901", x"14db6df3173e535a", x"9a18170f75b241cf", x"c231b27b3dbba5c1", x"8e9447ffa960a84a", x"b938e33d9ee7530f");
            when 22838127 => data <= (x"6e1d0faa985d9dd9", x"aca0fac10346f503", x"1355f559fea11102", x"c7aa7bc8a8688792", x"c42d4a6835496c76", x"b55023483d3d7d22", x"0d2b466e8d4e5d23", x"a61b1bb4a42df9aa");
            when 33451508 => data <= (x"2783083b46f38f31", x"43afbd13d0f11d5d", x"873832c5d2385eb1", x"9c1e65d4666636b4", x"c3ca1b7ee6ede15d", x"c3ca188ae1bfd22d", x"6dcbf61acd8c7878", x"a939546e8a0c4951");
            when 12934043 => data <= (x"e5be026f7f8bfbb9", x"a8bcc84f1ec68576", x"c006d5c945e72092", x"1837b438fae4621d", x"b4a29a9a9aa03cc0", x"b7985476ac33bbe8", x"d0cfc6052b7eb257", x"df2ab9548108663c");
            when 12315912 => data <= (x"c6950151f7ec7cec", x"6e2d1383b7d24451", x"fc6000cd5e5a07a7", x"ee05165a3d283471", x"b84bfc6df1bdd71f", x"727664f5a16948f9", x"e81de737fcdec69d", x"86096996d7fcaba7");
            when 25409530 => data <= (x"908397099560f505", x"08e3d0c3e9d324e7", x"dd73094f3a6e5908", x"93599a5203d5abe8", x"c8edb9b62bf0c494", x"724d9ff69482f1d2", x"99046b401b827a94", x"af238756ebd06d2a");
            when 10914657 => data <= (x"00d474905ba0bb3c", x"f30cb8288bf16d0c", x"862d80e4a5cd6b84", x"1493dc4f8638fb5b", x"79af2fb75ced9b7e", x"5200d4e8b989cf0b", x"2abaceae81679bcc", x"7b534d09b1b39383");
            when 11823438 => data <= (x"ebbd9c0bd33d6aed", x"7eac2e0a0eb48e9d", x"2a4da3eb3fd7bf44", x"d9c0b3c1eaa8ff2f", x"c359ab6df8ed92a5", x"e370e1b63b25a85a", x"ff6b2bb604541736", x"71ef23778d9ae281");
            when 16613310 => data <= (x"e9a0387f2b2fc092", x"4fbe47c56f477cc1", x"963c3375651aded0", x"f5258ecbe3af83bb", x"254548d8d447f121", x"2d1cc2c43e9a6768", x"68619311907d91d7", x"76472f276b9a3683");
            when 3422560 => data <= (x"3717c64818035515", x"6a684418491fe42f", x"f91c749d8df155ca", x"a1a0c24e47f469cf", x"8578e897ee8d7732", x"b12fa0113f7a6ce5", x"91446ef0029ffa47", x"12c33753cd155699");
            when 31014331 => data <= (x"9d29a152ff2d3021", x"d0befc8149ac8f97", x"a30a7e42d518a508", x"4838c487dffad37f", x"12b2f907c213e070", x"1538d2290bbe788e", x"d4fdaff83f2b0af6", x"53dd5b58e767e81a");
            when 28680359 => data <= (x"f3fb0310dee02594", x"8f96b0ef81fd3a95", x"af7a519bc089abb0", x"34fe23d32ef568be", x"e9815faf5a392667", x"149dfab695bdc30c", x"1c88f6e335a7aa07", x"b30591764ac7081d");
            when 4520955 => data <= (x"aefc5c7c292db8d5", x"73375b32276bb6ce", x"d8d6e338ffff6cc6", x"d3da3561386516ed", x"6c746cb0cd7bb947", x"db595da1f6841c84", x"6723e978e9a672e9", x"4a07ee46de6dd33e");
            when 5230393 => data <= (x"a7bf5c85a8c5fa51", x"85b2206f3e20935c", x"f944798aa7fd0966", x"1fa915aa538b04f9", x"ca90561ff90e05e6", x"28df2fe12f866c7d", x"5c6065d4540e48d9", x"9ad659c63d156162");
            when 12856579 => data <= (x"29c9b0eb2ad6e0c6", x"eb439ab8c4519e7d", x"5aee7a51f90472f2", x"c5d35b88af48459b", x"f037e5fecfa08c40", x"6b1b961ee4a1ea3b", x"21678632e9ef7f3c", x"3d353ed4e61b7559");
            when 4091382 => data <= (x"b0861566354d914b", x"14e5ee5bb41eb21a", x"a513c55bce9ccb72", x"b0c889a0bf54aeee", x"bee26aa2bb0e1300", x"8a307ec81affdd91", x"d18ba3449b610c71", x"279634ad0bc63e55");
            when 16467860 => data <= (x"16353828dbeafa5e", x"fb8087abeb3a5a4e", x"e8f8c59346f43037", x"6aed9a653d9906fd", x"01c7c3f884b13b52", x"97d330e8f228c97f", x"94467802cec5bd4a", x"aac9eefac310ef19");
            when 11097816 => data <= (x"21c2bbea51187afb", x"f785c6ff45015e27", x"b78f88df0685da6b", x"9823389bf6453765", x"708e75356bf4b098", x"0f08991db878687e", x"559e662d481bfe19", x"0f7c41d15a7b5f8c");
            when 30147349 => data <= (x"067be84b10d99218", x"cefb4aba18268abe", x"0c227a5177854348", x"fa5bf414dd52c3aa", x"153ea8dd92fc5465", x"0980c55b6aa9de9d", x"b1ada3d4e0d7f201", x"a86dedb68404079b");
            when 31779565 => data <= (x"221bbcf756c54ec2", x"83f8107fefcc464d", x"50301bb2e0037c94", x"01f9367a48c11184", x"eee3608e54e7e464", x"026a9b2a1d12f55e", x"37062be983e412a1", x"d8a9ba13d981d5a5");
            when 3447536 => data <= (x"137b99134d4f0afe", x"969a19324893f56a", x"e9c9034ae8df113f", x"dd962549535376cf", x"362565925f7458d5", x"b7e3c87f22860c1d", x"d7fb7b79e5855ec3", x"45d7e4b1b0ee9ffe");
            when 9565321 => data <= (x"e5fb4a09986c23b9", x"bd90a9f69958d286", x"d51ef5b1bd7de26f", x"dcca8ad3f04aaf41", x"9ad77830b0773ae7", x"8a8c1b5ffb8d0083", x"ee5915f7ef7cd0fc", x"d0ddfbe766b70d40");
            when 9072083 => data <= (x"9920985518bc4c7e", x"86153e5c3a0f4560", x"c80a4b468725fd3d", x"1536aa77906a03a1", x"09846ca9132193c5", x"c9b9f9d4c4df18d3", x"86f7a7c87a049670", x"47e9cfd7bce11951");
            when 7874177 => data <= (x"816c7c6d92288ce8", x"63a95915115caac6", x"ae996c8dc5acc6f3", x"fdc67a2e0a31e141", x"f2a3bc770cff7587", x"a45a8931f16d5e78", x"6d670cb30b3afd09", x"ceed6f1bdca056ca");
            when 13021810 => data <= (x"f83652a1768c9913", x"38a6f05e83b8a298", x"890f6272bfc55360", x"3c0df6063f8db7c4", x"8917bedeb250955d", x"d7ed856d041cc32f", x"5b28b01ad1c53b94", x"4f3f43519fc775c2");
            when 12375418 => data <= (x"c3cff18bf5ab1553", x"bde11070fbfb6cb0", x"ea07c461a8806d6b", x"94ebc86215d5010d", x"d1eacc99ba056421", x"7439f1de9a95a199", x"7cb4432ff4add08d", x"6f7278e621c6562d");
            when 31201071 => data <= (x"3e6bcd27d4d15d4f", x"617d34aed7e2fd78", x"546585b66453de6a", x"7c82b7badfc11986", x"25de8c0defd4e77f", x"8a8a9d0d650854c9", x"6a13f7fb430f352c", x"346d4a917e81079e");
            when 11246212 => data <= (x"3eb606f32f426f94", x"7b0d60b5fcad92e9", x"76b9a8a2b08bf19a", x"ef531facf1942669", x"70b7387d1db81dfd", x"2c4e3c8e5c8b6a02", x"204fd3e2d1c95986", x"a1a2a653558fb532");
            when 11373578 => data <= (x"6a725940ff8e708a", x"860319e439af38dc", x"abcc61136647df09", x"7c2264c3b7a0d4b9", x"1b0ebdf988bb9ab7", x"661511f3408a4812", x"97be9b51439deafa", x"e7048264a7937eaf");
            when 26585398 => data <= (x"e3a87d609c854ceb", x"4cd32ea93c5a8c49", x"3ffea2999fc6d8ba", x"48591f6a653eabdd", x"1449dbb5afa843e6", x"2c0aa910ffb1ef86", x"1b5d8fe23c47db8c", x"764a599f1a032dbc");
            when 4686888 => data <= (x"35630adf0906dd5f", x"8856fdb8d5b6aab5", x"27b95ed78f20f161", x"8b76f040558f33f9", x"322595cba42e54af", x"9561b797e2f9906b", x"3e2ec473badd0745", x"d9d78400761c48b1");
            when 26942296 => data <= (x"caf116e9671d8280", x"bcff8c10a05f0efa", x"3c6dfef37aa02287", x"dab2baa932b6331d", x"7fab2695cfac51c4", x"e08b9d8cf72c0c0c", x"7ffff20577094bc6", x"8db142b3b253406b");
            when 19814782 => data <= (x"7a1801104518a55f", x"747a6dbfd8f1ff85", x"e4b135bfb925bbb0", x"d0804acb79099a57", x"fda87740795eae82", x"98cfd1bd0df84542", x"ce6f541856b73583", x"1709eb19469a6d50");
            when 33377487 => data <= (x"c871a5f284e70f12", x"2faecdf0773400bb", x"0062604464a8a8e3", x"9fc65994fd1182c4", x"4ada89dac479dc59", x"3945a8dd8546fdaf", x"681e67eaf2417deb", x"5a56a730fa56a3f3");
            when 3084875 => data <= (x"32f2b2b69c834656", x"c40cc04a9dfa6995", x"2cc266d121f56292", x"4899caf7524857b0", x"9cf63eab09329aee", x"034a715a52b03d39", x"60b7713694b420e3", x"736e19d9deb9a527");
            when 27390946 => data <= (x"6b8f4e6d38ec7f01", x"5d63ca4bcbe891dc", x"25168ac6fc99aa02", x"f9c56b6cf604d431", x"a7f9c8f43f873c84", x"14ce8accc46a1999", x"430a61ca8c1e823b", x"dd87307b8cdf6402");
            when 9541258 => data <= (x"294ae9e8f4007812", x"dc17824cbd1e26aa", x"f5b9ef280300bafb", x"bf6bec2a3fe1905e", x"9ac5463948c72585", x"8e3ad9de1a46a1fb", x"3079faab2a7a02c3", x"041e44b43ad83ff2");
            when 10634063 => data <= (x"5d6a348e97cd5d1e", x"7c5979129faba367", x"74e112a40299a088", x"39ac4396ffd7780d", x"923fdaa9c25217bd", x"76ac022606d62858", x"a3d5d7f4d8c6c2e3", x"3ad085c3ea41fd1d");
            when 15051888 => data <= (x"7f11ea0ecf6e2b60", x"44dd7de1c0e3ca21", x"ff961b377d8782d3", x"41da6dd3b2067e43", x"c9b1912dfa8b054c", x"8a93d627f30631a7", x"7ba8834fa44af99e", x"4f52f7ab2b132dda");
            when 29806676 => data <= (x"6520d101acad1dd5", x"6591ae872640c5b4", x"d489e2f78a29fb78", x"8de24bcf72ac79ec", x"b953571f05b7454a", x"ae15a9ec6c8dc697", x"2fd2893719b9d870", x"336f948b0f67a499");
            when 25680228 => data <= (x"73629f290ca1dde3", x"246c0c1cb6340a21", x"4985949f86be7c3d", x"ecc7653d789b7c56", x"73b169c7cb728fb6", x"d22ef679d1eb6754", x"adbd7eea6ed431c2", x"7490d1245544c74e");
            when 28607992 => data <= (x"ca7bc7d83ac0fb06", x"d5e0f93bb1e64689", x"e205a50373cae995", x"33a9d51a7372e2a7", x"b788e1d3174b39ff", x"b8b7ebb423825cef", x"4aca4e4f58a2d730", x"b4122d08e1a35088");
            when 2119164 => data <= (x"e7d66a846672d174", x"85c48d0b4593d3af", x"99a15b44a57f2252", x"6bd0f2aae8a46c7b", x"2a56840bac8414c3", x"e117434813d6018b", x"f5734e71949c30ca", x"1dff9735947c038a");
            when 31204406 => data <= (x"77eea1dbabb20eb5", x"0204353451566d98", x"dc917fbe8c53fe1b", x"b3a88d10bbc9ca2b", x"090b08bf10a742f1", x"526d9bd0114f7fd0", x"981355c2ef554add", x"7d3684abb4cd864a");
            when 14369692 => data <= (x"0712be52270c5d79", x"0af3dffcad1fdaf4", x"9daf014e01fed19b", x"6d444eca02e2b363", x"88d69827a264557a", x"dcb1c313c151cb56", x"bf89daff58db6757", x"bf5f60f829af723c");
            when 23569616 => data <= (x"e12c50fec1bf0f52", x"18fbbcb2e9bbeb1f", x"2519394374eef37c", x"02a1d43496da7f9d", x"beb47d6b810b381d", x"998daa4865029be1", x"0d4c995c69a0f25c", x"db6d7677f2439892");
            when 12803305 => data <= (x"651097fdf9a2cb44", x"5af6a95bb7bc6d9a", x"299b998da8a6aa96", x"e63d0a6087121e93", x"5f06d9224ba4a0ca", x"82ccfcaadd7ec41e", x"3e9a3e5eb394d494", x"21fa0bc60da384f9");
            when 5418945 => data <= (x"bb4503670421a1b9", x"b462c2b9ec774e51", x"2a01af8950d9dae8", x"17ae2d49568743e3", x"32f87c388cf6a352", x"e6c8019b2eb44cb4", x"81c17e6080b64481", x"3f271a78cbeac992");
            when 22688885 => data <= (x"80dfd368b3e13400", x"b28990176b049f2b", x"460886b48caddbaf", x"02936cb8889b5df1", x"6366fed49d59208e", x"62068495b051d5ce", x"d54d9c1208ef4112", x"e931a595f0679bfe");
            when 28017316 => data <= (x"b05f76a8ad86c20b", x"a6b61420866ba421", x"f3aa816ccc2868f4", x"d4ff24bbe51fa25a", x"12eb95cdd288940a", x"cbc8b7a5f36b6639", x"4af26c8e3d7adf5c", x"9267e6622507e415");
            when 33254110 => data <= (x"09e4f2531504b21e", x"17dbaf4f75ad3930", x"82a7e3e7eb6ac276", x"93ca54e7f0505d52", x"564b5abfd295c1c0", x"64313de4f3efb20f", x"5e58072bc4849ab7", x"5de6948e5411c796");
            when 19503792 => data <= (x"a4a1710579626f66", x"ccaac9139bbbae1d", x"717d7f6924a7a4b3", x"415208492e1b37af", x"2ad53eba48286a4b", x"5c9bc52f426eced9", x"d5fb60d9faa6d5fd", x"569dc2ddfd56fd1b");
            when 9808166 => data <= (x"a40f18024c408e0d", x"e10c231711300f29", x"71729a31115aaf5c", x"d6c5fbe8af353b39", x"a68131560767f932", x"30584ff211f9ae94", x"080ac73bd1ba7489", x"8d3d96aaf709ad17");
            when 22422735 => data <= (x"708240a1fdbc25c9", x"8a70978bd900876f", x"cdaa31db5b9a3525", x"72887901c1acf1ee", x"c73553f5e2051adf", x"9cf57d13e8309371", x"5014db6b7848f861", x"300e7a696c741712");
            when 25550210 => data <= (x"70d4723468478067", x"a868ac1d1976eedb", x"c5f85f79a5efbb1a", x"3d4976bb589e52b5", x"cc89f5a0287a0172", x"73f9c276b0a2a810", x"2f22ef06ad2ac23e", x"92f5cfac52fc3656");
            when 13205012 => data <= (x"292d9714b20fa782", x"1893b095b7d48cc9", x"1512dd22edfea824", x"2d64835276113e39", x"c73696198b0dfac9", x"eb2c071be5f3a689", x"260db1b25f597822", x"1f00d486566c3ffd");
            when 31780390 => data <= (x"cab483e135c9b209", x"07bfcac7523c77d6", x"c7d871fe78bdfa19", x"6c5ac476162da8c5", x"ca2a70c2b7ddc6f4", x"82945d93aac000a9", x"94348a1e61a12973", x"add360512bb4c433");
            when 1012907 => data <= (x"e86ad7d7eaad6cf3", x"e1dde63c90fc0713", x"17500339637b467e", x"e5b060dae35b4568", x"07af3890019a0983", x"e94c904400a268c4", x"ac4463732dee148b", x"31a7a9ff35632a47");
            when 1189796 => data <= (x"9f402af4394fe59b", x"c6561b9ec4dc4db0", x"43dc09cb66fe88a9", x"6188c6ed0b3d94d2", x"91a6093160b1688e", x"b11547995371a6ce", x"5979bb85c22d62cc", x"92af3cb1356e78e2");
            when 19598449 => data <= (x"e041c329525c7799", x"eccd5c71c35bfe0c", x"002cfce2cca00e46", x"8ec8e98eeecd2ac6", x"fb893c8ebf097991", x"29082821808e1356", x"0e39434cef058ef5", x"d58b2941c2168a4c");
            when 33117757 => data <= (x"a581430829d9aaf5", x"9b3e49a39dd4d926", x"954b67bcd345e0ef", x"34d08a7928d31831", x"6e1613cbabd5b9c3", x"f56159cae5e861f7", x"c3366609e5fe8e25", x"3885bcaf0dd932f1");
            when 6066189 => data <= (x"7510e2d133ab7420", x"7894842ee5991b28", x"38142c7c9e4e9283", x"403428463bec16b5", x"85f6eeef7c4a5171", x"e2a29723eab323f8", x"1cf0e7d4b3f520b3", x"6e8dcfa90adecf3e");
            when 7529550 => data <= (x"469b162136c48daf", x"289152672473c5ea", x"6945cefd8115bba3", x"f722c9f9cd968379", x"015a40999dc59f07", x"d0c07cca02ab4926", x"ae1ae536f0669d6c", x"a65f1ad74cbaf933");
            when 5848758 => data <= (x"d9b92648b48765e8", x"9b9a99571d8cfb37", x"6d8bf042e3197f55", x"b047216ed7cd2ba8", x"5c5fe10837eab270", x"b04d5bfc631d2879", x"fa152c1fe9383a32", x"c7c629053f7faac4");
            when 27341226 => data <= (x"a05db5ad7727e75b", x"29c1d66fa2b63304", x"565fa566f9ed398c", x"fd8e1abadddecb63", x"9d00dd56ae568c0a", x"4cdf1de5335939d0", x"c09987898da225fc", x"fce5fb6ba1ef9e3a");
            when 27502713 => data <= (x"90ea04e3756fb938", x"f4a3440b65da21d6", x"e0d1bae9dfdf2447", x"98c787c03665d8fc", x"d8cc2b62294dbb26", x"8d8b35aeebcd5751", x"56f3fb87763eea8d", x"6a50afd7aeeee970");
            when 19013126 => data <= (x"89759bdb7d232055", x"f46cdc8900e7115e", x"c412af247e265648", x"6ca60505ab8e54de", x"1b421426aa757241", x"7b3a2bc0d9656d10", x"b7d539c77cb90771", x"7674da0ae7b1580c");
            when 12714001 => data <= (x"6af08eb706fdf7b1", x"02d377e21e8ee8b6", x"399afa8f0c070bf0", x"78d57f0990061b44", x"e02a566e103e9578", x"c0a925562cc2c4d6", x"5d379a2412426592", x"bb8a8783d882ea68");
            when 11751468 => data <= (x"e411818c518286bd", x"63423c5117c8d6b3", x"7f348e88b8e4af27", x"8e6769885996f118", x"29217677cb727eaf", x"22a8b0b5d3805972", x"00e14e26d15f9236", x"36b8e26fcdb9d4b3");
            when 2254713 => data <= (x"e56a50410dd3efa2", x"e7ba21b2463ce73c", x"9bf2ef38284f3f31", x"d6ea4cd42e972433", x"e97a4f465d20bd83", x"b78f8a30186fb025", x"e2152ee87b4b19e6", x"d5edb697789f820f");
            when 23926376 => data <= (x"bbf4d4549b3790af", x"ce89ac8671815f50", x"d60be3758419f64e", x"834f743754a830e6", x"08d0261f2cf252ee", x"134f6132422cdda7", x"4aa37799fae37a0e", x"a007bbdf9c54bbbd");
            when 19811245 => data <= (x"264f34dab0b44e39", x"47a06d60eab66215", x"fa9b995f5c0b627d", x"0fcf63fe1269b861", x"7efa7749262225dc", x"1c3bb733686d6461", x"f6f061a4d91892f7", x"e8c299b050d554ad");
            when 18861033 => data <= (x"829d150afec3bd80", x"e8544a4d3e8b8090", x"a5cd2b8b0eb7be2a", x"fe08311bfc5f08c5", x"51523ac1c45ffd82", x"05c5f6ff633fcd2f", x"1b4609f24a8fb15b", x"9b9ba6236d8c197f");
            when 30012963 => data <= (x"0ba9c84ac115dc7f", x"de8962c28fbaa01d", x"e1ad90dd9a917a7f", x"7db321ff22494bf7", x"4589bea640a75c1c", x"4f91df375f22f195", x"08ad298cf71c6925", x"8b46073f58a76af2");
            when 1258251 => data <= (x"4fbfa5e07b1ba181", x"f7c07d670d1febf1", x"2db57df1ead10134", x"9562ede44e8235e7", x"ec8cc05cce32fedc", x"eded9ab48cd96948", x"b5dd47aa02c3fb01", x"ecda40030cc5b1f9");
            when 28834507 => data <= (x"f8833b6e9fe4dbeb", x"149064953b928e99", x"70e0ff2003a8fce3", x"2ad57d0586dc8b2b", x"c4c4ea4654ad2aa0", x"35ea5e65ffc9d294", x"08e01d989d641399", x"cd72b1d9f94924ad");
            when 5646861 => data <= (x"8c4990ced21edb90", x"38398e551b6b2b39", x"624876be7b904d50", x"9dca2388c7a24fa5", x"6a0480d559482757", x"fedb1cac36ad2a6e", x"393984a53579ceaf", x"af5a0033742ab139");
            when 11472503 => data <= (x"54b9687785680d39", x"a7189eb2a4781253", x"fa89d2b7745ed7a5", x"83ab2288f8f1c3a6", x"1083c9812b93875f", x"f0e6514cf544642c", x"5bd3f386c569545d", x"9644f302520fa544");
            when 24308527 => data <= (x"4384bfba2535bb4c", x"0253434287b54f97", x"6b0cae044007893b", x"783ec9b10447ad48", x"e926813e65685a7d", x"58d975a140ca13f8", x"f92943b95dcf4491", x"366731699f0a6a5a");
            when 22573809 => data <= (x"9081329e6bcaa712", x"daabc12c434dee8d", x"1ddbdd18084d92c5", x"9a040c5d7214d380", x"e0c01d1e5d9f6d84", x"3f2f3b63aa3ac2b3", x"ec2833ab9afecb97", x"573f21bff77e7b08");
            when 26050739 => data <= (x"6bac2fd728b20249", x"29f84ac02be7c11d", x"9240811df607ed21", x"7eed7f37640b6cb1", x"fee8f3d111f30262", x"2a20950c2dda92ce", x"e419e16e7240b932", x"6485516207dc5f53");
            when 9820582 => data <= (x"141bbc890f1d800f", x"0268bd4f6c2b8e6a", x"f3e9450ec38391ea", x"b7574788a3c76dfb", x"71813ac66310a4a3", x"760ca2e730b5b58a", x"432aa997d76393ab", x"b158a1e51822a946");
            when 13217152 => data <= (x"5957e6c6e4446a09", x"3d4ccd5767059c53", x"bb858fbdb9697755", x"a5d0d7c49d734067", x"628e624292ffc356", x"b7846042906e3ea4", x"4d7aa0f308507833", x"e37229d83487b129");
            when 2757958 => data <= (x"27d64191a69e3796", x"cf148512288cee3d", x"b6da5664711ad663", x"804b601dfe5d95b2", x"ba40179986b66a38", x"f85b690ee54374fc", x"20fe26e88045d7c8", x"9a28a35758edd085");
            when 32172891 => data <= (x"53cdd99c03f1c983", x"c1bfa5a8fdbe5756", x"1a75c7a67a7fa650", x"df376e8d87f234a8", x"783a802002394752", x"36effa058139952f", x"2e38b7632caf7b24", x"7b17dcda0a1fb584");
            when 26199214 => data <= (x"be534e24d49398db", x"f9ac61a652b33c69", x"6712686c49870838", x"ed2c56aef2426276", x"47bb8b88367d13ed", x"5c4d78b238b18fc6", x"e5b839cbec46d979", x"c60796acf90b911a");
            when 19203916 => data <= (x"01eab5a7b95dc51a", x"b32c438a7068dda9", x"e5506a652e91dfa4", x"4fe97da9ca3a0b3c", x"704ad06cfdbc7140", x"6f0a7b14acb09dd0", x"000909c5addfad1e", x"d38974c612c239eb");
            when 10655854 => data <= (x"707eb0f76994402d", x"36e43030dfd20f98", x"e108efe620d49c77", x"71dfa7c060d0963b", x"6df84e5d0ae3251e", x"13ef878708c47a8c", x"89bf1644cf28ec31", x"35d0a2137d6bdf10");
            when 3955537 => data <= (x"8f6d234e960bcbdd", x"6e2900d17dbda741", x"4b7f5d99e1771d03", x"aeb50a042686a1d1", x"16b33b4548d68a51", x"51cdf179e6fd1e7f", x"4fd07e8027f09b4e", x"f19a775a0974a9f7");
            when 11682208 => data <= (x"bcfe79499ff1eb57", x"29f411329a4e57a7", x"b21483444d6a99ef", x"5189ca8f505dc86b", x"452b2d94572b2df5", x"ecd0c957712b7fda", x"7756cf7b06dc54c6", x"5a9c91525ca9ab70");
            when 27137609 => data <= (x"ce3c114ace668fdd", x"d002315fe1568995", x"fec19c1a0913d7ca", x"d12b478730d38454", x"262c3b0573533a7e", x"67f52be8bf9c6129", x"ec15dab529ddae24", x"3f972b5482f36f4e");
            when 4380591 => data <= (x"23ec2da060a8db02", x"c1e130a2a68e7d1b", x"466a5fcba4e7967c", x"3f204e817990fcca", x"a9aa0316777de9f2", x"1f6e25c946060d5f", x"a1c2b1ee20166d57", x"0678faa8c7e653e5");
            when 30497580 => data <= (x"2be9fca3f12c1352", x"1083557f3797d6f0", x"aa7d386d01c889f7", x"37604dbba4e291cb", x"090b779fb3a98a38", x"6a631777dab21207", x"396ab2e61c1bad9f", x"ebd880047e3946e4");
            when 5874852 => data <= (x"5acaca1b8e0e6b86", x"5e52e3fe768d3da4", x"95da103e36123c71", x"0e78756abba30323", x"e00f3c235c9413f8", x"e52240a726f62978", x"17865b97da0d2caa", x"76339004d3299e3b");
            when 6670463 => data <= (x"b2a6da1be8a67f2f", x"baeef70173104280", x"69fe700cf4d77c93", x"ffc011b404c64bfc", x"c4162f24879a456c", x"cdb6fb25fcd09150", x"8f226ac1891e21b8", x"c56e3df2b0de9c83");
            when 20821054 => data <= (x"d37cc5a23cce679d", x"27d72fd5c8ea5a28", x"4cc4f1910df1772a", x"52373b181bac21db", x"b6911b1a299f9099", x"c1c913e25700adf3", x"049a8d12cc7372b4", x"1e92395b57105dfc");
            when 19019740 => data <= (x"54037d58631e1d7b", x"568516ac707c4f24", x"a7dba5bc6f2ad518", x"ef8779ba7295eab8", x"cb26165e16b0b091", x"8300dfc47fa807fe", x"c871e2382e357589", x"a68e15b4ce14e7b4");
            when 8272871 => data <= (x"f5b008b4f1c71e59", x"e26d3cc9e16e8cef", x"9f193f6ebf809a19", x"d3e8bdb683fa39b7", x"d5d8eb5fd184239d", x"95bee4de0625b0d1", x"a01faab5a43e093b", x"894ba15295391b68");
            when 28075568 => data <= (x"75ff29545b795443", x"02f6de3e9cf5d839", x"6b43e29bcde8b5f4", x"16cb9339b966693b", x"7686d71cdab64711", x"5ea0d6ed97cc5a66", x"d9503e985fb37aa2", x"6e274b21415c50ff");
            when 13989298 => data <= (x"808ce1a84981fb50", x"572270f67e9d72f1", x"15e17d79eff17e70", x"e7f3e5a83e3a8775", x"58eddf1bb9c56764", x"7012d68b728daf60", x"c9a742fa4ccc4dcb", x"41bc6dca512c8347");
            when 26093790 => data <= (x"ed56746c07fc1c2c", x"b3a7a0dd64d2d4c1", x"ab7dc3cc9ec19aa3", x"282c8954bf28e607", x"1425f0aec2442e7d", x"d1da96d9652afc0a", x"cb0439982edf453a", x"bce87fb7a3dfd7a7");
            when 14376589 => data <= (x"d15787fdd85c8c11", x"f4a6289cebc75519", x"6ecbd300b5ab55aa", x"d58b9f02a079eac1", x"74be15142b27c186", x"2f850ca1d443d9c9", x"ebf6ac5a0b9078d4", x"4db4193bd5495d4c");
            when 4099865 => data <= (x"be795a505d2a4bd3", x"ddaa8cfb23bb1fab", x"348f2e3b9fe3c147", x"7224a05546cc54a4", x"ddd11d934fcf3dd8", x"5644cbd4fee1fd16", x"11eeb496caa1496c", x"c7a247528944aebd");
            when 17005302 => data <= (x"6753c5660aa5eecd", x"7d9a094bc340df9b", x"a19d02dcf659680d", x"b8c19590ccd4c4f1", x"c14f8816de33f18b", x"7f211a1b1d572f7c", x"318bdb2138bcc32a", x"cbddec3694e9abca");
            when 26716032 => data <= (x"e84370fdef8f0181", x"e198e4bedd0be217", x"731a8cfcb6fe6290", x"117d40ee0efda3ae", x"3e87c8c1db203180", x"eacfcf569a1a80e5", x"916c166aac3c95f9", x"70db59287277feb7");
            when 28249374 => data <= (x"14d299b6698c5a99", x"c008f8673030d124", x"c9a92f0454d042cd", x"5a8a094151368e3b", x"c1b73af2165ae46a", x"a4c89b6b87cd374a", x"03b2edde83e2d6ee", x"3d6b46d076ede5aa");
            when 25819033 => data <= (x"113d53b316b3332c", x"7844545eca20b481", x"f0c43173b8fd756b", x"c08041f987f91f02", x"b9035efdfe462bcd", x"a8e369e2dcc597ae", x"ca2249e1f5febc74", x"9c01ada80f9a50ad");
            when 11039257 => data <= (x"bfc2d093bdc7d162", x"cafa9647e47806e3", x"34aa17504e60913e", x"4aff9c6054080668", x"8e3450461bc3f9a5", x"ce1c8e6c57549818", x"8bd0493f3fc2f27d", x"6ac5d2a9143d11fa");
            when 4411552 => data <= (x"b5b3f0cdf9ec1d80", x"aca2053013fbe061", x"7b09bf888033d8a0", x"faa3986eec42e967", x"d9056a4d270d84e6", x"10c12315655f3bc5", x"75865f6213bb833d", x"40a5c17ac9166bbc");
            when 25971025 => data <= (x"086d802f5d7ec786", x"3a2fa870976afb00", x"15dd460895a07ef2", x"30a01e53edca608f", x"b93f9d1d48688674", x"b0e215bdbe991633", x"c527769a6d2105f1", x"e7b978801424e4d4");
            when 987731 => data <= (x"83f5a7ae2b2319d6", x"4d0a1ac1467bbbf4", x"5dbef05531d496a5", x"03abd1c042e151cf", x"c7847a8403a585e2", x"a9c8367e5dd63b43", x"7bd013702c889e70", x"ed36a68d95e391b8");
            when 27208372 => data <= (x"c04fbd6cdb5f4052", x"29af2d77d3425817", x"18df5ea6d5526402", x"55a9e38ac0023b3f", x"3b49dc4875125207", x"11dca455ac0a7546", x"bd017cd01936fc88", x"b4ed732f5efaca55");
            when 16973284 => data <= (x"b892f8a042ec03d3", x"ead536f6b1f424fa", x"a3768efd7652aedb", x"349bcd033d8929d6", x"2ea713a190f022b2", x"e3e5dfd8f6ebe5c8", x"61976bd92b77f955", x"07a57e729e0239bf");
            when 2718204 => data <= (x"231a833796b1bc00", x"e9a53397939597c9", x"7c6acd1fe18b4401", x"372edf247c3ba20a", x"7fb915475eb90992", x"eb6316e5498da991", x"d09d0fed6bd715bb", x"4c0f1b57bf510da3");
            when 17830950 => data <= (x"640a9622c48271c0", x"8f67561af4883ab4", x"472f781d7c5f0546", x"4d9d369b5c8daa9a", x"f32b258f52c5b3d9", x"357fdad37d6cdacc", x"934c19ec244a7bd2", x"765775931865e4d7");
            when 5893308 => data <= (x"aefe723c5e532460", x"7cb69d024c4c6fab", x"59629a5dea33772b", x"4b5bef258fafa54e", x"aec452194277cb9c", x"49b69d5faed4275d", x"ca949df4af5d7886", x"f8bddf2000a144e4");
            when 530042 => data <= (x"35cd7978ccff090d", x"f1825fd536fa511a", x"683df0172f567c4b", x"869267a65f47d076", x"f4a5d33cd2de2361", x"b787654c6ca010b5", x"4417bb680dfd52f0", x"88ee4baa01a73f97");
            when 6559271 => data <= (x"3a91e472d8fd38af", x"7b2b9f7abb10a1a1", x"0863a8d4f66370a7", x"a3090e13a002f6b6", x"44a143683b82529a", x"ad06d1ee50c64275", x"5a8f3ee917e9b23a", x"6972cebf2a286927");
            when 32345246 => data <= (x"12e101dcade646e0", x"4045ac52390d2eeb", x"877cf71b7655a601", x"7020fb36ef24568c", x"109e2176c3a2d164", x"38b984771e6b5f3c", x"0860cd00dfc24fd2", x"698552a6c49d2fb4");
            when 23990170 => data <= (x"bace6f70fa566142", x"e5dd86e7a80d881e", x"560baf06cdef1608", x"39f05e6ae3d72559", x"e0e14d0f041ff79d", x"6ebf6a927e6ca6b6", x"eecb450e8b98a853", x"b62f5c5c134cf651");
            when 11024129 => data <= (x"edb6d80849c02992", x"30de531d301e340c", x"f57a0d0d80be35a9", x"5fe623c74599d5f3", x"b9c498b511ad2e3a", x"1f437e2d31687fc6", x"aac4da3f41d704d4", x"feaac34f78a5880b");
            when 32040317 => data <= (x"f840130016b99a2e", x"5ce9b531e1427964", x"673b924058c78586", x"fbf595b148d000dc", x"2a7322c6366bdbeb", x"82adbebde8de04fb", x"75027e2907844cdc", x"eec6da1c98d6f2ac");
            when 32885687 => data <= (x"58edd0ed7a23bddd", x"9bf780a7c10b59f3", x"5ba450182eacc8b4", x"5634d706c5cd522a", x"965cd337657902fd", x"82a4b113761f76b4", x"ffb790094e227215", x"46134e863e356f81");
            when 24707972 => data <= (x"9b77d2ad5bba13e6", x"ac164fba3bdd3693", x"580f664e672c3b59", x"4f10b5d433bfbca3", x"df357272866ffaa3", x"e845a72143b23a17", x"30ce5c836ac6654d", x"feaf334ddbf16778");
            when 30352935 => data <= (x"f620c69a1a3a1c56", x"cd77df1a32139c91", x"d6599e6a7f5a0875", x"5db946c0ac10ad9b", x"6f0ba4a5beaf09ed", x"8877afdc7f1f0a7e", x"d1b19eec08963d7a", x"3ea1d05c2990cf0b");
            when 11074565 => data <= (x"3ffb79c93857a03a", x"7e1fe1d0ec82786a", x"8dac3861927faa0d", x"f0fd30259d7b84bd", x"2c3c06b211ec1b91", x"39129c392f4400b7", x"794077afd3486e67", x"c5bbc77d79ff4470");
            when 16419571 => data <= (x"b28d830f295784c2", x"97bdc48bbb3d962b", x"aa9a9e89495f7022", x"e548777ed0dd0a40", x"25380a172506b700", x"b3b6435607477b7a", x"9cbeead3f7eda9f7", x"0a814ae971f9ed64");
            when 22132082 => data <= (x"29c098d1635a5c56", x"3e2beedce59a157a", x"130e72c418d4e373", x"2950f815d7c1ac8c", x"2475ecb3fc18ee60", x"cecebe9cb84b518c", x"4b7396d0e7f99308", x"14ce68b7f3a0a9ce");
            when 19580613 => data <= (x"4a539a59f9c38f93", x"3c32a03a4dd33d4f", x"7c95629218e8c024", x"183422d80331e157", x"7196d1fee64286aa", x"1ee6bde918a8e974", x"ec8aea5f19f8472a", x"6f36d8a5a406b6e1");
            when 21495652 => data <= (x"7cb9c39c2e5b4e51", x"88f8e5d922208b7a", x"70be1c066f5a1ac4", x"5fa7d29dece7e347", x"41ba8e76fcc144ca", x"2ad9ee95fe3459d3", x"daa32054341b4a53", x"cee0170150551f34");
            when 17174422 => data <= (x"63bbf1efc24fa322", x"fe9a08709618c823", x"542383a683bf383d", x"c7bcaf674a0c6940", x"f746194ea2b6c541", x"c5621a68fc86a026", x"ec71a26b01908418", x"81dd439261d31734");
            when 777484 => data <= (x"810039c5e3a622ba", x"ba0e9463174e1c05", x"e39a8226c8b90fb6", x"81babaa57e28676f", x"26abb7bcc63125f6", x"b36c62240f0b4752", x"5b2c968d7284d772", x"debdfb03fffe14af");
            when 27762821 => data <= (x"14fe7567891b4009", x"493fa86d5c7928ba", x"b3c5602ad040f50a", x"6dce068c170e69f3", x"46c0eea79a7ef5b1", x"c530a59a90b3a040", x"e429840bb574b067", x"2606483b94ddc46b");
            when 1237208 => data <= (x"7bdac90557957a88", x"04dc71473bfd0cab", x"f2a944e8cd097054", x"6c88682f2d266069", x"c894faabbd14200d", x"fbece9b6604c3bc7", x"ea1d008c61a890ad", x"9392ddf0c7a4eafd");
            when 27114787 => data <= (x"749f5ed2e80402f2", x"49811ed36a47cc48", x"6aa448bc7f1a5e41", x"d384284bd311a5d5", x"d429699525640342", x"fa92aa1bcb4d3248", x"a5179efcec311645", x"42639fe36f683ca0");
            when 6383405 => data <= (x"271a975c6a671ce3", x"35de3e5ee408dd1a", x"f6def6460761025c", x"ed603cfd9fadd8df", x"d6a18fc1eaee7ddd", x"a4c041593ba66872", x"51a19b25e1054e48", x"7eacfe1d247fe4d1");
            when 13877196 => data <= (x"3b1ce586a41d131f", x"f955e035a0c912a2", x"64ba03a11fa8ff86", x"e281a6c85b371214", x"0427ebfa984904ba", x"5573a8ed4ea61201", x"6854617784f6b4f8", x"ec02c5365304703a");
            when 4789530 => data <= (x"3340c52b0d418939", x"788351349deb70d2", x"01ad28bbd15358c7", x"d0a6b14e41eb3ee7", x"2c67b4fd96d8cc4b", x"955e0c8848b65633", x"a77893fa3addfcc7", x"93157a047e3bb08a");
            when 21777027 => data <= (x"e3d8d82f2022562d", x"32f18c56c948afb5", x"0f401172bb3b129e", x"a514a727ee128738", x"66596de8d6524cc8", x"ee0b30abd8fd48fb", x"711d64d5e33a68c3", x"727f5807c7a59676");
            when 20580978 => data <= (x"0c61bee7d02a5c90", x"5edb4dc9996a6c33", x"3397aee7c66062aa", x"52ebcc6fc5f49bcd", x"2da2818fa0b235d7", x"e687bf5d905f6c3b", x"a80e54846ab156fb", x"a62dbfe4e4329574");
            when 33154697 => data <= (x"e7669abd22619231", x"15d73c003a1090b1", x"06a62cc0ed59c1e7", x"fa5e83d271c09196", x"373b4b14e2e934fb", x"9c53aec4ea77c6f7", x"93163b58cc364239", x"a60e7e52e237d428");
            when 11216394 => data <= (x"effc59d0980880bb", x"9786f372e8806934", x"e0477f6ed6c11660", x"dfe93b5f5e2c4757", x"63b9be93eae3503a", x"c49dbe842389fe91", x"07504f6208454a43", x"2a94976e977d933a");
            when 8154424 => data <= (x"635d87cd93b07eed", x"e9669b613696c1b0", x"9ccab106f898ebad", x"9099c1e9b9b0a9fc", x"dc8a99db1ff52e38", x"950333305dc2935c", x"eb4db2ad6d2d9364", x"513ff5bca5a84cba");
            when 15517841 => data <= (x"98bf9dd63166752b", x"13cdb051c0d84273", x"5a78ff382097651d", x"12b67d074b5a38e4", x"8b992e59fafd9c14", x"704e2d5a9e335c4b", x"8926b46df51269ee", x"8aef30b6213d1df2");
            when 29904692 => data <= (x"38cc8b8824c2a03d", x"56cbabbfddbc07ed", x"39bf42749b0927c3", x"3e962000ef371d05", x"6c0fc6cb38af3ecd", x"18e10ff93b0fab83", x"9fc51669176b6798", x"e482fc190bca5951");
            when 30922947 => data <= (x"0f3445d80ec8eca9", x"bcd1b33789817d61", x"788a3ac44b3af930", x"9d98fde4250a74eb", x"d31c80d491936b14", x"4fe0b811a503c96a", x"460ed6be32a10b7b", x"5e136c6c4b825d82");
            when 25032961 => data <= (x"840dca049f6711f0", x"af31b915f5343109", x"cc0f361cb83a85b7", x"d9e09e61d24a61ed", x"b39888e9d806ecce", x"35555dfc5e563ea9", x"043b6bb75c011ae7", x"5153c60c32bfed5b");
            when 20870663 => data <= (x"6612408ee87dce7a", x"8eddf7d0067e3e0d", x"718c3342d0395fc1", x"c78276535c68d9c4", x"d7a9768399367ad9", x"77e98a3326eca1eb", x"04a03d056bda8eaf", x"1b82a1aa0f4b3b68");
            when 425048 => data <= (x"ef0d8dbcd3c18d11", x"234cd808a42bc801", x"76527ab19f4f3b2f", x"c1989f73ebc45fa6", x"dce2353f28a7c239", x"675cc153e26addba", x"e03bb142d75664f8", x"1e8bfad7b9c3ab05");
            when 18124138 => data <= (x"54c4603bf889ed28", x"3e8ef2a5d6975c40", x"14897070ab4f5f10", x"985d768cffcb0dec", x"124af6098aedd2a7", x"ea89b5fb6f2cce37", x"a25c1b59e1778f22", x"c8c504b438dd73fb");
            when 2751755 => data <= (x"3f511a5aa6ea1a16", x"c45a749e6ba6ccd1", x"49b1bced5b0322eb", x"8ac8616f074b8325", x"22fc2dd1508b02ff", x"3d908145ed83cae9", x"97447e5231cc9008", x"c20cadfdc7bd4b56");
            when 17810209 => data <= (x"35bd78d228b45441", x"41548441e7e370ef", x"642632bb809da069", x"057bb32150a8f0cf", x"0185cb4d40b9256e", x"58312c00b749eb7b", x"96f00a7cf825929f", x"ccd98c48df61b775");
            when 19198853 => data <= (x"f37f0309fb37d6c0", x"83b437dc7c70cc6d", x"8383434bd52b2603", x"04b3ae9b65e3260d", x"eabba24e2d656341", x"a98f64f2b5657f3e", x"757ec2ad74c374a5", x"b9a4e8bc186e275b");
            when 24714497 => data <= (x"20ac0198b3035e91", x"5f601ceeb5835dfa", x"597c03ac9bb05eb0", x"82a6e4dbcf5160ab", x"b2ed01c20eb9d138", x"a1bbde080b7bcdd9", x"c34414720f1a28da", x"57e603676f559d97");
            when 15730096 => data <= (x"7a260d4e6c53ea74", x"2cc1e7c5b87ea06f", x"3288898649851767", x"e75494403ec4f89b", x"73084e1362bc6da0", x"38703665c16dfefd", x"79b213267baf8b37", x"0225e6dc9cdcb417");
            when 3872036 => data <= (x"b0435f0ef9e54209", x"9cc1037d443ceeca", x"65e2d23fe15b0428", x"d69b209677470339", x"3727fc0b26831c21", x"9fbcf044315a623d", x"a3ab46736f1024dc", x"bc0b80cbf2ad7dd2");
            when 6463822 => data <= (x"5db8902c6b003273", x"dd62f37a1cf5f09f", x"4d8ed0d0fd11c4d2", x"2e0583da503207f1", x"9fdf6716873b7c37", x"d48409afbeee036f", x"e88b082a9fec2da9", x"15533353702826c9");
            when 14373223 => data <= (x"b82ec3ae48a441ef", x"be102856216da90f", x"67965a3ed89fccce", x"9431aae3e3f21cf5", x"753c90366190ed7a", x"1a4b360640b01a9d", x"e5827b02f74d9b44", x"ab8455fb8fc7b336");
            when 14704395 => data <= (x"8c7ff917e0163bfa", x"902c4aced0cf6c89", x"cffcafbb18f6dcdd", x"9b1b9960850520e2", x"6126bcc4dcf937b8", x"5356ce1e93b61df3", x"ba78ed07c0561636", x"b569e9662c8fc85f");
            when 816677 => data <= (x"9c1e65c3cd8af6e3", x"ab3d3d126dcc7b63", x"3629a71df68fa7c4", x"13c63bdbc8bba24d", x"7e2e2ad7e5b04503", x"c0505975573cc265", x"f63f7b5f8cd53717", x"f05214810b77b686");
            when 3902096 => data <= (x"1c612c9c7986a84e", x"3628bc3c6216eb6b", x"19d3df0e5aadc204", x"9c8fdc4cb7c91f36", x"95ce5913123872a9", x"2b5483f7fbdffc10", x"6803a434bfd9454c", x"b942fec97bd83bb4");
            when 25164834 => data <= (x"12188be3e8001a21", x"9ae41748bf580921", x"fab6049d03e3700e", x"7f110062ee81b4f1", x"565bfaeea6d7adf4", x"ae19cb793ab9c8cc", x"2159ad5ea121051a", x"582fd8a6e864e86c");
            when 27962153 => data <= (x"d97257c7d9c6ae25", x"0e4310490f32e6f4", x"03d8c8c8ff4ccf60", x"a4aa19cc3a00a91b", x"4c471f42078903d1", x"3c07d2142423d369", x"3eed5272b7d259c1", x"ba8d0db6509fb2df");
            when 14433131 => data <= (x"08e20eabde30cce4", x"2a60c9f23367f86e", x"ec248f4bfca10d65", x"451b58c7ff2c0f78", x"3c938cfb3af54d23", x"3882edee882e7d9e", x"106396843e2d348d", x"2ea087a4c5a835d7");
            when 25792216 => data <= (x"ef4fd4adf505e418", x"78eee66379e51085", x"769969423d618ec4", x"5cf6734d06de8a4e", x"80cdd844de94e520", x"0cb3728b6c1cb3c6", x"6ba5fc04eab1bc8e", x"0cae9594bca7256e");
            when 1142612 => data <= (x"e1f4fa5a0b442b21", x"b497d004bb955486", x"dc52bdedd70cebe9", x"e489166a32bc3067", x"59f0cf5c081be62d", x"698db11b35895f50", x"ce2f7f396454397c", x"6062a1676140d274");
            when 10699075 => data <= (x"e038b2f80bf059da", x"4da6d55b328c21a0", x"94584a6f452d27af", x"602d7caee8a36423", x"014bcbb9781dec63", x"54581140b4a2b629", x"ab02ecb0c8d28431", x"5bef2eb04365b97b");
            when 22245581 => data <= (x"5e4222f9c58ceb67", x"321e5a86e9460906", x"7246d496a01e2f0c", x"0a11b6937791ae17", x"28720f448f2baec4", x"d765d1c757ac3d60", x"9e5a670e96b72e81", x"aa9b0f42fc2c78cf");
            when 25748590 => data <= (x"6a3c4a6e71521cf4", x"1cf2de449ae5e12d", x"ea1ab1681e43cffc", x"12e7f0f662992a61", x"28dc5fed59a0e40b", x"c9f1e155d48cfeb2", x"04911d0a36998d64", x"2bd8cda0128ceeed");
            when 3807355 => data <= (x"e9b01623812ba803", x"b6bb86c4465edf71", x"d94c398c854ad35e", x"6daa1f0406749151", x"a4823d47e738b610", x"dfb88dbe2c5c68e8", x"d49ef13d4cb446ea", x"3af22164926ce60a");
            when 22543125 => data <= (x"7f0c1433617efbf8", x"b188479b2d175119", x"5850de3f35ad61f7", x"5353f8dba7443359", x"0142625f7e5e12e9", x"6301b8cd179a5cb7", x"15a3e979d93734bc", x"a744bf6c3b8db08b");
            when 29994227 => data <= (x"8ecc5145a4b1ea0b", x"c87570c58493c403", x"6e47eb6f99d5ac31", x"a270d7ffcce7a01a", x"da1f324927a5e6ff", x"f749bdbd1012b944", x"c95c58f6ab7ed157", x"d3021ca6688fb3bb");
            when 26670440 => data <= (x"326e554be60a13e2", x"1323760cab4ab181", x"1ef0677b636a3ac7", x"2fef9ee22ddd7abe", x"a8a45d7cf9174be3", x"386c08d5983eecdd", x"60ba217b27521a62", x"0c0b15452d6c913b");
            when 28218361 => data <= (x"369401a6e5fbda3a", x"0c15f95a468eb0b4", x"f0a982b785843e8f", x"2cd2c26b4fb80ab3", x"b197f88400443c17", x"b916635353f4b37b", x"7ff4ddcd624f1094", x"8712494e225f5c9c");
            when 15274640 => data <= (x"3815baad0726357a", x"b0daeb4b9dbabd1d", x"be946088fcd2af76", x"1d3c72964c7fd3f1", x"5a4b26b8f4f8ecf9", x"5012be12e7cf1e9f", x"b9471c4e56acef2e", x"5d97ed8ca8463f7f");
            when 2676022 => data <= (x"674440eac7d99364", x"cc5091b2ff39a756", x"6df05bb39178dcba", x"e747dc8422f065f9", x"7aad0c5bc48cbd48", x"b02ec225fe6977de", x"16c384870f9055f9", x"d9c863e173d0a035");
            when 29933580 => data <= (x"cd98e9fe18676bf7", x"47589b2210f93eed", x"e908d72fad5748eb", x"b8c57ad7c33d81e1", x"f199a8a6971c7676", x"ed7b1903c2a8bb1c", x"01883f5867d00e59", x"9046dfe734d9b682");
            when 2374965 => data <= (x"a51814cfba871bcf", x"071f9c3630938d2d", x"c7932196f4af6e7e", x"7de417c7cbe05e52", x"42cc811e1f2d0851", x"81a264f8abe5b174", x"83ccc0a08068bf8f", x"1c8b41efee1139ae");
            when 10647537 => data <= (x"927a8ec8c6e3a918", x"917c6bbc26456db4", x"15c15fb74151945d", x"717638ece8eb694d", x"95960e6858849dd5", x"57240edd715ceacc", x"55a9276c39c654ea", x"1271bd1f9b98e9cf");
            when 19257680 => data <= (x"28c1036a12238397", x"b1554d617a292d5b", x"7851618e551968f4", x"856406b4cb61e2b3", x"3682cd5c0103a91d", x"13040ff890b82786", x"f67435f54eab3d03", x"160b807163ef23f5");
            when 20070333 => data <= (x"c381a8ca69241ce2", x"3c96b1af5c732286", x"410f607d2b625449", x"e38387727ca0ad17", x"4b2f54a5b81d256a", x"47c9c6d3660921a9", x"e33d2be695cff838", x"785dea9cd37796b5");
            when 30245197 => data <= (x"e4ed44e22a3f253f", x"f6b82c376f7874cd", x"75eaf45621824c2f", x"4b7a38ca06f93fdb", x"3abe9cee61564a66", x"c1e91c2307cb83fc", x"24dac2db6bd114c4", x"b7a135384d76c758");
            when 33456657 => data <= (x"daf100f7dae70323", x"c44383c863bea7bc", x"9b2ca7c5c53c148a", x"cafbec261647755f", x"6520bb82e9bf100c", x"7bef418a28f8a50d", x"e8ccabaeecc052be", x"09619b23f9e6af2d");
            when 11582071 => data <= (x"5f316d921ecc4f42", x"8c8d3a14522e0672", x"c71586a02a239ba3", x"33e4eb0a5e2310a0", x"4cd3c0b04ef30eae", x"2c2c8d47f8def25e", x"f811ceb1141922e4", x"73ccb9569fbd5608");
            when 1040222 => data <= (x"506dc9425c36e090", x"1406df1735ced01b", x"b550b8e6adbb8fef", x"fee02acf2f9e58a1", x"86735aea90d33b65", x"b2f15eec7555ad88", x"8f51c73e392404ae", x"a9590b4e36123005");
            when 8394060 => data <= (x"3ecd970de6302f3a", x"f168055ec6f2a239", x"1ca95625227d54e7", x"3fa70d7236d0cbb2", x"b40ec0d53d599155", x"e03243f13e8d6bd8", x"89b8081322cb612a", x"d8688c618eae8a94");
            when 33083836 => data <= (x"969dbf94dc2d0d12", x"d8c9412f0aa29046", x"cd61cb5a6fecc944", x"44c7cfb18dd80fe7", x"db0f073495b231e8", x"ae3a57cc46253a38", x"ed9a3bea6cffc29b", x"5b0e29f2ab3601ef");
            when 19684321 => data <= (x"a65cb8f3931b166b", x"7991efdcb851a4e1", x"cca51b45bc6c1692", x"b3e9375f77984a0e", x"48389f38faa5eb91", x"55dab9fe65d5f8cd", x"aa84eff93cdaff52", x"7d69a4b3d9a6f49f");
            when 14228352 => data <= (x"54d5c9690872bc82", x"b86dcd55ee94e2c1", x"fda3430d315c5a92", x"052195e11d6c7664", x"92e5d05eb637d45b", x"5011c2589fbcb57e", x"131666bbb8ba4f1c", x"b70b9e5cf216119c");
            when 3198265 => data <= (x"03c7d1dc7c16146d", x"8fdeda2a9f929fd6", x"0d88f2e11c25fc64", x"e8c17c73846c2464", x"5279096324b59450", x"50d6e18758d2efbb", x"06e97e7cd65ce8bc", x"6f7e442e0a0c853a");
            when 16296160 => data <= (x"e86200397a9fa4a3", x"90c5c704d03575db", x"bd520bc5d17cfcd7", x"fec5b2e2e2c39130", x"b402fbec60867725", x"fc28aa76a4c7da07", x"9fe827e0e158fd0d", x"78ed579d4fd146d1");
            when 27686670 => data <= (x"c9255fd2a280cdc3", x"f644b0cc212b8a1e", x"7936d852fa1951ff", x"8f347778512c94f6", x"f6226141865fa3a6", x"9830047d42e9fdae", x"593ad0d3677cf83f", x"1ddacedeb0b6c990");
            when 29554552 => data <= (x"8bf2bf6137c6e2e0", x"3451b6ddc900c95b", x"7880cc80d583f3dd", x"317aafd7662197c1", x"f3151298be0a438d", x"805ef636e62dc300", x"4667e609e8a3ca12", x"909497ea457345ba");
            when 21954034 => data <= (x"182a306cf7a6f669", x"63a03dfc965b1aef", x"f2cbd30ef2d0eb5a", x"26e39a946c157d63", x"7ed674949e15f05d", x"8f946d610d19d3c3", x"e4d9288337e4b3b9", x"8e2bebd56fd2a5bb");
            when 16747005 => data <= (x"36fce1950c9eeb58", x"3f5191c8f677635a", x"2c41ff440c220487", x"ae03c2338464977a", x"cdc6afb482f42c57", x"a830d6c4227752a6", x"7100ec9601de556e", x"a9ebec9139e1ad89");
            when 6102005 => data <= (x"cb74dbaeaafc6beb", x"2b15b61e47432f63", x"517d8af302b135f4", x"ccdc77201df75094", x"501b535f432c9315", x"eccbb194f24862d2", x"3065d9e54a521dc1", x"e4f2b5083cfb5c36");
            when 14344259 => data <= (x"2c99872e29699342", x"8ae82335cabffc33", x"0d086542a9e44483", x"6397a20a5b05e712", x"b3fd765d9d0705d3", x"7cb0a5b73f90bdb4", x"b55a34cb29eb0422", x"f2c5f0d184ec6ec3");
            when 6743552 => data <= (x"dc19779bb1bd41f5", x"b3afff8c92311e09", x"9e409dca42d7bf13", x"a5580404b3298162", x"d2852a30c5737a7d", x"f9fbdf2e1810fa6f", x"bb95340e414fbc9c", x"cede290ec483c283");
            when 3222559 => data <= (x"2d7c956ebac47583", x"eeaf9c49cee736f3", x"0c0f10b342cdb94e", x"fb07ae35e581bf36", x"1e64d3dbd905eb68", x"63bc1bde81911cc7", x"102019d2a3ea2007", x"f9bc741136c88e6a");
            when 11959113 => data <= (x"ff041270cf4d0fc8", x"a538001f0409613e", x"798417c75a251255", x"71fa05a96094b718", x"1882cbf6d3c29c89", x"481d4cfbaa6f4eaa", x"2342e8380b3a06a4", x"84ed2aca4897f320");
            when 4411707 => data <= (x"81b322ef9eb0e8d1", x"0db9fa998dfaa42f", x"15af06e9ca00f73b", x"c6c4dbbb6a0aed74", x"6a2626fc6ff6bfed", x"b32ef9498f0befb6", x"e6b849e02022b756", x"921cd0e132c4097f");
            when 3645445 => data <= (x"c51c39f59d0ed441", x"43f92777ceb0c491", x"2dcd5a0612ec748f", x"ed516b36e3ee42a5", x"27a60039d4eb118a", x"80a88474f7a97ddb", x"5ed583e20778ce5b", x"8e8c9b9fe1863109");
            when 3534318 => data <= (x"81ad30af46077b6e", x"cbd875ce1ed34b41", x"0a5c61e042d7f02a", x"44cbdf49fa2d2eb1", x"c5d5dad4a2eef102", x"ae320bbda692c516", x"f3fe02272fffab2c", x"49fafe19c0c409c3");
            when 9916790 => data <= (x"7e3ce835b3de224d", x"74a361f09872c1f6", x"7e03eb6eab283f22", x"2cea7dbc85ff406b", x"9b53639932a9ef60", x"6e74d49d2a326fc4", x"da512e8fb92a27fb", x"6fe36807b35c2b06");
            when 29741068 => data <= (x"6475b2c902fe9bf7", x"edc4484d5d1a24c3", x"514382c5b6286f08", x"1f87610ec5f0dc40", x"1ab185912d547ca3", x"e8b26f77e027764a", x"d81803d6c903f977", x"58db67f76e441aec");
            when 1660807 => data <= (x"80301b4e4cdabe41", x"63641cefaccda912", x"0565607082fa19c7", x"f4febf8616de125a", x"67aaff90c4a4d775", x"8eb7447f8a3cd803", x"695b128d78bb63f7", x"cdab9b7728f361f0");
            when 1531468 => data <= (x"4c6c4f979885b45a", x"6a892527b77ff230", x"ce5a27b909dde2bd", x"45c71b8036ea8860", x"8f179315611bd276", x"685db9062ed4f233", x"cfd329f701962ec2", x"f73c278cdd7eb2df");
            when 27983414 => data <= (x"f500d83beb08a973", x"a6320cb5e6292b8f", x"a92b798e476d4ad1", x"e3ab407eec36e621", x"977527375477a47e", x"5ae00ea4b95712ea", x"2225c974b5332d08", x"8a05b0ed35bc588e");
            when 26771045 => data <= (x"77b00d1de35b668e", x"11380306ee5c0deb", x"8b5a69d9e0b3029b", x"e32277d7d1011c10", x"bf795d09aa683d8f", x"1b865d26e4cd7ea7", x"c2859a59057483d7", x"e42513388f2456a6");
            when 1571419 => data <= (x"b3a4bdd8dcb21672", x"3cc098427f2cdce3", x"48cb4f612173dd45", x"9772db7bf9257e9e", x"035101bf0e908a61", x"e53be4d14a5ee7c6", x"e6d19bb79507c4b6", x"b27be081c90b2f72");
            when 24199899 => data <= (x"0d50984eedf112b5", x"b327e814b16ab05f", x"b61525a3a763cc1b", x"5f2f475a69d56c87", x"74235c9b2185dcf6", x"66379df5ee2d6b8e", x"9c15b6b4c975c2c4", x"dac252c3be9b29ce");
            when 6798861 => data <= (x"53fcf3233e59819f", x"2527aa7eca2aa2d0", x"9e824152c8d9236b", x"3521cf0b033980a3", x"793221e548885719", x"686a7695885657fc", x"affd88fa6f991b2f", x"6e19a0f2ab36b882");
            when 799471 => data <= (x"3028e83944033bfe", x"3f157a6eaff8fa3e", x"160fa1feacb211db", x"5e9921d96b63d554", x"49c2467e84e7526f", x"08a4eeff810ad3f4", x"d9584d4304a64a9c", x"6fb47b3c09f3efd5");
            when 29949085 => data <= (x"c69ea449974feea3", x"7c8582caca7a5ace", x"dc73733c3290096d", x"fed4ee85eb67e797", x"138198c65fee29aa", x"8aee91d80f86da26", x"ff207d1bddbb7a52", x"0c52d401e37696b6");
            when 21532986 => data <= (x"b7e233075eec2944", x"9d235b88256ae5a2", x"e270306a87eab2e9", x"e1ed2f42092f1f52", x"882e0adb59567086", x"42b3cb441a8944e9", x"ae1c1fef81f2035b", x"f8e45c0b6023eea1");
            when 11881788 => data <= (x"fad553743ded240e", x"83850d883e3d5ffc", x"05eab927fdd43e87", x"c8e79571956c38d7", x"5214ca73f966ce91", x"e1b72d2c65e16335", x"03b06757026eaf91", x"7e8ec4942167ce1f");
            when 33314755 => data <= (x"df152e67bfe47b40", x"7a67055730b172fa", x"eed80ce407e52093", x"eaf3e357618d5f56", x"ac6c46ad821de91d", x"5eb961e22bcabfa4", x"db72d685655b09d1", x"83b41c9a8e76b840");
            when 1194049 => data <= (x"e4e89f76c5de12f5", x"156257d85b6be58c", x"d7c739da9bbaa879", x"4c091e272e56b19b", x"7d3407e7de23ba14", x"ac55a7a05072c55b", x"5bba710e4fe967bc", x"4b57648fc18f54ab");
            when 17385417 => data <= (x"2a66d7f91832c4ea", x"726c4260afb342a7", x"41ea9afba461dfa3", x"14683c3f4ef9f7de", x"19f35915dc96751a", x"3a3abbc27d7eabb4", x"7323ab504cf6e15a", x"bee958d4b8dee2cb");
            when 18611252 => data <= (x"ca88235051ee1588", x"4b82b35f0dadb66a", x"2fe824120c4f5481", x"de57f30d8e70935b", x"962fed8e25797c5f", x"f6d8b858e2d7979b", x"37c847371330d031", x"faa6672e36a490c2");
            when 20088581 => data <= (x"df5ea4fa7e6fd6d8", x"82788f33e787f224", x"293be601b8dd384f", x"ae212a4abdc046a9", x"5dc461ba13fe6604", x"b4b228de6d36dd19", x"a0b3d3eca6837e92", x"640fcc3752c85067");
            when 7550323 => data <= (x"1474aafddd44ec0b", x"95a830ebf147354c", x"b178e2babdfdc963", x"928d1acc25f01395", x"0d317ddf5e252639", x"dc2724933cf1dadc", x"71afb137f09e606d", x"5acafb73cc3aa204");
            when 4945976 => data <= (x"e65b03336fea5fdc", x"11e61836f6148943", x"302bda18fb8b2840", x"07f44e1a6d64ab71", x"0953806dfddce255", x"cd707ecbb77704ed", x"67f8a12aa183309d", x"4192ea880a5b0ed5");
            when 3481068 => data <= (x"a88ee237e710bc18", x"6fdd5f89a964e8f6", x"9b1010b8ee8ef79d", x"5ab0ed93d3ecff42", x"9f4f0a350d39432b", x"16c8c77521e04bb8", x"9101b87fcc14c0bd", x"3b2d204fcd1f36a2");
            when 20790135 => data <= (x"894bed6b18e555f3", x"db6e9f960d75312b", x"6b0a5f6db6bfd96f", x"a708e00b5e1bfda5", x"da4cf5042faec783", x"a2034e776f03dd5b", x"20617626a90896e8", x"b2c86ba3cc0c950c");
            when 22923254 => data <= (x"4b0f627a22ff159b", x"73b631af6ea4a1cf", x"590233070cc27a41", x"efd2f9312706eed1", x"101bbc91cb46ef28", x"ff503029db3f765d", x"babe131e61f71285", x"9e883e837ec04cf1");
            when 12438263 => data <= (x"e8feda0c209b6ae1", x"c21c47db1bdeae26", x"ebdb6f8c43a129b5", x"5221079e9266d542", x"f50b2818bc26d087", x"13ab96c648f11749", x"92d815fbd653a542", x"bf0474be25fd7ea7");
            when 30618096 => data <= (x"2dec29e331ee4e4e", x"7b9e9c8853cbee7b", x"accc2025d0b1263e", x"9e0a7eca826685bc", x"5c305a4de21601f2", x"e410ba6b371a7ad7", x"ffe4b62339336ef0", x"3fea932cbe825c6e");
            when 11873445 => data <= (x"53455ed4aff01d2f", x"b611883ded70d0db", x"51b9fea0b44890ce", x"7116b94ef3c08adf", x"44957d9688e1fd0e", x"d50cfe6c42f15f4c", x"7c71195ff8991e32", x"d1586ce92c9a3ebb");
            when 18518430 => data <= (x"ba868f88252e69ca", x"867b4c81f043eb17", x"69d15945dedc88e2", x"114667d2b37bb9e2", x"b0dbe7246037735a", x"b1d13686ffe3e647", x"7d1155049e354305", x"f3586f0a915c3be4");
            when 19742824 => data <= (x"4d990b8a3ccf4e9a", x"1794fba878463780", x"4d73c81b85a62f30", x"d61a4e362d4f9f4b", x"d509e2871f9e00b9", x"c78e15e59cb8d0b7", x"9f810fa06d8f6635", x"fd9f966301a95347");
            when 15574959 => data <= (x"a01314f024de02ba", x"c9e986f76b2833a6", x"863c4b0b4d084458", x"b2c639770fde2fc5", x"4983b4f6c7851009", x"8def459f7eea61c8", x"5764a2751d9a16be", x"5af9cbc5cf78a86b");
            when 10878021 => data <= (x"4a7a52bbdc75f3a2", x"12dc3fdb426d506e", x"0551dbecb628e09f", x"2a4069065b75bb50", x"cb11777a9e6b8933", x"d34e9682f39c5cf4", x"4c55b8ff90a3ee68", x"5e4f2d3ee9d4abce");
            when 27486364 => data <= (x"9bd1e5f63ca2a6a0", x"8cb9b1f4c49f5bda", x"d00400a39ae62632", x"c4db5cfd637815dc", x"aa84ff7e9c373e59", x"1e16f8fa9b7a05fe", x"3b842171a581be44", x"8b54e3b1ced11dac");
            when 20569459 => data <= (x"0775731e72a68c77", x"7a80582618378994", x"c660ec0ad26b0ea7", x"39bac73ab5064a0f", x"62b4e29ef7de39cc", x"2b2c437a3ff3de7c", x"34a90211abd7d775", x"f70c07ff3da2e415");
            when 19445672 => data <= (x"e7a6cf839cb91436", x"031796869a113274", x"9bc1430425f4c94b", x"7ed94975a63be219", x"4f147a3ee0e7ab89", x"d32abbac38463b60", x"639fe79822bf2093", x"c6ae1558701f709f");
            when 33117727 => data <= (x"1d42a75498c6d48a", x"9ba3da9af2cbb018", x"5a6a2ee680708f38", x"317549d1bf62ddfa", x"49f12c88e71cb974", x"2a25024e03bfa5d4", x"054f69d46c478118", x"3879ab64c55d3978");
            when 595694 => data <= (x"80ecbecf1590848d", x"ae7ee73c779b576a", x"6119c84c4484fed3", x"c1ec37ec3a65419d", x"6c212426e22014dd", x"aae8ab87def9a8b2", x"61d4c8c81beaae13", x"8c856ee20f1d6772");
            when 15413378 => data <= (x"a21efd9219b5afb8", x"5f5f52059a5f15bf", x"2bfae06ee41301f8", x"3dcd2df45914c276", x"752f54adbd52b4a4", x"7e02d5ee6c7e1dd1", x"66950412090e639a", x"ec318797b2a68d4f");
            when 26295682 => data <= (x"ef560d7dcc54f843", x"fe0d1c29592561b0", x"d70fe1938bf3f99e", x"58c131019e65e51b", x"7f926c16eaf53de0", x"edf135966d217746", x"f2a2e4a11e91e6b9", x"54662bb5719a7047");
            when 26181323 => data <= (x"a56b8e21277958b3", x"0004f234d622a363", x"63daaa32b13aa58b", x"bdf67d01869bb52a", x"215f4ab4d1f39ceb", x"0e0351a0d25b7d02", x"672742094ba261e0", x"262b13ff2dd57215");
            when 27418190 => data <= (x"e1b43e9f1813b629", x"4ca03a9c856fc640", x"89e037f38b84f874", x"09e0af13cd5d42f3", x"b6db674147451f6c", x"8660dc568740e056", x"8f99b0d58358ac7e", x"4116719fee6d25bc");
            when 21628957 => data <= (x"8069b8c63033ca1f", x"ffbabf83d6c2d973", x"012d914a27ef952e", x"14d1b099c49d3d88", x"55368202a982d366", x"80822777846baed2", x"72b3749c5347768b", x"c1b3fc6e5a6d50e0");
            when 31635806 => data <= (x"26653b9cf8dbeeab", x"50f7fe1d7710e6dd", x"a69481fb09a0c212", x"1ed4dcdec46fbf56", x"635c06f4deab069c", x"992b8672f00a5477", x"e0958881648bbbf8", x"e38f24090467686d");
            when 30099362 => data <= (x"442257920c143ca9", x"180d7610e4cc3240", x"b681e134c499cf63", x"b905ad038a83bc53", x"2e7bcb6e3313b187", x"1a75110773f8dc0c", x"d0373e069afbb275", x"7d33a1cf51487ed1");
            when 4086375 => data <= (x"1c46204570ac669d", x"c6d19c4108d86900", x"e347cae54cba1352", x"813614c84ff13aea", x"42a2a3d8089aaaf3", x"dac3225adcf79d66", x"8dabeaa61f60a047", x"03ddcc2740890278");
            when 11339255 => data <= (x"c6de9d0d78aa036d", x"83ab0634667cfa7e", x"e93b14900a72f99e", x"6498a8ea1b9182ef", x"1dc1ec5132364f2e", x"65396dd01caf2d5f", x"32f7cc8b49aec291", x"01553950b1cc3826");
            when 10128822 => data <= (x"7be90b54960dcbbe", x"9c4f76cc9e5b8b0c", x"32bc4849b6d919e4", x"508463cbad6c1115", x"c0de2e205876a611", x"ae8c8aa453da94af", x"1a474474b0a760d9", x"164847119678209c");
            when 29332503 => data <= (x"fe4f728a76f084f2", x"c77170fdb02086c5", x"26bc23dec407b0a6", x"546f949a2368f00b", x"37bbd9747b5d3492", x"d71c9d220ffea475", x"208a8021dd20a27f", x"55723519cc2c0670");
            when 28607745 => data <= (x"fb797c6de7d088f9", x"db425d5d8d3d3a93", x"e9337d7fb322b747", x"5fa28c88e5c9ea4c", x"e28687fabe728da8", x"35f42ae3217f561d", x"bda7ece31377e2e7", x"26db98dd5a167707");
            when 31703683 => data <= (x"a532ad4454aa0129", x"aef9f638a8f5ae24", x"98baf22983ba58ec", x"bb75b6f1f7bd73ad", x"4c3da879b8d9293b", x"888f36753e30dc90", x"c025c915d0f7b813", x"8ec4cb495ff712f6");
            when 23462448 => data <= (x"7893d5a1713cc31e", x"d713ef6d89b51557", x"5012923003226c6a", x"e674d2fedb16ed72", x"81599e2ebf8e60d5", x"7aae8dd66539a5d1", x"7602426c11fc638e", x"742a46c814f331e9");
            when 6703857 => data <= (x"3abd3c31bb9f0f8a", x"de569b9ad92cbdfa", x"d7e901a469700dab", x"b99fdd3df91ce1e0", x"e4afd9d0a77e263c", x"b4e5c70abdb65290", x"0c70d49968293a2d", x"ff0528ae287abd9e");
            when 11686496 => data <= (x"c2ee2279da959520", x"e6eab35e160ab0ad", x"bdf4a6a895f146fd", x"68dab0157d1c3b80", x"27f52eab737ed0e7", x"3384a58f68492d41", x"63bc870d8011599b", x"5c03c7cdbccc5b62");
            when 30393653 => data <= (x"25179f20b4b495f8", x"0521961932b8da8e", x"7d42c1c350044ff5", x"cc42524205010560", x"3785bdf638e7593c", x"599996610f67fa85", x"10fcab0cfacce42d", x"316a19cead547235");
            when 25278537 => data <= (x"9d0c124da9e67450", x"875d23bc6214b1b5", x"dc3d1c47f51c0e1e", x"5e30871e01c5c14d", x"4bf7f2f49ce78e87", x"191356f048aa15c7", x"456ff4a6cd7cc17e", x"c3bc7085b699285a");
            when 15071806 => data <= (x"1a81933712d17b48", x"b0be4d40fd29f556", x"a58081b18fe44ba3", x"0ad9a06c80792315", x"5afec448768a4014", x"0d76696d61c2bb2b", x"15be87b078677da9", x"029d18cf6531f455");
            when 30149567 => data <= (x"649535b97cc88977", x"fdfd52ebd8f43c8f", x"549041aa79495974", x"da961beace7b2db3", x"76d016b277bc5c19", x"adddb60d8b861e1d", x"6dcf694bbf292f46", x"0667199a26a6a43c");
            when 33475365 => data <= (x"5462d75eb2810f61", x"eeeecf97c78b2467", x"5a6e02c59c893d23", x"6b0b8725a4c948c1", x"146ad67649d58c3d", x"7dd1e92fe9ea2e0a", x"53bd29857a505f03", x"1502439082b24b60");
            when 23592386 => data <= (x"300b8dadda441cf8", x"ba9102bdffe1e4a9", x"6668a4edfdcc43d3", x"fb503ffc3219d1db", x"eb1d97424b4ecc81", x"8af9fb239bbde55b", x"fd1a80f976b75f25", x"e12d6bb6fbbc7ae7");
            when 11718273 => data <= (x"0a042f2c3d1864fb", x"eec757610feda7e8", x"78817d1fe22dba21", x"2cab192dc11d6370", x"e4ea759579eec2f2", x"e139ca42d3eb9fa2", x"0cd4d88cb3fad7a9", x"1f65a03e52864077");
            when 17734679 => data <= (x"9e1f3ab29623f44d", x"c11f4fb4f76555ea", x"d832a3e4908ebe5c", x"c723dad0d17f398d", x"e905dbe02965e90c", x"3038ccfdf3c94142", x"b3e7f20184d16184", x"49654dc96ca6e6c7");
            when 17057435 => data <= (x"d8da9a4bd4bb6e52", x"2532c18d42bcd1fa", x"12679e3729c1a00b", x"c5a4b092e8a1e2de", x"45b96815dff444da", x"893a8bbb3b964dd1", x"633bc2e46fc17e70", x"5badecc6944eb649");
            when 13825761 => data <= (x"69d04f525acb428f", x"bf865ba0e82449cd", x"f0d6742b487e7545", x"52a772359178b684", x"7dea6693bf026cfe", x"d54a2f263c36ee5f", x"17fcddedb4643949", x"8f43f1195508e0bf");
            when 4739461 => data <= (x"4278f8ad8f52ea14", x"813a625c6db15d5e", x"e1883ea00990f091", x"e620a5b3117789b4", x"f9868720c1d74d97", x"76dd11db0ec8f09f", x"59cb5996d6fca49f", x"54181466831bf0e9");
            when 15036644 => data <= (x"826cf24864471896", x"8117372a359ecdb4", x"1904d99369ec9167", x"0c8fa72181544dbe", x"ad7c8554117cbc74", x"69cd2d0b79bbc552", x"1fa2eaa9c1950869", x"cc7468e5de588c00");
            when 2345938 => data <= (x"0fd42f62eb76303a", x"1dca5df16c70a2d8", x"486c4ce67b87b45e", x"999c32d1163d5ed3", x"6fe143353cba36ac", x"639d338513b56f3b", x"d960437c1806fa71", x"77c3a2978e13f525");
            when 1762006 => data <= (x"e93f9ccf2a647fc9", x"96c3167916c247e2", x"c6614dc38e5686b8", x"01ea23028708609d", x"4954395514008a43", x"a7c18f9e3f61937a", x"d96dc555877487ec", x"f192623b784f0b4a");
            when 17642072 => data <= (x"6daefc7923bbe57a", x"6fb9656d9da56aab", x"229daf514d613586", x"0763231f50f771eb", x"cba3ae25d7c695ca", x"474c9600764e0354", x"d43baf961dc80ede", x"c228120ec42a267e");
            when 3419903 => data <= (x"3cf85d0206bb6894", x"24bde6961164d99a", x"77526ca347bac6ab", x"a924ccbfc904529d", x"867a010b57885d81", x"59aca5d0bf46b97c", x"7cca7ce2958abf6e", x"40eda8c226e1973c");
            when 26466864 => data <= (x"d88df6d84bdfa0bb", x"e0c419e9c3429997", x"523df442d1dd2cf4", x"19680282fb29a6a7", x"fceaa355406d71e9", x"e47061a92cab7c87", x"580b473d5c380717", x"aa9ffb09aac029a0");
            when 18537630 => data <= (x"98c6c13f5c139bf7", x"b670355caf0f8b5f", x"0c3f043a2052f9d0", x"cdd1c413779a651a", x"56ed3c306d6d8953", x"29079e0deeeaf3bd", x"fd5500bb38518db9", x"4f2c89fcac9614eb");
            when 9707321 => data <= (x"e3f83e27a6dac729", x"a5c2801a628ec997", x"f03dbd3a54ed68f6", x"e19e2b9f0cc30c64", x"c89d9aa5e35075d5", x"fa527f722d94f9a7", x"99ef7290cab02742", x"928c1d464ebffea0");
            when 15620275 => data <= (x"2ef2456de7fbd77c", x"7c6ac102dd23e410", x"e20720dec34d9f5d", x"e2624d7d9f3db3c7", x"6cf2dad4c272dbfc", x"5f2ea53722d7e3a5", x"b80670bdf6149699", x"de482b74f5a6992f");
            when 26986125 => data <= (x"6cdeb4bcbcf8853a", x"bf6bd3d0810f5959", x"898c0540815f4347", x"70111ae604827a09", x"7ce9c8eb1535016f", x"3445e97a8070614c", x"9204e754ea985a1b", x"509333d3698a7032");
            when 7540721 => data <= (x"bb00d2fe87fae2f3", x"c6d73bd1864d2811", x"5274dbd63c48f8da", x"9246efd42efe27c6", x"36c2fd85a0748124", x"fa74e912c94f5b45", x"a63cbaa029a64756", x"3792b6cd375d0e80");
            when 17780057 => data <= (x"a9d31011c3389f69", x"65c76fbdd334f8b2", x"157726aafbdc7a64", x"376d0985c219b825", x"edac9fed1c66d189", x"27d9fe5a3520c905", x"5c59d1f2ecc665ac", x"28b71abf71a43147");
            when 18724518 => data <= (x"18de2ef1aabd8ef3", x"9d6cb9c97194c97a", x"4363e6d2903efc79", x"04b7d71b21a5f261", x"c3466ead8a097313", x"6b24ead8dcb03158", x"1ac72c0c3fd13480", x"8d130d0a6e15bfee");
            when 23600674 => data <= (x"817bb24824fa9eb5", x"6dfa1be37ee35cdc", x"df2f83a08a571fff", x"3b1836ca1002c759", x"9b9625d56284d273", x"5836a4e3038b6df8", x"c912a8e1e49b53a6", x"51f11da1bb924722");
            when 25436261 => data <= (x"fbc1bd80a90c9103", x"7dcb151439c5c2e3", x"c6f11f6f3e78b380", x"f4ace526ee0e339b", x"3780db861b7b0181", x"e8016cce9a883fb1", x"0d11cec4cc8dcbbb", x"49f91f9c4e1c3656");
            when 8783948 => data <= (x"36f4b591c4dd35e6", x"5dc2522e80f7cc25", x"5418d8d74092fbe2", x"2eb3ff64fa36370d", x"15d6315664fe6fbe", x"17d77ec95a17d4d2", x"2ed31ec276728b61", x"3716e16dc4b2d8bd");
            when 27596088 => data <= (x"b6ed2b0f8a94741f", x"63732a0bface95f4", x"e7d24bdf233d5d09", x"97ffcbfa19f92eb9", x"dbed5277dce9a511", x"bbf911e5fd27c846", x"d2a1b0b4d673d86c", x"04a4d104c1f80cb6");
            when 31259388 => data <= (x"037d6b15a5c8accf", x"ca505497d97bd2e0", x"14a952897b34ea3c", x"9b7aab81e6ca08e8", x"20ff6bb92ff84e05", x"30732ffcf80c8c4d", x"10525ee481935bd6", x"6be10ccf7a5e4ea5");
            when 23319066 => data <= (x"a8a61b0163870010", x"7a45ef17491a8886", x"dc006562cda2a41e", x"7d59da5d141b6ec6", x"c5d78af8573eb199", x"9ff896a447dde5b6", x"e44c502e0340b05d", x"35a195cd7a0364f5");
            when 25956853 => data <= (x"a4dc8fa02311fdf4", x"528735cf0a233303", x"c139ea5fdae73bc1", x"44739ecf1d6b7894", x"a0ba9697c5fc1284", x"4d2a002534d00ec0", x"611e1344a53113e0", x"e52ab2db4ddd1bab");
            when 15911146 => data <= (x"c35e13df0cf0d145", x"beec2acadb2f95eb", x"6c8e7df457982943", x"22fc775a8435dc58", x"bd1a37e2256246bc", x"858bd1bd92f0f617", x"7ee3aa302e3c50a8", x"a6280d458124f701");
            when 20413777 => data <= (x"1e0a4ad0b1842459", x"5349aec582564ad7", x"59de00bca27d5132", x"e88350e86e5304dc", x"25ca15cd63ce4a4e", x"247d6a4a35c78bc8", x"71c2ea989a5ebdc8", x"bddddce8ca1d3131");
            when 11348137 => data <= (x"fa838b9f633406f9", x"6814dce0c00f96a9", x"1d4c36e36b961d8e", x"82fa5c5f8ba57f5a", x"ed42ec454eecc50e", x"f086dc48ce038f14", x"33c17ae472f1c416", x"fdaf11b2189089b9");
            when 11688108 => data <= (x"9dafff68e503450a", x"e94a216bb3b2e9b2", x"a8bdb105095d60fa", x"e0a314e991275150", x"74e2eee7001ff3c3", x"533b919567e389de", x"be31b36ae4038bb7", x"a75f95944dbd5fe2");
            when 32703076 => data <= (x"0d46e55ae5ea6bde", x"8928b2be6f045aeb", x"614ee9c0ac9f6475", x"e8ae46dc50890fac", x"ca514289aab9dda0", x"300dddef1e52096f", x"30d712a9f4da8eb7", x"5b2c3c794739d531");
            when 30435118 => data <= (x"41690a3430904953", x"403274d1bc47d816", x"94e2a7e61437bafc", x"050708cdd23e8ac8", x"e99399b066b91b88", x"7c84cde74e436ebd", x"49c7b980598b9935", x"8e36902100029e3c");
            when 32122826 => data <= (x"6ed567a108b43e7b", x"b0a289ed7cf4283e", x"f9a63143153131b2", x"78a953071f96b543", x"4355f1101bc616fc", x"200c5662a241bec5", x"4bd14e4869ed34d5", x"edef4e8402ed1d2e");
            when 15869991 => data <= (x"ed7745c7b56987e1", x"0ed73247f33e826f", x"8db63245c0e79975", x"57caa118815b467d", x"a65d45eb606f9b21", x"aa47625793d0feeb", x"b84472b303532596", x"3eb4dc01cf0d75ba");
            when 6312268 => data <= (x"b7e94f26a5dc838e", x"52a8081eb25171ae", x"3e0f48e942d472d7", x"c3f2da1b10e07aec", x"de1519fd5eb29845", x"ea3ba1950842cda2", x"24ef91fe9cc31b66", x"99197b999fc7b84c");
            when 18507889 => data <= (x"ed225d3e84d594a5", x"4975102958dc64b2", x"73b4933b10c14d67", x"9263faf9c900b249", x"143f73513ce39911", x"0c724db39acac7ef", x"c69345e36e96a004", x"d7a0c28b9c92afb2");
            when 16587371 => data <= (x"d6ac805f7fe5ec7a", x"a803af6ee10ebdb5", x"eadab3aac90c3474", x"d3676ddf8e437f4b", x"a0edbcf33f126710", x"92fb1034d0baacd2", x"47ff25f3b6fb520f", x"5007e6a6e0a387c5");
            when 1727610 => data <= (x"782027facb0cad29", x"0dc7a095d7edd8c9", x"a445e2fd6a116363", x"001aa62110aaa27b", x"4815de4815130159", x"e73c93da248bba15", x"031f9d4c8e9eb6fd", x"038642eb2e12f303");
            when 1461518 => data <= (x"d9f4f3395ded763b", x"db6106ff767ae303", x"c75b556833568e3c", x"3e3d3c7ad6196733", x"e4b750d65d88dfd1", x"eb1edf58885f484f", x"2fd7cdead878bdc4", x"b1cb83f6e0d50c60");
            when 17601030 => data <= (x"bfe4414650aa61e7", x"e98b1c3518f3d103", x"c4e40f79e568b19d", x"0333b81496a23d13", x"671c28480af735c4", x"ca3072901d40690e", x"b06b6827cf7ff810", x"776bc1614fe552bc");
            when 13240582 => data <= (x"b220a1e9dad33d61", x"53127fa626b73d25", x"40af16a5cd4053c3", x"f3c7ee50115ff13e", x"ac58dfffe07e1948", x"f942d67dad915a65", x"589f81ebb551fe7d", x"a7c510eb494c3dc9");
            when 3934710 => data <= (x"225ed58d9a2011f6", x"038cd3d524fdac04", x"d499b520c8232b4d", x"3bbfd437dfb23b7f", x"80400aee9fdaf651", x"172376fe45aabc7d", x"97e0db3fff3c5ff3", x"2397137cf4b2cb19");
            when 15003034 => data <= (x"8dc08d40e7bf3e67", x"c3661cd9157e95c7", x"53e25cfdfc113159", x"29b2173ba78fff52", x"e8ce3c5f7264fc62", x"a5c2257f71983384", x"202d6d94d1bbcaa8", x"e1f5c7f3fe5ff165");
            when 18690390 => data <= (x"9534691fe89c9fea", x"41886284e6d01197", x"be2a9ff181e6a256", x"05f1ab10222b8cef", x"92530b359f3d2824", x"471eb5331c5d6d02", x"f2d6beaf5f97134f", x"0c0e59516f1142c0");
            when 15816810 => data <= (x"a3d1d8aa7f25521f", x"4bf4e3e553cf0321", x"f7a5ccd61421ca0a", x"02c3a1994cd2f3db", x"9b1a40a0712e923e", x"d86600ee3eb53613", x"2812fbdebd9a1522", x"67163dbbe7af2ae0");
            when 31750214 => data <= (x"5d33fb416f4ded71", x"400bcd8ad6e3c8ab", x"d0726856cf79948a", x"9582382ac857d66e", x"565565ea47a4e079", x"3e284ca180506ef8", x"6a1f1ca172df7f2a", x"955d36ce384484cd");
            when 8904218 => data <= (x"ad8ca68ca4a860dc", x"dc6a5d5665d1f36f", x"0a9e326b3de5cb3c", x"ab0ec83ca8d45ce1", x"391d43ea90a90899", x"555927b8a487453d", x"146562d90e14edab", x"31389f7a533ab715");
            when 13407684 => data <= (x"fdbe9b335cb5b976", x"8e16bbb7e79ad1dd", x"08b75732b99486fe", x"e629c174b28f8f02", x"f17e19b4fc403f35", x"0c6a9d485c05911d", x"93ffd611bcfa92e8", x"988e67b6f52a36e6");
            when 11467249 => data <= (x"72846444cf3394d4", x"5c0763c0e92fa874", x"6b71cec2f33f427e", x"25bcf35daf8d44ba", x"a4930238201a092a", x"f87935e1e3cc35d8", x"efaac22e9119c0bb", x"01e99709cd4e1eaf");
            when 23504983 => data <= (x"e7c9d572a2d7bdb5", x"f60671c64e732c64", x"44b20f50c573d8f3", x"1002c22f49543266", x"bdcc234e21385238", x"e1cdf644457ec2e3", x"adb1fc86dc9b1aab", x"00d471760ff20376");
            when 2070307 => data <= (x"1c48215008e1fccc", x"ca997902895c7ceb", x"f53cf8dcdbae5e3b", x"478eff3296365db3", x"fe4a92a77a564b04", x"0992e8fa95e09c34", x"6585faf3b26d5f81", x"2941b75deb4b1be6");
            when 7907561 => data <= (x"d912aaca5b6fa1ee", x"95ef9d05534b3599", x"d21bf671108d8afb", x"ada00553666792ab", x"7b578415232e2122", x"9b9fc1393ef8bde7", x"a1dee9a452827596", x"6e5b2758c65e3508");
            when 23816390 => data <= (x"9feb9ff2911adcdc", x"0f4d32a2337d860a", x"b774e2b2084ddeda", x"bec6f3c5aeb7e12b", x"1b0c609a758f2eac", x"08ab84b0b9eccc00", x"e8953c00a85b62c9", x"5a7b19062257809b");
            when 18925491 => data <= (x"22458cb785be9dd5", x"febca78f7579b6c2", x"a1bd80cd2b1e0843", x"33e2016de9c79368", x"5ad2e3d70afc42af", x"25f4f6507d908baa", x"7ae4d77e6ae5d7d7", x"5f92d32eb4331743");
            when 23301247 => data <= (x"18f076b1bb15ccc9", x"372be7a0ad3132b9", x"3d26cf7bdcc2d277", x"881ab80823cfbfb3", x"f3f161f3da7f86f7", x"fcca8b94aaa928ef", x"a3f487be7289240d", x"5c058afe4ee30407");
            when 7902665 => data <= (x"325cf8a531781b5b", x"e78e9ab470a07d89", x"22b3156ecb40d337", x"813821318a3b8e22", x"3d19d4ea4b2772ae", x"c16ae5ea4782ad25", x"f3b0cd3c668ef3b9", x"8c6ed921447717fe");
            when 5122967 => data <= (x"aa79489de30b5d77", x"b10f97fe0e0b3ab5", x"59e23408de35b7ea", x"17afa6799a58db50", x"36a40014ee8bf4dc", x"be7d4946fbf66436", x"c074e21869934e6a", x"edb6583a094de699");
            when 29718963 => data <= (x"8017aca2ea032143", x"97dcb9929ab13aae", x"e5af35d4c83f9cdf", x"66151c11efbdc822", x"73df74d667078f8d", x"c1297b7d8d71aa8d", x"89eef0ad9a56ae5f", x"7361b3e098966fc0");
            when 4004393 => data <= (x"bcc1032e2379c365", x"7e3b9872694ede02", x"2dd264ae054b0c3d", x"903017663d38bcee", x"dcf64ee542e72902", x"17a13bf660cc5110", x"61796b3c99a71a76", x"7e6800bcb131dbe0");
            when 12849909 => data <= (x"60ac28c0e0568f14", x"5c4ea69b484013e5", x"d41dfc391fcf2382", x"5617361332838a6e", x"81328d0411706f0b", x"9cfda0a0715fb04f", x"55435f09a70d6ccc", x"4ac0171355a1b777");
            when 19199497 => data <= (x"84b15efb49404acc", x"4435844e7f860196", x"90d4eb531748d5f3", x"7c8564d68937fac8", x"c18c0d4fa4c47969", x"9bae11a4bb593215", x"62a22e3e7022f3a0", x"c04c652ff2adc668");
            when 8227129 => data <= (x"3fc54744c8089680", x"fc8f61177449d2c7", x"8ca21000bab81dc6", x"70b2b8904acd813a", x"76ae8fc02044e257", x"d00eb49f8a72fa9e", x"3ca82814c810f91e", x"8a3e1139de307572");
            when 3696764 => data <= (x"e093634d1d1ac2af", x"1f4c457db07ecbfd", x"cc9952d05a519e0c", x"b6e29eff348d93a2", x"e35d5d1b933d4790", x"02b651dec2f1deff", x"fc46e6d7f4815690", x"ee2723959a55ac3e");
            when 2364254 => data <= (x"e4c78ee8310231e9", x"76740444ccaf2946", x"78c22ae120ed9cb7", x"79de0223dfa65816", x"b9c36ed99f2fa0d8", x"0a72bd17b9b3f04f", x"a53fc987b95d70f4", x"35c784f18a787d00");
            when 27127596 => data <= (x"7ebd462c6130325a", x"6c6329cbb974057d", x"f7c144b25e460d8e", x"486e660d7206efdb", x"6d318c70b1f1d5cf", x"cd8c43292361323c", x"1974bf6cff0006a7", x"4a3c8b143da53c04");
            when 3009371 => data <= (x"70330d9b6a195904", x"51a5f9f3da1e3520", x"5defcb2a31007588", x"5b36928ba46af79c", x"6656e13b8dd0102b", x"860203b2baaabac2", x"8a71c697478d5ac6", x"310194a6a6bc8069");
            when 803140 => data <= (x"b93267faa8c8b69d", x"d67771be36bd36a4", x"ee06f6e41e074baa", x"385f67e63fc70d6c", x"c18a913201237b13", x"366de35924b3e521", x"720cc6133fa45b16", x"7774b3b89a994ebd");
            when 16015372 => data <= (x"0d72b149cebc5e3b", x"a78e15e828deae2c", x"15e895d85ba2bd19", x"175c822091525978", x"683a4cae3347db75", x"aba6446c673eefba", x"a926a8631b13088b", x"6eca94c277134fbd");
            when 8819075 => data <= (x"cdcb7db93bc1b0e1", x"a1c4b25621d72735", x"ca8f6d758ea3bf97", x"b891add6bf3a4985", x"8222de9f92712971", x"de6476d1b553f8d3", x"d233a4d4b4b9cc73", x"8f1dc77545c745a8");
            when 17186940 => data <= (x"9b09e79d90de9e37", x"d0d615a0d0c6055e", x"4eb9a82cee9090ce", x"4bc095a8d4cb9a1b", x"27bb4a4099675cea", x"81d305c38f431c91", x"383527f52dab66e9", x"d9c0579f4382c753");
            when 24323240 => data <= (x"eaf8b22f1ada33c4", x"fcb92ccba68e4a28", x"7026cc2fccd9f791", x"c2e25d44e2b7770a", x"46f4cf0379d788f6", x"9d2dae71ba3fdb3c", x"bf439d3c357fe0cc", x"792070c6e7ea0dfe");
            when 32933559 => data <= (x"ddfdf374c158a105", x"a317020ccf1fe94a", x"df3b774876341f9b", x"e0ac050d968222b6", x"d3201f95a27d52c3", x"5088a3f4603a75a1", x"364f9c2f997685c8", x"0cf6f34025d6fcd5");
            when 16655854 => data <= (x"215f41ca755b54e7", x"66a9ac34b99452bc", x"92d23e90b849f87a", x"58e3e34693cf194a", x"e5aa6df33104d5bf", x"17bf6f8b4ec419c7", x"70553334e645ac0f", x"d7584e9992e1eeff");
            when 22895077 => data <= (x"c33635801bc0b7d3", x"dd0f3e8c98235726", x"b3ac24d2e0b3b1cb", x"27d7d91e02773627", x"5bfc02164245ca63", x"0c7a42188e88ee59", x"e4419b9841e3f47e", x"541d4c7206bdcc88");
            when 31958102 => data <= (x"7dacdc84ba30b9f5", x"36508cbd84915b22", x"aaae37e3cf93568c", x"a0134e031f275a59", x"440a900ae507b7b3", x"34628240755f0ae7", x"e266735df9f9446a", x"06b1ba8bdb65718e");
            when 13461657 => data <= (x"c11a6e77560f2fe6", x"79bb03baf0ecbbe7", x"99e8a44714d866fb", x"642cfbeef12aa54e", x"a5ad6eaac346e8ec", x"c2230619ffb070a8", x"2bd10bbdd44f0ec5", x"57bb826a7c216b8a");
            when 627646 => data <= (x"0310835484332299", x"d7b4bb14faba5d5b", x"87ce15b1f10a0415", x"291806405202ef57", x"b669f9239e028285", x"30b696e91092c656", x"f8a2eba22e9ed04a", x"3feac2aeff93add5");
            when 24780069 => data <= (x"3d75773f92433912", x"cabea511892875bc", x"d263b130d94727d1", x"c29da06fc7a870da", x"6b946c428b388122", x"e7849c12777c4ba1", x"d2fa2debe3325b26", x"df97bd5e3ccb359c");
            when 9674792 => data <= (x"c87af5456f53c7dc", x"a3787ef1d7b49640", x"31f21f7a072ed39a", x"791236c673376f32", x"cea2332519060e8c", x"56a3d6449d34b848", x"10262ddc00e02762", x"492f43dafe2f6eba");
            when 32695393 => data <= (x"82056121aedb5bee", x"6c2cb805966c304b", x"13c77dffee300d1f", x"a345dafc4c964e3b", x"c61152ed3d3e6912", x"19f7ee80b0d2b53d", x"2fcd0ae5d5ed3581", x"5b7f2672b9072391");
            when 32406013 => data <= (x"0522716723617702", x"900e3fe3a6ff140e", x"aa6f717ccbca18fe", x"d91eb637e55d3ee1", x"7bde2807e5d05bc5", x"6b442d92d45f423d", x"3dc54726e7bfdf5c", x"eae9abef21ad5b68");
            when 17901421 => data <= (x"c46a9fff76cf9c2d", x"d34a1cf666a19ac5", x"626a35d63735c94e", x"1d7c821974d5dbac", x"50ede9dd715e99ae", x"e5cb1e97b97b3bc0", x"57c0db012110a9f4", x"9c11972939391e52");
            when 32739991 => data <= (x"6bdd3ba3268c336c", x"ba24c48f6fcd93a6", x"816ea210c056bb91", x"7eadc08f99ed6302", x"f6c66e3a643f6247", x"b6d000b23ccd1df3", x"0e16ac0d63e78e91", x"090a1c09913501db");
            when 12018534 => data <= (x"ffa75e17793b0963", x"914ca905eb117f07", x"6780f8e17f7ca301", x"281d8fa47d7367de", x"0ed8de171bb1584c", x"a568b089dfb10709", x"62977318a0b0ceae", x"eea3f2f88d1ca014");
            when 27922667 => data <= (x"714b135663ee0c6e", x"bdb621e6e57f3624", x"7c1f153723d40265", x"850564951c901aae", x"a8307c58f407f301", x"8230ebd7523417cb", x"4942c2859d782691", x"28d12b415b81f1a4");
            when 25378288 => data <= (x"1ac204118dc67ab1", x"d9c6253f8c22caa9", x"91f81ea484c6f3a2", x"e209d677b0686783", x"fbc3b0783eb9fa58", x"53ff07f4b46399b9", x"84d0b8764de166d3", x"c2b0f8c2fcdef99c");
            when 14578841 => data <= (x"b026a4d5a319b0b5", x"1c8f391d22ba9a10", x"eff7adb276b770a5", x"7248a2d052dbd9a5", x"1315650dd4d7e33b", x"7dc36128a0c65483", x"4525f85d38330f3a", x"9d11529ab7da907e");
            when 18147835 => data <= (x"ca0ac8a274644180", x"3eedb8f4ac1e7768", x"fd4e331c5e67d6a3", x"f5b88860f954beaa", x"6c95e2f267431a1a", x"c897b652ef4ffd2a", x"581605c6b611d5e2", x"c39314b0ad14e190");
            when 8556752 => data <= (x"ceea288f105d85b2", x"c1127095b1c73d32", x"3c3d3729424d2153", x"9c2b0a9d02ea6f24", x"61d7f1887e521834", x"1b87fd317c458859", x"4d86f7092bf1ba96", x"8d493e34f27f6d59");
            when 24308033 => data <= (x"a197d8c506a36674", x"4f594397fa111694", x"2a16ee370eeff018", x"351a31dcf495b2ee", x"103a4ad9ad915859", x"07c8026cba3c8a43", x"f95d880c9d4147d3", x"e9c22dbeabe11060");
            when 27447611 => data <= (x"e84fbb85f22f2e85", x"0de91aae11a456e6", x"6ac973c442790914", x"c75675a866bf75de", x"bf3ff5a53fa9a314", x"ef1ee463fe206aa8", x"7773548aeee8bd99", x"86af672dec8ce0d3");
            when 21495530 => data <= (x"587fede369d7876b", x"fb331b5af7ab285d", x"8711a56503a23fd3", x"d5ec54f287c8b143", x"8586e10f8dcc4b9c", x"5af48f010b0b192e", x"41908457b4069e88", x"c6c1695d00873c73");
            when 32557494 => data <= (x"a0f6de326438ce73", x"ba77a3831ac836d6", x"54839a6600284750", x"a07262ce32c73530", x"19da8cf298d7df7a", x"90bbb0a5778e1dd9", x"0abae92775072549", x"6da3e55ba3296e27");
            when 2734601 => data <= (x"693b573042ed39bb", x"273871f99c344272", x"238b09fd61e92796", x"716ccf6ec8c22029", x"476e0df2bd55bbb7", x"15afed2714218924", x"6505cb7b51a2de7d", x"5cfd7f1ba6cbb81f");
            when 7895400 => data <= (x"9a35e5355e5afd38", x"831830f6da0e03e5", x"fcda7460ff93b162", x"5c31bc98a1b3458f", x"05b101bc59a79959", x"e61ee2fddada3704", x"6c09184524876f0d", x"1dea17edb455bc2b");
            when 29145154 => data <= (x"af73a271ab6c08d5", x"59eac68f2b1ea0cb", x"b3384dd8ee569c66", x"9dba916525c38f8f", x"998b2f9d75469d49", x"d3b1f5d7719cc49a", x"07a65534059ff813", x"3875830c26747399");
            when 5714195 => data <= (x"d70753e30ff994b7", x"2157607c03fcb558", x"01ceb4fd92b500db", x"21ccac204ed03f78", x"2ab0c8c02b482fc0", x"3fd6d153226a0c16", x"32bd6a4b495f6fce", x"2168645f3dd134b3");
            when 13536167 => data <= (x"018dcc92c5dafd27", x"f2ee5887e37a9ccc", x"29bd411d01148a6f", x"81f1c7c6ff57ae5f", x"55227cc5b10838b7", x"90b6f8adb420caab", x"13ada74dace5e1df", x"ef5274381481eb94");
            when 14750175 => data <= (x"0714314198bda65c", x"7d205a90b181f682", x"204e2f6f033e3d09", x"310729a515e38a1c", x"f3eead6dbcf19a32", x"53d3f9a74dc9b50b", x"aefa913e5e7a8f51", x"d7dffa93462b68c9");
            when 8036674 => data <= (x"278597fd7882c58c", x"e951c855a26e95de", x"564e61f0a3f136fb", x"f74d0cd79cce4458", x"eeea14ef23ab6fb8", x"6ed78c6fd77b6d5c", x"f94cf12644c25777", x"620237acda3d048f");
            when 28393984 => data <= (x"15272db79c0b3069", x"a4e3fa40d2fafe86", x"36c4ca10d0b927a8", x"0988f98541bd2de2", x"6c3155b4f7a80565", x"6000bb64adb58a44", x"bd9c7fa3575dcac7", x"3572aec94da33bf0");
            when 29946049 => data <= (x"fc5ebc2fbf51cf60", x"b2eb487912557588", x"b8d6e2153810a133", x"bf9ab5b742935c4c", x"1c1e4947bd172e21", x"ef72a67c57dc9d21", x"477030bf4a01dae5", x"5de7c910647281dc");
            when 10866910 => data <= (x"b91270f07b2bee29", x"e13dd367529b0bfd", x"fda434bc97ac8a1a", x"cd39f8cfd6091519", x"12893c38835dbc67", x"af9e992c602f2b69", x"eaa1f5e7bc3c4328", x"0b0ec026b5c415d0");
            when 7639053 => data <= (x"fff607bf58750d58", x"4438a6afb05ca54f", x"5732e62d703ed07c", x"888e4e60936b9dd3", x"dfc57a25972bdaf7", x"505a62c2fe6d717f", x"538371402bd5b5c2", x"52146d44f5796aaf");
            when 14213931 => data <= (x"0bc5bd99df00e07c", x"3a4a882b93b3e62e", x"92c89e89ead3537e", x"a54b8c1fe8e74c85", x"dae4bdd69d5c1d69", x"ef8c77b442c3c45c", x"2a6b941275dd3b80", x"d69edb332510d240");
            when 10616220 => data <= (x"f6368545ea15aa45", x"9aa8420baadd704a", x"92c39d573cf38cba", x"5cffea002731ae0e", x"b3151c80177fe7c8", x"7a4689c23252f10a", x"0e2fc806d55f46fd", x"a936b5cf87b0bcbe");
            when 16601558 => data <= (x"4fca26faa21812a1", x"ab139034e8b27309", x"67b9e302907e664f", x"fc409d09dfeaa4b2", x"88a9bfd6f84333fa", x"b5fb352de7b81488", x"841293e05c75531e", x"6384565fb68e24ef");
            when 29035039 => data <= (x"a4673beb558f819d", x"a710362bcbdf1011", x"d5ae92c5fb4be513", x"deccdad3849ffc43", x"10d92f87c5caf083", x"d1ccd99095007c98", x"a42f771299f0089b", x"e45ee8020d771a2a");
            when 14890724 => data <= (x"d6eaa610db757e80", x"ddd15361a9e7bf62", x"1a68c3b99253403a", x"a6a79d64dcf5b380", x"a4d607a1d0b83f71", x"03f5548302236fcc", x"37f491d64d1fc975", x"5753465299d49cf2");
            when 25363508 => data <= (x"65453e580953792c", x"3d8c7f00f4c2023d", x"f87e0aee2387493f", x"56845b74a10cb25e", x"95c5dcef6bb3342e", x"5e1fe9ea99f3df93", x"b99e725a042cf727", x"aad44311099dd5a0");
            when 23426066 => data <= (x"424a919cee910d1c", x"484018ad2addf064", x"c75d2bfee5dab81d", x"348db6719f8ba9ca", x"f9a5fcbf1ae5b81c", x"355c26485ae26db7", x"254f5e7d5689f2d6", x"78264a37d004711a");
            when 16390999 => data <= (x"05450d6aa835043f", x"bf904982ceb7b897", x"e9809176984b3ed0", x"ef5b02afceff1ac1", x"df9dca80de92119b", x"33f272a9192d3c3a", x"125bd91335a74ca6", x"4560a22a993f1886");
            when 32408654 => data <= (x"720ee3cbc74d12bb", x"de80265ff04ff06c", x"ff198beb4bddf6cf", x"8cfe990ab84f9618", x"ed8aaf94b42f947a", x"ab164185bc5434d0", x"7b5348d8007eb9ae", x"d9b5f194246937a8");
            when 5436763 => data <= (x"d03a73894b216acc", x"a1bc88e5e4860c53", x"ac75f23ad6a45447", x"e155dd20c356fa2c", x"230f03f50a422057", x"66e29817c40963cb", x"71b1118726cc91c3", x"1402a1078ad7256c");
            when 1972747 => data <= (x"f5d03c151e82bbdb", x"cf21a816c0fb197c", x"e045761e14a56b5d", x"484623c233f82252", x"a27f09a53bb133e1", x"32f7e4f008a3abc9", x"57643bbb222bcbbd", x"05426bb2a0636e37");
            when 4465594 => data <= (x"f35042ee49da0d89", x"0d3986df18a20597", x"d54d88437fd6b097", x"eca38c33ecb91210", x"8bfe6587124328ed", x"da96d196ef051df1", x"bafc6493d54b8acc", x"f2bd160182107128");
            when 31146957 => data <= (x"e91d113c9fcce97d", x"9d6e1572d724f5ba", x"715d686fc8704296", x"3da497a2869998e3", x"8b8d0c708b21c394", x"d2d3755824024ab3", x"779119a732285546", x"25666ebdcc191f51");
            when 7864900 => data <= (x"ffb6bce6ac48558f", x"d4a75f7ba3c8e29d", x"85ba1e5d2fc3080f", x"cd89148dbc657554", x"ce27ba529ffe2370", x"d05c246cfd32afff", x"52a39d78946a1079", x"aa900b683d8a170a");
            when 16084946 => data <= (x"4214b19843dd2100", x"857ee082c2ef58f9", x"68f919318478bed3", x"1a530a06308839f2", x"f683902ac807247f", x"52f86d8973370066", x"7bc929ae2b735b19", x"7366965177e10d0f");
            when 12910107 => data <= (x"2f7f764755879e2b", x"0330e7688eb79f7b", x"5b2b2b3312c4dcf8", x"24466a42446b800e", x"b9b4fd671be40cfa", x"c4c840802c3218e3", x"4455e51067570f27", x"7092db5a44ae6d87");
            when 5438354 => data <= (x"16d31c0442c9362f", x"e0c1ee8348fec191", x"9cc3747eaa45f2c0", x"b476a97511e57d3b", x"de946842c4daa457", x"5bd79a5aee37ff9a", x"e83d4f4095bb5fdf", x"a2a45bac18fe87ae");
            when 30304066 => data <= (x"aab0532ebf8b5f7b", x"fb18f13b6d230ae7", x"473e826856ef2f0e", x"9b0dc6ea5e4c21b4", x"3b477b65c5131d41", x"d3968751a59d1cae", x"be64ecd73d3776d4", x"9dbe1c89041e2a18");
            when 18631688 => data <= (x"21fd622554de049c", x"3aab26a3df02ea5c", x"e60a83ac98f69081", x"332834d3134d39a1", x"a2e56ae51c778c54", x"0bcb89b0cc02e82b", x"4deff8ebf88ebfa0", x"725f4790f491c4c7");
            when 32322313 => data <= (x"87b653739325573d", x"0852a42e175afe13", x"9e0e0e18b72e10c7", x"0ee6b59a33204915", x"00ebbe023997c349", x"14b7eb9df61776ea", x"59ca546360b7ed40", x"a28d18699522e6f3");
            when 28202822 => data <= (x"c68d4499750f8e5e", x"452726c83879de34", x"d382c93500cdaa27", x"7743b0ec7984bdf6", x"78b0b24c26df19ee", x"55801bee08165894", x"35903f20ba95190a", x"5938460082eb4344");
            when 25179064 => data <= (x"e8c78a2b4ff45b2e", x"e9842afc3dc06343", x"d25f98c6168feeb8", x"9963b7e7bf17027e", x"957e2dc8d0c2adeb", x"8c27207913605b7b", x"7e6aed92faa9e197", x"9b07656f49ad6780");
            when 10836267 => data <= (x"4fdf58d5e88a4122", x"009d12ff9f80c608", x"63b86e678f7e7f97", x"5966f9c2246839f1", x"fc1c1f1b414101c1", x"59c66b5abb5f85ea", x"d4295d47d8a6b7e4", x"4b732b397a27dc15");
            when 8362822 => data <= (x"f3a6af7f0cd7f006", x"236bfe88f8e13e79", x"d48dc91f5ee759d3", x"1d9635f3b6f305e5", x"e77c605c4e17ba52", x"f3299c6f72255186", x"fbdda17ee29374cd", x"b57e513b115ec64a");
            when 32129611 => data <= (x"3e10ac17a0667dc3", x"b2ae86cd79a2c558", x"e2c3408e16307eac", x"c81fcf3e02732351", x"84b9aa35c8590f26", x"b9c39b81d0476ac9", x"7dcad49b4374a75c", x"2a9f20d1481e9372");
            when 7295372 => data <= (x"31ebe91485af80f5", x"75fa20efdf0523d6", x"daed48947b10dcd4", x"10dc223b99e905f5", x"5fb210b5070832e8", x"c4ac8a623219f59b", x"5f33f0b36fe7e42a", x"0dbafee78a0c6923");
            when 21684055 => data <= (x"0ae72224009c2c1f", x"11b29f180f250f2d", x"733bd3e8675aaf3b", x"18ed503b5f301dcb", x"8398602459ffe1fc", x"c26de50f2faf10c6", x"c1e510f25589c6bf", x"c7151fa6b5a8b2c4");
            when 19490104 => data <= (x"121b584c483ca953", x"538f0a2031a22eca", x"298775c514da8199", x"51ec53ae8cd8ed4b", x"dbef0925af6d507f", x"7be5a8aeade5b998", x"547f88411f8068d7", x"6b70f90e1ba3a9f5");
            when 7101323 => data <= (x"bdfd9ed27c1003c1", x"c1636c1a554fa03e", x"a01619580f207835", x"764d209fa134d11c", x"32cd5744525222dc", x"af74f9e079e7e5a9", x"fc686a2816493a8d", x"9d9bb3b69c065d8f");
            when 12929911 => data <= (x"a9bf0061f6c4f683", x"98176271b2f5d1a0", x"8ac9e77f3d2f1095", x"9d04cb0078cef8f8", x"75cdf36a90141133", x"220a3240d61d1d82", x"c5073ab815ba5e19", x"aeafaeec15e372a4");
            when 15494022 => data <= (x"8d2b3ad645c04952", x"40b393d1b6b9a812", x"ef966ca7e1749dc9", x"f50fd1a108921e45", x"228deb0e37f092f9", x"1316678428921e8d", x"f15dcebfaa48577d", x"93f9f4d5efb6c637");
            when 15718593 => data <= (x"ee9f661b1dbc92bd", x"68b7288def6913e9", x"2f8d22aea5e95c4e", x"bd360892096fa4b7", x"e2f0b2e61d8d81ae", x"d2dc01e26c963d7f", x"1e2969a03f9459fa", x"6edfdfc656e4cdcc");
            when 33698247 => data <= (x"7b6c56079727639c", x"af79b6393473b8fc", x"5a7b331166db477e", x"25205e225cb0295d", x"f32f573bd5d65dc4", x"6d5815703089c13f", x"01cce753d0064f01", x"cc0e40fe59bfec59");
            when 32228423 => data <= (x"07b5c691ae6deb0b", x"14185aee29b52eef", x"96e4b597ddb8774c", x"968aa5bd037daeb9", x"030e2e615228ab81", x"550766feddfd36f0", x"170e19d4f65ab302", x"06c8a3bf6af9eaf3");
            when 4368187 => data <= (x"4ac6dfe3af3134a6", x"c9f67b81e5210bf9", x"706d9df3b3863d32", x"14b5e8210e38411e", x"b4a75d2a0c17e70a", x"e0860659fccfe8a6", x"a28771029a5fc75f", x"9b7c96c13b3e24ef");
            when 20050699 => data <= (x"2660f02cb89c9c2e", x"cc81247ab159bea0", x"e08de3f1b84395be", x"34d6d4160e1c4bc4", x"0136c10abb8862f6", x"c7acc66c125a4c43", x"5f5195d832b6c5d5", x"7e881a2476798ff8");
            when 9871020 => data <= (x"e620d486ec46d3a2", x"378b03d85e4c57ce", x"6b3c2dba3d653e02", x"fb56ffb2c2d73d47", x"7ba75caccee2a390", x"9ad49db5554554ac", x"b74ffbda4134fa3d", x"1411a7e30b210675");
            when 22903571 => data <= (x"6e4a0a7245eed631", x"62a0040e9f91621f", x"7227ec99c9d33e0b", x"1a536c4430b7c2fc", x"66a18da12467986f", x"dd9a40a89b49eae0", x"1a11bd64fd465e7b", x"6940af9526f4e6b3");
            when 29128196 => data <= (x"077b264ef17b71d5", x"c1c3c941b583c475", x"6e5ab06aaa04ca36", x"a86671a739633801", x"82bb34f552332a75", x"14b0c6d260773a67", x"eb92d026aa4a0896", x"09a63630284cff25");
            when 3304343 => data <= (x"69c9f1126e042ad7", x"91ca5750e12bf087", x"2ceb44abfb8660d4", x"5b16833b2e639140", x"21dc8032af3a82e5", x"1759c8403b29ba13", x"2a81cf9d0a77bcd2", x"a7840e85525d5225");
            when 23951206 => data <= (x"273ce3497911937b", x"0515c8e456f271c7", x"a14361aea0434c13", x"a5032175afd59595", x"98c954c4a104d279", x"db005e04a1a43b6b", x"0dbc0e56036874b7", x"4ec25fd330d8c152");
            when 2390125 => data <= (x"f058a7cda94e949b", x"1aa2a22dcce13bf9", x"4b7d837367b18457", x"2d1f30581d6b8cf6", x"e7c566d129f55830", x"0f4ceba4c76c7416", x"2f46dc6f1f54c6d9", x"aee321759b709179");
            when 13024770 => data <= (x"9c9e0448ab3ab987", x"06df4fed2e3cc7e0", x"e6ba072756425236", x"106f4ae3b2f88bf4", x"1f0de9c4a8ac8af7", x"1a57306a9b21c1ea", x"1fd19f4a3f187ad0", x"8d041cd777ff11b2");
            when 12102478 => data <= (x"0ed1634b3dcf3cf8", x"f9f8a0feeba1a0d1", x"848d49f4950736a9", x"d6328d3b53d7d5d4", x"4f19dae7784ca3d8", x"25e3bb5354328193", x"27fe5095544b7056", x"da3ac42847c0d7b6");
            when 8623076 => data <= (x"5e4b4b692ba5c9f8", x"e127651b0afd4dbb", x"70136137effd4c6d", x"445aafab75f4032d", x"1995e04fefb33bdf", x"94cbb836054fb978", x"25d5b87a847fe765", x"cb1dbedd48e1f6f7");
            when 21865054 => data <= (x"a5101ee05eb68d31", x"7f25d2151469d7d6", x"2c204ac70fae7f59", x"666713e99a2b198c", x"ca3d976ceaa19b54", x"deab91587711020c", x"2b695a5ced29616d", x"e1815267e7771ee6");
            when 3943010 => data <= (x"2225e05146c274fc", x"c5d1f54759623524", x"3f0f1f038a7ab52d", x"bd395fb9a3f184dc", x"2a3e49f3b89018d7", x"13bb94a1943a4969", x"80984730e94bab9b", x"2f3b69a25aeb71aa");
            when 17340227 => data <= (x"11f09f2af1adc798", x"4e716cd660b5ef51", x"1992ab0c898a49f1", x"3101c6c1e506c1ea", x"97e565ad16b8a071", x"b99e4e82e43ead99", x"17f192c46a33c856", x"002b11d2a2505034");
            when 12777261 => data <= (x"a1f6d087502ff52e", x"ef926e16c56ca938", x"8ee3d9f32b60d5b5", x"9d5c37d269b6ccc4", x"433a6296c14f19e8", x"585960f53db25c32", x"2dc1d1b7c3f62076", x"2086acf2bc02c6fa");
            when 21066173 => data <= (x"3d41405ae6ccaac0", x"0396cfb95d0c6c57", x"ab347932454e36a7", x"b7b1aac2a99ee50c", x"d0c469f8957ec0ef", x"6635ab5d55af6cb4", x"4c438025b34eb35e", x"bae96c5d5b9ef6e3");
            when 17139771 => data <= (x"740ece5f5cc76102", x"44bd5a01eb447861", x"e2feb2f922101cea", x"27f21f2bc5243e88", x"40a2984c8225d9bd", x"2c806bfaf4e7449b", x"5e6ab6e029ebd29e", x"e92bf5270dc1491f");
            when 2020868 => data <= (x"822816ad8384e553", x"bd9995bd94de88d4", x"0b8b18c0b6d1f4db", x"09aeb940e3e8d19e", x"fb72c1a8c33791e4", x"8b596a779a258019", x"2e1935ba27411923", x"7313aece063c0371");
            when 7527053 => data <= (x"5e3812d23da6efcb", x"da010f36475356bc", x"138df98a16e0925f", x"823bc1350008d346", x"ee633f04cadbc65b", x"80ccd99e32f31573", x"21b5a020439aa315", x"baa30004c7fc716a");
            when 32206972 => data <= (x"2abf0831f68b5aa3", x"25e368d74fc65a28", x"6c9319db929fe2c6", x"b4bc8b9a0af12b6f", x"a81c716c0f6c4a90", x"89f893fc8ab2a59a", x"0052b94c1ce83ef6", x"29c68669b340d8ab");
            when 17397962 => data <= (x"1d7f632bfa7119b7", x"d7813d567f2f03b6", x"02ebbb929136ba14", x"53fe7d5f5537e5a9", x"f31ecdc051cfef9d", x"59980f864a0391c6", x"aba78f6f2d23455d", x"622315207d1cc6e1");
            when 26642437 => data <= (x"fe191cb68217f967", x"d924e7d85271f725", x"55165d3506953d99", x"ed8c3496fd86913c", x"5013229bdc8e5143", x"c1b8da3bbbc524db", x"029c88a82789b44e", x"06d0b357573fbf34");
            when 21861963 => data <= (x"8f4db8d23247beed", x"228991f63d170b13", x"44bb6467d22c55d6", x"010b637ccf70bf9b", x"8bbae0e512455a84", x"30b53816fc716061", x"da7ee2c37f63d952", x"24e0294013620898");
            when 1116337 => data <= (x"cc4d3d13c549a133", x"7dd847e9bb60137d", x"a48359246a0704aa", x"64b4732a202e03b4", x"317e016b49b67138", x"5a61f661a3a563ba", x"c4f13e65762b9c30", x"844da4d1f6e370e8");
            when 22637073 => data <= (x"98238b498e7156b8", x"85b605038da8059a", x"f591cc792add5ba0", x"4c9eaa4c601459aa", x"d8fa7fd0dcac5d3c", x"3ecaeee9149e9858", x"d0d627158ed66a70", x"f30562128d2b5813");
            when 27904269 => data <= (x"8f453c9446601826", x"15c9c92eede52cb6", x"9f8ba89f145d40c8", x"c5515e5964b3ad52", x"551a617c05265012", x"07680b301df7d1b1", x"fffe7271eabeebc2", x"faa13aebc97e3642");
            when 13346033 => data <= (x"769eead3e572d40f", x"7ad140ad962123cb", x"69ec409e205a16f3", x"77c30cbacd46b68d", x"3a6b43ee5ab3393d", x"b523ebe5af09f555", x"d6cad07f27b4c2e5", x"161f6345d3e6448b");
            when 22118772 => data <= (x"089a149a50311548", x"6152ee19ddf08536", x"fdef30fef562e2e1", x"37e9d2df0bf6b1f0", x"98373e59c97f8190", x"278aff70e19c3dc4", x"672dee6e848001fc", x"c96d8f5b677d80e6");
            when 14081567 => data <= (x"a1827439da477129", x"faab952d4ec9f8c7", x"6559f2539712e612", x"f71f84f65561dbf7", x"cd3131122088bd63", x"131c031741e4a248", x"96e6339162365d7d", x"4ab2db966160063c");
            when 7282892 => data <= (x"613167371fbc065c", x"c712b128a88c9f3c", x"812fbacff948a2ba", x"276a874f27569ca5", x"2783a950a2338de0", x"a3c2f0066ddc34af", x"ebd6251a09ee8b9d", x"7f93336772ed7a66");
            when 26349561 => data <= (x"92898154909e8905", x"8dbf99c28973699c", x"54c1a8f4468f4183", x"d05f495ea9397e6e", x"dbe8c639833f013b", x"36ee89d285c51ff0", x"7cb679041b85cd94", x"283237a581277369");
            when 15046417 => data <= (x"84da846d54226aba", x"8eee7b109a6e2f11", x"cbdd096eae2d2ddb", x"8c8c0677c67c8d27", x"58fb51c5cf25f292", x"2e4c5fd0933c971c", x"0e374c2d856ec74b", x"b263f939e24c682e");
            when 28533709 => data <= (x"25e18f47b18af1ab", x"26b553c866d85f23", x"a00d0473e2e0a4ac", x"93e3cf92901c9af8", x"5c6fc1deaec026f4", x"4d12d8d808fd7428", x"8d15a9228cc1b77e", x"067b37002390b6f0");
            when 3068806 => data <= (x"1ddeb4126584b380", x"a0272f7adb529c23", x"8c0447adaa95bdd1", x"0d66057673ea5717", x"6f09d6326b97d0e4", x"c63fe52286ac1bfc", x"7111b90dbcede6b2", x"9b90798705dc3c6f");
            when 20401837 => data <= (x"c696399dfaa50255", x"399cf232e8fb25bb", x"aaab908b0f2f0e30", x"869eafae2af3283c", x"8b6455b90998252f", x"2c94b8dccb1bccab", x"89c5fb76cad0edcb", x"f96e978e36acf969");
            when 30716733 => data <= (x"918c2c7cf9cb2a69", x"07d522ceace4dcb7", x"487e8dc850193b39", x"7263ca7761d99c18", x"38840147c374b31b", x"ea66537d42f14a35", x"04f5e67a777cc698", x"12ac601ae7ab282b");
            when 30541592 => data <= (x"ca1685d7783ed306", x"189edc8a1c2a0103", x"d76e932c28440a5c", x"0964665914c45d47", x"a8018c325a8bffe6", x"e4bc3c68629ded0c", x"2ec0d6bf5599a52e", x"7d2bd8cb510e049e");
            when 30438408 => data <= (x"e10a4a5978085290", x"3d1b69cce47a86fc", x"ea69b32e3cffc625", x"f41a6d1606d873c9", x"cbb5147b72452a90", x"98c199cc33b2d3f7", x"924ec7d3c407f922", x"98d2afbd9c696197");
            when 11616193 => data <= (x"5e66dc741fcd4411", x"580cf6809df83d16", x"e69e6922411cba80", x"b5331a9392fdf19e", x"bf35b922a93f947a", x"3ab533543d3a9916", x"7e2a0f848f7fa50f", x"7546a102c34606b8");
            when 10903781 => data <= (x"c8dd9cae56d164fc", x"9ec73831c919b201", x"6e9277998c04144c", x"274a19bef13c7b91", x"d4ac4cc62ef6a435", x"7fc32c90ea452c3d", x"68a7370cdc8a32a8", x"5ae62410e06ec196");
            when 25800526 => data <= (x"8be18efb091ec1d9", x"d83f31faac136d83", x"e8748951149dad3b", x"d5f996b681e57af1", x"8d346ea3cfe7c1fa", x"2a31a7f00af58c84", x"76a9de6b240f90c3", x"6b170dffe50a5d77");
            when 25333783 => data <= (x"93d2d6232596712e", x"3de7d31d1372fcd7", x"56d6fa943f444396", x"6265cc38cc6d9c45", x"7c3afb694f61f5f9", x"67672da818fea476", x"5d91a450d30575ef", x"14ed60d5bc8a2775");
            when 19339462 => data <= (x"66325621d3a3ee55", x"fda0800b76cbb058", x"02cd49d5339f6f2c", x"e52da1440f13f59e", x"5e87450e5822d859", x"ebddea719826958a", x"cb6342fd7db33f4a", x"a711b23aa036ddfe");
            when 4224312 => data <= (x"8d72f77e287aa19f", x"c4c6a3fc5a6e9406", x"bbf6b4555465ca14", x"89823c25b1b2c30c", x"ce4fa3f8d68b146a", x"f90c48628520fa04", x"9cbbd3377cd4f387", x"07f13f7698f7fedd");
            when 7093516 => data <= (x"61cf14f2627e9485", x"0f6a30dd3ff8e484", x"5d2beb0cb42de198", x"a480b97061cc0ee7", x"26c75d86599131a1", x"34af29b69da46b62", x"2325f92360ad54c6", x"1e47454b08d47e73");
            when 32660546 => data <= (x"523ff236322e1bdb", x"923cab60667ff9d0", x"1455cf4f799ed10c", x"3291b6553ddddde3", x"1ac4dee74cc841ba", x"04ddf638cde660d5", x"12aa2cec3ca69374", x"75161b4eb8ca02c8");
            when 19391056 => data <= (x"796bb6210ba16aeb", x"6665c0dfb180dc8f", x"180a90beed949958", x"5a1d145b81a17992", x"80e3462259525cdb", x"eadb67638096659c", x"9930eb86d9bbd8d1", x"e9f2b3f8fee0b273");
            when 28897036 => data <= (x"eeaa62d84b23e15e", x"989efab713c018d6", x"d0a6b64aa330f55b", x"cbfd3b18b08307c3", x"b8a50f881ce7da07", x"fb8c80af1cf68715", x"c993d3cad15f599a", x"f4ec1626025f2af9");
            when 2393752 => data <= (x"0f5081f015d32dbc", x"0beb1ffd89793bd6", x"db0e3ebf17fccb96", x"e247fcb7c5dc20e0", x"9121ac72dd0950f9", x"fdc491dee5442319", x"236a49ba9ada8873", x"c169e4049a503474");
            when 31589509 => data <= (x"f37d61e9d2ac0b29", x"4de96f16d97f0566", x"b13d5aa94d9e4cd9", x"ce6270af26498198", x"689d8a36416f7582", x"56eb748eddecf09c", x"cdbc29211b75ea78", x"c041e7991f740f5e");
            when 16836318 => data <= (x"bf8d76c425dda015", x"8222d3551153ea5f", x"7e20e98de32fdb60", x"ec6527c080ffe464", x"40fffb0ffdb2324a", x"2e5eea7a95d7e0ae", x"a8cfdfd92b59f034", x"4994d8baa6a52689");
            when 27870201 => data <= (x"ee7cbc9606fdea39", x"89865966a698c2f4", x"cefd5c744c1eb5c5", x"df686c82fe595d51", x"a94d4713f58e6b39", x"7157dc1740d4f1a0", x"b0000dda71d7ffde", x"e28e7791f2e9f8cf");
            when 13853901 => data <= (x"f5c14071d01b5fcc", x"66cac92eab54e8b8", x"5358ba6d83651156", x"a0bd3ccb4f47a058", x"3384d9df9e0ab276", x"a85a4a278a34fadd", x"f371dc355270cc3c", x"540a30e642172c48");
            when 14873705 => data <= (x"c9cc1cc40e63a3c2", x"e848e4ac7e7fbbdd", x"34d9eb45e4a228ac", x"f5ae3da07a3e9c73", x"9c19f74b7a40e5f3", x"3726610f734fe38c", x"a178fa29e24fdfdd", x"0327f6956a1984b2");
            when 20152621 => data <= (x"2094f21bf3bec1b9", x"86b61d22512b200c", x"c1446567b0ba6529", x"3370a3deefa02b8f", x"0535b0ce3abb2ffb", x"d03a418e95f01323", x"62bb2337f597593e", x"1917c59e7e880583");
            when 32164966 => data <= (x"51b28fd9015a7b4d", x"bc4db2afce709463", x"5d0e8c49d5ea4688", x"9362d8779caa7562", x"8e94e70a44316b4f", x"17d7ffd4fe958ad6", x"df497c10d747f069", x"f652d27a5b2f9ae7");
            when 10719813 => data <= (x"4d8c4d810c190f89", x"c20cb57852a1cf90", x"05a8073a4719aebc", x"422fac1331486503", x"d7bbdd659dd4747b", x"a294b0d2dc91db3c", x"b671c5daa725ad4c", x"842b174558322fdf");
            when 1795900 => data <= (x"5a346ee42213388f", x"e6b41b7c193f392a", x"7775dc7827c39a01", x"82e40df6b756ec35", x"93008dfb9bab6c06", x"26a313caae06ca15", x"e64decae0c0bb1b1", x"f37fd3db7d66520e");
            when 948232 => data <= (x"de446e7d5a2b0361", x"4aa5888acc4bafd6", x"0e5ab85fa84dd616", x"18347eb4e1cadfab", x"bc495daba7610f45", x"0502cc46e8e3f7d1", x"65e2eb6a74b6e59a", x"bc5edda28291e098");
            when 16158194 => data <= (x"9faaf3dab4e96f81", x"59a79b537f5499d1", x"84269f508eb75fb4", x"358ad7f0c3c0a9c6", x"ca293e0bea7e0c28", x"65bc54ea15b5a30a", x"98a7049d89c16f97", x"8703dd7d3ab778d0");
            when 3512837 => data <= (x"ee032f3646b7686b", x"fa135f7fb765b897", x"d3322676f945eee4", x"313df8576cf51404", x"f5ae5c183b08bf28", x"46ed3003d73a9314", x"699375fb8069c3cd", x"9ff75191b6132756");
            when 20788342 => data <= (x"27c9e8aa7045b649", x"a98efc0792d575c9", x"9a171c2dac1fe904", x"0635eec2358f864f", x"ff1cb3707112452e", x"f4a774dd303d8aff", x"a27138139157d689", x"c38d06fb44d7e356");
            when 5164888 => data <= (x"e5ef15549895b45e", x"365e8cb066041e41", x"e9aad6093455d71a", x"b62745e78f8b2d6a", x"f8185baaa07f9036", x"6dcd8026aa93d8f6", x"4be8811eda53e5cc", x"6fb23c4a09022ba8");
            when 22205821 => data <= (x"fa0e0af7e95f2e7d", x"3961c3f3165809b8", x"a153a22f66f7643b", x"d0a07c0446e8af5f", x"1ec6ca67b3fd768e", x"b4ddba4b8748b714", x"3c1c982f4dc980c4", x"b971b4b761566638");
            when 25290133 => data <= (x"bf1b670dfd95c529", x"25e8bdf55dc77a53", x"0d2b68e271014b67", x"f8b3c353d30222f9", x"b6bada01bfb84399", x"25e5f4ad93745392", x"1c51662695917727", x"701728bc232badc4");
            when 6028066 => data <= (x"46b3508a18c4875b", x"e34bf3fbd08c8a90", x"2c5d79487111194d", x"07cb2fb133269ae7", x"210ddb4024d51605", x"a491c2ddb6165371", x"d105015b83fb004c", x"1dbd63980793fdd6");
            when 2168537 => data <= (x"c917339f2ef0de07", x"6f703e013a9b8055", x"419d3581103de0da", x"67a1f6d5d7fe4fcc", x"f88837353f609c4e", x"b1e31f21188166ea", x"6a65cf33d8687771", x"20c934a149715598");
            when 20644804 => data <= (x"d7a661839ba6c298", x"fef241beaeda148d", x"bf2873a61e6a9146", x"855ffae11f7a1638", x"a5fd7fa37012fd22", x"28406c4a30c5fe75", x"b6ca2d1ab42f876a", x"5fafe0665c307d89");
            when 33559397 => data <= (x"c496bcef645953e1", x"1540ffe852a1640e", x"51a831b00d354e12", x"3b5cbb91aa24f150", x"18e45dd8761e72fc", x"d20be52450f66cb6", x"f8d03d0b4b835060", x"d22d918cc7995f76");
            when 13477693 => data <= (x"4f09a56142cbc8ed", x"d91565807b762685", x"85f70a919a9168f2", x"40215382170fe999", x"5683bbbe03995fad", x"1d80adb7787cf20b", x"77aa5e51fd50976a", x"7284a74ad21491a9");
            when 8197870 => data <= (x"639a0da6bcd4e878", x"d4f74a3fc4e1a3e5", x"108d35bc0558a5d8", x"b0aa2b220b5fd91c", x"f982a7ed2b750e96", x"0595783ccf38e5ea", x"e768729a1af41f38", x"617b812d501d351d");
            when 33210452 => data <= (x"6a5c59e0e848ed5d", x"15e47cda355f9d60", x"fcf8c16b4297ab34", x"b574b62cdb076a28", x"d1a9794e17653aef", x"cfc1ef4a670c041d", x"d253f9e214b52be4", x"c83aa1d2bc524153");
            when 27337034 => data <= (x"bd7300868c98ae80", x"a4f717073efba7bc", x"c195772548daa47e", x"78037616a7142e1d", x"63f270a93251d8af", x"3c01cee9beccd32a", x"35d5bbf955eeb5cf", x"4a62731924a4ea8d");
            when 7042234 => data <= (x"d27fd8ac3d27857a", x"600a5598cd4e91cc", x"1dbaf9a66d345e23", x"45eb8f9f0da2c2c2", x"7cd0175eeb53f833", x"a8b5eb90e52fdc84", x"7da0f085b4e1c766", x"da58e4faa8877799");
            when 27539762 => data <= (x"a35a18bb01b98373", x"139723ac9deca287", x"ce51546e0eeb8bc1", x"fd1e93b6996c4e3a", x"e93f7fc6390877a6", x"f47b05220cf91976", x"9f01d1d2cf4d7f83", x"177e49359e28fbc1");
            when 22148291 => data <= (x"f4b8e22f0e4affa5", x"110523668b47e9f2", x"0d1daa7a35d756ad", x"1ab7a75ace82af59", x"804f3d4ef514a81c", x"ab88c27da4513203", x"1cb72677b8355c46", x"ad5c09a03877ce1d");
            when 23174339 => data <= (x"ba5c0d4bc506a724", x"64194768849609a7", x"1fbce24a91f6a8f5", x"a437247627597a79", x"241b15d0edaf63f7", x"25b5868b361c5498", x"d789e7b192b59855", x"930c927e7e01b4f3");
            when 32735601 => data <= (x"843a1b7db9b918ab", x"0d7825cefd02fbe1", x"736b955529fb9d19", x"925e400d3df4eeca", x"c1d2c8b4c2da44ac", x"542ddb4fca070124", x"db9a2c3580e3bb54", x"5a04e02fcb0b1d91");
            when 28312521 => data <= (x"279c8c31c37a7ce6", x"d1d46d86c35f1c59", x"06492d4aa75e9143", x"e6627bb84a1bbdec", x"1d6ca0044cc1b9a5", x"3667bc3d131f55b4", x"0f15526b5f510332", x"e064414bc82fe41c");
            when 27281984 => data <= (x"7a65d5d5ab3e28c5", x"3e1962c7f6342c03", x"dce88122de6e7c74", x"339c16d3ad5424e6", x"d4de3f5e19b04beb", x"3d2e647399537ded", x"70cfa68c0a814753", x"a6018605029089ae");
            when 656410 => data <= (x"161aa88ea0935914", x"d42c566ac30ef162", x"1be5f4b50412474a", x"8d67d35cad6424dc", x"468398d7a73e4427", x"e0ddcbbc755c16aa", x"964e51af5b6304c1", x"e620e66f5483dc8f");
            when 18456948 => data <= (x"daed20b01a19af75", x"7ff9ab7a497e3fc1", x"d9c0143d6c2a42c0", x"59417d2277fc4efd", x"e71617cc01874151", x"6bd1ab033d6a0dd2", x"234ef50f8b90c05d", x"d3f892a2cce0628b");
            when 29450197 => data <= (x"f2723e5d46fbebb2", x"e2ba99611d68a444", x"20f696b300cbde6a", x"57775abe96edb448", x"41782caac79bde63", x"cb723ac5f1fcf94e", x"74a03805c2272926", x"cced65b6f9125db1");
            when 20766334 => data <= (x"f462a02683fb1d8e", x"affa64192061bb12", x"004a45245b40dfb0", x"6943269e76500e13", x"1cfb0fc4218e886e", x"baffa2e3ed8e7292", x"2d21cb5938a7e4fc", x"76e650c37b3baa9b");
            when 23739536 => data <= (x"52d1b3077a031d78", x"8f897f7b779469ff", x"f78c919ec40a6117", x"73558f4e8c628d2c", x"05369821fc8de1d9", x"2d8b355a5f3b8971", x"cdfed36af0cee504", x"0c0f14541250081e");
            when 6003028 => data <= (x"887a476e1ce06473", x"5697976a82bc3c93", x"4dac0669ffe3de8f", x"1f80b5ab2de8ddc6", x"ee1eb5342975ec61", x"b61cfc40829cc864", x"ef7a6df5acc28b40", x"c48304db2deb58e6");
            when 17694967 => data <= (x"9ede68234c5db219", x"1f3c1bd53e6421c1", x"db26d401920e3940", x"46a8cdb3ab2e1e61", x"7c260f932972b314", x"63ba251687acfb01", x"cfb7badc06b79075", x"ffae43f5287223c8");
            when 7055508 => data <= (x"9dd7e60c1cae5442", x"f4318d967dc65a6b", x"da39e5de83ed1540", x"d282148821a7548b", x"8ee80fc1074984cf", x"2d46fc2d5f5d7b96", x"e446a7d3c8997adf", x"057ae0cc336a43b1");
            when 1730613 => data <= (x"46b3c38497bea650", x"dfb15b4d569fa530", x"253aa4c2676c1eb6", x"1edcaff2c1eccdb9", x"cff9d89a79715837", x"90b324da4f6d1b1b", x"3367891915c909d8", x"3de54dac4e3c53c4");
            when 19584203 => data <= (x"7f5412c2122e7357", x"d947da0db71ac4be", x"9da2700ba2e816e6", x"96360ba02236f9c6", x"737deb0b453d94c5", x"1b9088cd90f5a5de", x"a550eb7d2c023957", x"ee60c728c5f4924b");
            when 21913479 => data <= (x"1ecb6c49744f51d8", x"7710f3a777629d71", x"7f6d82d36948d42a", x"e7c0bf27b74bb6f6", x"4d947f2d5785ef15", x"bbb4818c67f46499", x"6d0caba3c068c3eb", x"c89c52fb51f9b11b");
            when 22961438 => data <= (x"b0cbd5427bab9162", x"3446a7412b4a61d7", x"f3f1b98106067336", x"836ff630ed7f33d7", x"136d2acea172ded9", x"15c345257ff0ce32", x"8d1caa2b4f64652d", x"d7d95e289b132129");
            when 24184044 => data <= (x"16f252d5a4c6c541", x"fc2b8a4d74323f67", x"8141cd2bcab1aa16", x"225e378e91c15917", x"6b574ffadd0542aa", x"8909edb314a2b236", x"6bfcdeb34b868c44", x"6c6093384ef0c43e");
            when 29801796 => data <= (x"65b44e1903e4f9de", x"f91a99c9c248df75", x"a934d16aede40d82", x"25ba928bc374f9ae", x"bb91c7d000d8ca85", x"576c7dfd67aab65e", x"3e1aac1b1cafd0d9", x"04d390409cc61def");
            when 1773884 => data <= (x"7b0f5d8037c498ab", x"0816b7870692de1d", x"294439e533f4da2f", x"deeda9929135bc1f", x"c91bcb0e12a073fc", x"3c920a5bf225e22f", x"cd162488c27b70ff", x"a455da073ad67a57");
            when 14645945 => data <= (x"02c3952d6cc2b394", x"c25e37d94c183806", x"bf69a3058b989c79", x"1c3008aaf91746fa", x"aac05e925a2b3169", x"c40f6139832f8e0a", x"db986ca1cbd681bf", x"5c2c39e6f294f2b2");
            when 20896798 => data <= (x"9b0e2893248bd147", x"1dc7c703d38ef4c1", x"9f1f0e69987744d6", x"edef3cd1e2ea082c", x"1fd28b8829b7f657", x"e64f804605217e2a", x"45203385b27f7b96", x"f43934e2cd328757");
            when 18269572 => data <= (x"3c5b17da60179bb8", x"b96277adcc01da30", x"6f17d5c8b1120c88", x"cb03f8396a13e6f3", x"2863ed0cc98cec6b", x"5fe977e34e2f347d", x"4ab4189d6b143869", x"ddc3a7ad82d33033");
            when 3685588 => data <= (x"0aefb35616b3f417", x"c6716f2c53e859b1", x"1a417fd4cf9d920b", x"c9e64e56774348b8", x"e40e9d7ea98c584b", x"5e9eb44bb41fd8d3", x"03a481c3a93fb428", x"2065266e79f75e9e");
            when 17588051 => data <= (x"4b2f3eba68e8cf03", x"0b8830db19e0d91b", x"ccb9ae454101f5cd", x"6abe851d3cb5a8f1", x"f9037cf737ef1ffc", x"e73f069528c2f7bb", x"f5269049e4aa7641", x"315cdcd94c811ed9");
            when 12335682 => data <= (x"520f6866ea5852b5", x"9e512527b43cf593", x"f28c5f7065072272", x"37097996e8866109", x"57b0ff6b0d098f1a", x"dfd087d60a84ac96", x"b2e6a7ef4d1f1979", x"095b13345e7b2d95");
            when 27334602 => data <= (x"b9f550fa24d53095", x"fe0f9e60474dfa65", x"042ddc4ec66906cb", x"637b6f455453c4ad", x"8a93bc4c39521b9d", x"cf6d622e599b1bba", x"72b276c6636f6eed", x"b1434ac80fb06db5");
            when 6170734 => data <= (x"ade5ca5e2fa29d0d", x"26e53a751a749d7e", x"da6e209ccee2834d", x"3980f13610198f74", x"948f17ae3d71fa35", x"13db28127dcab150", x"934d65b0a9b5a377", x"af9863a204c57212");
            when 12950574 => data <= (x"09e8a3a039e91495", x"02b7dd7fd5aa4779", x"40cabea4a869e041", x"db2449dd4952f0ab", x"33cfc19c45fcc1aa", x"a989f4808636c2db", x"27d14f6d96562428", x"92c6ed0688a108df");
            when 2599784 => data <= (x"91a8fdef5fef8342", x"507d13c08cf63538", x"e14b7090856ed910", x"cf9c9af1a560f5b7", x"0463014ac075fa3f", x"2443104a77b25802", x"9ca8117fe947b7df", x"a0d12f450d551f27");
            when 18557386 => data <= (x"6dd729d611366282", x"3cb8b78678c5b444", x"1d346b109d376681", x"841cddd1b4f48e8a", x"2f28d36f21d43e58", x"3f1e5fe80d7a32a9", x"da4d64802b70a531", x"249b873c6352a28b");
            when 1631986 => data <= (x"d8fbdcc913d4b02e", x"6c0757ce309bc1ec", x"431162591fa2bc90", x"2969442260266c4a", x"aa35dca134e9af8f", x"e3d280fe6d9ac2ea", x"5f4a7e6f9f27e829", x"f4b8be5720966b76");
            when 5124752 => data <= (x"831b7e87f454a9b8", x"5ef8538f971a165e", x"c757d2e7ed76a72f", x"db29ef9ff207806c", x"2e101062eafc5124", x"2ee54b9aa1b41bd1", x"12b1f190358423b9", x"994887ea715e0b01");
            when 4232231 => data <= (x"5716815e562b034f", x"c2902a3c3aebc082", x"27f0a2857c9e9c10", x"e5bf65428cfb2a43", x"8a62e27fdf51413b", x"fe8a30eeca38a309", x"2c0d9eade2aeeba1", x"ce859762eb2614ee");
            when 1089777 => data <= (x"2c5c2a3c82cf8dc7", x"7e9d03f466374602", x"8b9bf348b4db5499", x"271c68c77ebeaebe", x"a2cb31d462293f2f", x"27d780b0f5632b04", x"be9c66bdbed794d3", x"b5bc66335c93468d");
            when 25477805 => data <= (x"78bc5e19003f37f1", x"cd21437b4ff43192", x"1e91abc78174026f", x"1fc11e9265cb9243", x"3805bfbc87a92ed7", x"deb5692e2983c914", x"a5dfdc65a3c33a31", x"f60c6d5c6eb91d24");
            when 4339298 => data <= (x"c90ed6f9cac12f32", x"2896a8df5d389cb9", x"477d13cfdfa7bb2c", x"9bcc8da221e6bf18", x"b03e0a2c64813836", x"5cb84b128575c99a", x"2458aebb9a8ea581", x"2bbc61ce5c176fce");
            when 3413178 => data <= (x"1b812becf197f24d", x"1fa6df5acd15d56c", x"d7e3a51e1f41409b", x"eeeaba724e1f095f", x"9524c68c3b126493", x"dd4c5c376e3a4f5e", x"30722aae592e2039", x"b78a9d2b9d42e2b7");
            when 20882454 => data <= (x"0b6271fdf9f31ae2", x"565b3c4e719b7230", x"ce43d3626392b80d", x"f518304a5b88b170", x"a06b732913c6eecd", x"769427e679af747f", x"68d06c50d687902f", x"e6527177793f4618");
            when 19455541 => data <= (x"befde46ac03e683f", x"0724ea9f53396ffd", x"e0b366f211f9e37b", x"06ef55adf5d9d907", x"5b5a092ea3e609a3", x"f3e7f1a06d9822ec", x"d2a6f701e453cceb", x"1ce39b23796a7aca");
            when 28931959 => data <= (x"1856c6ef315617de", x"dd54dba70c0afc05", x"b70d7497f03e7864", x"0d67ac78e4b0099f", x"5066ff28e85e15f4", x"fcff98a56d3cf5d4", x"cecca9d769e13352", x"3f3cf7647611eaf5");
            when 8453494 => data <= (x"1fc251547477af27", x"1a39f785aa252bcd", x"56ba771e97ee8a36", x"93c92238e00cd33e", x"d03e85302091dcfe", x"ba67bc1e1b8e1304", x"560c5851424198fe", x"31c7d25eb855bb00");
            when 8964829 => data <= (x"add0dbe01a2e50e2", x"3abc4494e3f96927", x"f7eb726789f48e20", x"5a1c045527ea803d", x"eda01a5e5f707a74", x"0048a61b556f3272", x"1aff10eea2360c74", x"db306716f5180db9");
            when 12004042 => data <= (x"01b8c0c506f7878d", x"2ea8119cd5dc23d6", x"376d4de7c069385e", x"9abdd5f664f876e4", x"4ad20eefe472f005", x"e4913ed0ec0dfd83", x"6a28123900361d82", x"16bc4037851c34a6");
            when 11567615 => data <= (x"d49843cbaea5af86", x"07627f77117c9cb1", x"1c26c5602292b665", x"ff01135a991e14e4", x"0e45d2574db7271f", x"0b0613626652de0c", x"7707422e5dd69c4c", x"f0af5fd34852b5f4");
            when 26613135 => data <= (x"ecb3dce2ef99ff9f", x"e63897875e61c645", x"4dcdb8b184dc4fc5", x"8a1c7d691c18d44b", x"48e88ae7bf78eaca", x"e6b5c82aacf14b85", x"09fceccebcdca987", x"23fc98b0b1ad738b");
            when 18050700 => data <= (x"bab4dce1deda8b07", x"5a16035849a7b3a5", x"a58ed7c24e44f634", x"a5e7263625b81bd4", x"efb7e8c9298ec5f8", x"0443837170c46596", x"3adf9948bcdcefca", x"1b95e7f1fc1eaad5");
            when 14790511 => data <= (x"3692c1c2e82ca7d4", x"d7bd9b8d240e89b2", x"2b06f0b5d8dbd380", x"557084c7511a9fca", x"8409c5e2904a1e03", x"911e6fe2fbcdbc25", x"9a78548a221d460e", x"24080692415ee70e");
            when 30503661 => data <= (x"f743633f691d6a39", x"55b9ba0fdea3036f", x"ff23196032db9b98", x"27f547582bd8bdd5", x"ef429ce390544f35", x"c20b0943f8ea4b86", x"05c18d9a0ede82ea", x"c9e96a9d2495954c");
            when 18443963 => data <= (x"4a3703ffcc5d1eae", x"08b01a24d1854da0", x"c0d974177dc6b79d", x"df766f6bde515244", x"b70455d623d069ca", x"f8ee0dd1f6be5859", x"1a00cc5cc37d7b6c", x"9f521717c54ca6c1");
            when 25578891 => data <= (x"2fe96dd388d74cbc", x"82dc318dfbb26851", x"7a5d44d812e6963a", x"066308723bf052b0", x"fd0fe0df27ae6077", x"518691750d38f35c", x"48451c1e260496a2", x"1aa9c9a2e590e95e");
            when 22295771 => data <= (x"83f26e7d0f3d6e6c", x"2b29f698b1770aa2", x"94761d2bc60bb48c", x"3c83148da7f9b5e0", x"9745e60eda961908", x"7bf6ce04d02b73a6", x"dfef43718a4bed07", x"30ec965b7f147588");
            when 28304443 => data <= (x"08e3cc39ca2e797a", x"3e3c7ff0dc3607fd", x"778107fb7fc65e72", x"7d3e93890dbec136", x"12da150f1baa3e9b", x"c26d5940b49eea36", x"36d90c86be0c4820", x"d03321269c60d974");
            when 10542421 => data <= (x"a86c17af6cc0a793", x"5f6d7a3333ae2288", x"dafaf2329f90fb04", x"26bd6a3c1c142869", x"0aeca7e970db275d", x"4ea2f295803a68d1", x"73d8d44a5d3bb4c5", x"c90ccb56575e1e4f");
            when 16482995 => data <= (x"60308803381a6d62", x"b3b4f0d2242f64c6", x"757f16bca8be27a3", x"3624595ced32cbf3", x"568882905e828e26", x"a5e93803f52ee595", x"fdf7679b8e3a50d4", x"7bbc9dc7392c4cc0");
            when 15243680 => data <= (x"03c19c1a85ae94bf", x"0b1ae62f0d43ee65", x"dc0bed6ed7e06ebe", x"cbbdfaa8159071e6", x"799720135fcade60", x"5abd1ac51403f2a6", x"2dd592bc2edc3286", x"aba55f3d3a59f52d");
            when 25904383 => data <= (x"a6959113c253a4e6", x"54dde2b9619a16b4", x"cb52f02d5c07b443", x"46d9a256db885500", x"527fbf5c2e7c9d51", x"7e631aaf52658c30", x"586e7151a3ea2767", x"8d5cc4a689af85c7");
            when 31386642 => data <= (x"68fd1c05a28f74b9", x"5bb37d80cefe6bf0", x"756860d96b4219b5", x"aeb9293a54aea545", x"8b58ffadf74ca2c4", x"cc4d0fbe15ff6c74", x"86dc21597dfa907d", x"ec4996c9cd7d5082");
            when 780087 => data <= (x"ad4fea541369dd3a", x"1d355281036f609e", x"5c8e26737dff657f", x"5a77a7b48ef9bfbe", x"35b59cf2452d88d7", x"7747b61113e0a2bb", x"0d45f6f869643d50", x"c803adaa4fbdd6cb");
            when 2872768 => data <= (x"de5ac7b55ffa09c6", x"eb0cca975fbbaae1", x"4f94d576ee5bc055", x"fd9e660cc4ce8487", x"2cc9822ef2afe221", x"65eee2fd892df8ee", x"24758733d4d52b71", x"a1ce1e312eea4f3a");
            when 624416 => data <= (x"b7eb4dc590dba02a", x"6e97ffa23da4abf0", x"68b9b3fdee6604c8", x"da9c4cdafa410974", x"5a05b0b33dd079c1", x"6d9e818f3fabc143", x"17363e4b4a2a0181", x"e3935d265510708c");
            when 19972512 => data <= (x"edb7946e15317156", x"9213a2da63931595", x"f2c0359c494c1661", x"fd950359397cac66", x"8a35671596d4aa76", x"983cf7c9d914ccb3", x"9b1574dcd72564ec", x"2aed3f4bcb74fb31");
            when 13447825 => data <= (x"38abf60f52ae9aa6", x"17fb65aced5de666", x"9fea2277e4d34f28", x"5484946b08e0db1e", x"fa73436ba2787bb0", x"9900e1b1c36f8a99", x"0662a43ea3dcacca", x"ff71f72cb3674309");
            when 3679782 => data <= (x"3c87f7190fe16b83", x"9146c7b873449d6c", x"9e79b9b55bd431b4", x"267b9d44d4014141", x"4984bd1dc6b89bb9", x"0e193f8b835cae42", x"d35b7f0ae1ba745b", x"f40868736facb9c6");
            when 15907946 => data <= (x"d881ac293acadfe6", x"1aa9931db7b498e5", x"a81525024a4ac5eb", x"7d1c0f8a61da4327", x"511edcb7250eab52", x"ec59ffd6f9467be9", x"477d7f2d0d071e92", x"b9dd8655d87dd8d7");
            when 18545540 => data <= (x"a9652e76698ad1d3", x"608784c612c82115", x"0899df76973c2c3a", x"c9982fd460aaa2df", x"c0d75c0594855f74", x"89b9b1bfd3d55f3c", x"776202d55c00fd8d", x"6dbf37850bcafa5c");
            when 14035587 => data <= (x"f2f46d52aef72939", x"45335970bf1d6d18", x"dd595440b5eaee72", x"1b93cf48ba8510a6", x"a99c9155fda482dc", x"30b9e3f6ce55554a", x"d5df7bc456c3039d", x"7f887f5ca9832a5f");
            when 7117721 => data <= (x"152472e44227d666", x"2a8d5006015669b9", x"3e95dd16bc73d4db", x"1c9c586389d40847", x"3ff3d0714fde8020", x"2344f066a6ebffc8", x"e897d6990dfefe80", x"9bdedc49b1aad332");
            when 5593467 => data <= (x"8180b4d307604d51", x"a21c91ed1b968f40", x"97fa767ba1f1c361", x"1a2c824c94dbe9a1", x"41f8957578225735", x"3dbf2098ff17b060", x"0ab46df1767da5df", x"45186093b442da6c");
            when 11945598 => data <= (x"7391b6e8a65f7ea8", x"3964b2934d451a9d", x"65d42d780c7d2423", x"b934c248db7607e7", x"db670cc89db76056", x"536c383eb213ee04", x"1a6fdaec2cf29a4d", x"1c01366412dc000f");
            when 27843411 => data <= (x"e5ff132abf022b24", x"a71e150c9fea7204", x"478a150b3838e26a", x"fb09908213f85423", x"fbd0f1276bc9ad1f", x"d30933a5944d60a8", x"99eeb5c670f3703a", x"cca31d54620052a3");
            when 12741160 => data <= (x"1e43d47efd3d5f5e", x"22eb13787c0a6609", x"d8c6468b99030e11", x"6e90ca37e97a9ed6", x"b0ae92cc2cd3d5d8", x"0c78b478a3fda46b", x"26febd6e320e665f", x"5a0c1394c0e80ad2");
            when 19277993 => data <= (x"99f41c7e14498c34", x"e44c9d925eade6f8", x"2b549e9520394e9d", x"498bb541b64ff1ed", x"444d88451be40c49", x"8ae85d3db80f583a", x"c034f79d40d3f6f0", x"9cbfc88daef6a291");
            when 2292256 => data <= (x"0f42e44efd8484d3", x"42dd2ba1260ec0ed", x"5dec214629f0c91d", x"6aae93ed02b3aa1c", x"31e436dae2c5c507", x"a56dbf5f0a533f4f", x"3ea66b68fc450812", x"e8a251480c607d16");
            when 19956839 => data <= (x"739359a4f25d8895", x"2a402197bd92b0a2", x"6206efea53b1694d", x"46bd1c5b0a38d7e9", x"086e8da45cac900c", x"42a7c93ccecff618", x"c1b8a3c7a061908c", x"1d91e6d05a2d7fbb");
            when 15499191 => data <= (x"dfd107baa9249b07", x"8c9d5c77922df2b5", x"6eed923b5d2e217b", x"6f89231ca52e29e4", x"057274af7774a261", x"e8307cceeef826ec", x"03d80f74e8290103", x"3259bb2258d06e33");
            when 25278084 => data <= (x"cbcc75ca50d806f8", x"c207e27ed608e8f2", x"43cc46470765380b", x"647e4ea13ff17099", x"00db806c4e5cbc23", x"7d3a568f47a74e62", x"8c9ce55881cc6e7b", x"34f43167acdadbd1");
            when 27702678 => data <= (x"b57691ecdb91c71e", x"2d970220da3b02e3", x"02b970817ff10720", x"ed3e8eb8f4c50126", x"4d7916095b985d99", x"4ce8f156467b2830", x"3ecc0a8a64c1e00e", x"afebafd868e5dce6");
            when 1873821 => data <= (x"d796099c1625c8b0", x"c152ffeced649b6b", x"5c71b92bdda0b06f", x"63543eb324aebf52", x"c28ce7f05b3cf211", x"ee8f418e3a950d4c", x"4da31146a02d53dc", x"d66f3ca2e3da3f32");
            when 11808268 => data <= (x"e68a18663bf2ef8e", x"7488542b5709dc50", x"a7ba5238a428a364", x"4a6d7b05df41c027", x"db3262196582b77f", x"2440d7c2b0b9e200", x"dfd21220a6367233", x"b16edd1288d761dc");
            when 14816519 => data <= (x"fcb3896e5827a01b", x"33ffa8fa32ae8ed9", x"347113ecfab73adb", x"54d48a91d13f6ef6", x"ad3155234ac46274", x"8e624d903c8daed8", x"b542d80489867b4f", x"e756ff5d827d3251");
            when 22540588 => data <= (x"29b1501025342de6", x"87d55ec740668a19", x"5db68b32e654731b", x"bc61fb7262220fd1", x"311c87f782f59864", x"337eafa386a43d12", x"c3c9f2ccaddab795", x"c2be448c7dddd597");
            when 1550774 => data <= (x"0a7e6324d5141fbf", x"f1b75821be5a8822", x"066d8d784dacf893", x"9b26d457744cb630", x"0382cf6908c80746", x"99d14a1180a4957f", x"b3c6902eabffa10d", x"cb2450cb3be1e061");
            when 16210050 => data <= (x"6a2858655446e788", x"b3a40ac0bf155cdd", x"bd435e1757e58ce5", x"e7c6190d76409e54", x"d93bb03e0ff4e629", x"0f71432398139852", x"e60f32cb33659790", x"9a279bdeed55d13c");
            when 26970460 => data <= (x"80b69f499b03d95e", x"d38c92dbbc00c883", x"5384c79e12c85e2f", x"6d5febd6817bc118", x"caf8adfea1ec1596", x"afc11885494fec3c", x"6efdef2cede3ef91", x"baeeb2ad508eabae");
            when 20018910 => data <= (x"618a293add5bbd92", x"3ad489af8eccf68a", x"fc22281268942cea", x"d5ed032c0e81c38d", x"efca1796f3b05432", x"724b21671d01540f", x"1fbb1d25598b40a7", x"90f8eb39b14a5b4a");
            when 25688586 => data <= (x"9734cd7785fdcc1a", x"ef453727844bfe10", x"92eb79c0da0e5bb5", x"51d9234a3c42f639", x"31143062edf2021f", x"bf222eb4df561c3e", x"cc542ae4aae9c108", x"99e008ef9721e98c");
            when 31354062 => data <= (x"c014d071f4ec3344", x"589f760ce3a48e68", x"0120761889a3e516", x"f777d5d23e719789", x"4b5d1f75afea5f6d", x"3ca4419cdd57c373", x"a4bbe97677fa06e7", x"8e99420ff0f69b2b");
            when 8148422 => data <= (x"1aea757cff4dc4cf", x"9e4d5778a968250c", x"c5a4df380eae5e0d", x"ee6c75bcb160b1c3", x"c7dbba7a34f4222b", x"c5988b4219922345", x"cc20968b84924fe9", x"3364f5a3f184a5f6");
            when 32140193 => data <= (x"e3012047faca64ca", x"eec7c80b0b65955d", x"2313bd0e19e293dc", x"33cb59eb4e14ecdf", x"c8a68deecbd0b36a", x"497251f6f70c3a66", x"c7f4830678d1cd98", x"512aebc7d9114bfa");
            when 12453785 => data <= (x"b5095070ccd1ad70", x"b1d34165e10c897a", x"fca6f7245dc5551c", x"7a5c904425b1aea2", x"a17c9fdf74f11e46", x"6f899277b0e02454", x"58de72957849e73d", x"4cbec2adc20e7819");
            when 25764333 => data <= (x"fbfddc91f292d08f", x"dcf4cfe4d4e2410e", x"0f037d02754aaa92", x"91defe4986633ace", x"5e168749e4fd9ca8", x"b2984b3b5274626d", x"b7306f6e5762f46c", x"7dbb20b15927d31c");
            when 26193465 => data <= (x"eec3b5719fefbcfa", x"936f9f98b6ee8749", x"5a71b4e93a52be1d", x"992ded561e3e939e", x"9b8bf058c993cb82", x"aa851d7afdd61a78", x"c988b3914b63dddb", x"321bcb63396b638f");
            when 1425736 => data <= (x"016d4be485826097", x"0ab446ded02eaff6", x"09231461813f5efc", x"d69cc232454e589f", x"232fd189daab6986", x"4b1799e0deaa5364", x"92bb96ab34d99fae", x"353be0272e3a3953");
            when 4248736 => data <= (x"a682bb6915dfbd54", x"99dc97924f998883", x"d078970b10a9fe57", x"e71bc40ede9d2a71", x"c6157feb5451fa46", x"de94da8af83b87a8", x"bfb60451a68f16bb", x"3ca5488045755c3d");
            when 9014486 => data <= (x"b83698557af4f915", x"6fb343ee1514c0e5", x"bed21e6210c19eb1", x"8b806a67c440b885", x"dbe1ada66faf4360", x"e887ae9ccc476773", x"3398d23799f2309c", x"979e9885afe0e66c");
            when 20979221 => data <= (x"16303846d7c1e8fc", x"e21f0c392e2f2381", x"0bc848b19ecff0d8", x"be96b4e191fba9df", x"8af757eef5cc0b7a", x"e6c27b9ed48e7af6", x"e5fc60f8a20aca18", x"0fc82e351da72860");
            when 8315497 => data <= (x"34116c2e1544b16e", x"b8c7ab2a6b2c66bd", x"2bacc073090c448a", x"036eab1f63fffe4e", x"eb58f5fad55b8a82", x"c5f556242de3c3a3", x"05745dc0fbf6cd73", x"56aec6e61b0366b1");
            when 13488080 => data <= (x"0d5a4b8ed9f38f6f", x"6428f923abfa6ea2", x"53084f694aac814d", x"8a89c53067a79119", x"fba1204f8cb6d40e", x"0ead80e2fc6df8f1", x"d781db47e5e0c0df", x"c0f60e08ab0dbf4c");
            when 2521621 => data <= (x"927e99114b8fda0b", x"4fa341f925317bb7", x"68df293a9fc707aa", x"87376b9198624f01", x"3914a2138f50b2ba", x"570d0b9929e566b5", x"208bd25585131053", x"ec845179e21584d5");
            when 21726569 => data <= (x"dbde25322b160293", x"37b9206b9c0d65a0", x"586801d8761d1bb7", x"6b05f18619288f9b", x"6a36e5db48a3c80e", x"bf6f6996d5be2ce6", x"535a20738b97dcfa", x"bfef1e88fb5dba90");
            when 17378336 => data <= (x"fb25bc9cc78c686a", x"3eaab27f5eb0b591", x"bf296db40a264aba", x"f5a7536668ba737c", x"c76eef70e3552fee", x"bf74265bd92f4a32", x"3ba6ba623037bb0d", x"33ce0da1c1b803b3");
            when 6648651 => data <= (x"7b6b66fe67b550fc", x"98cf31c24b1e08ee", x"2349424b353fd352", x"70abb9b3ceaee705", x"9a6970b861036695", x"2502ce22e3ffcea8", x"7f822ad7879f2ec5", x"fd8cc011f8b16f85");
            when 18451495 => data <= (x"87cfa336a59dd04c", x"864b95b00e797bba", x"eeb07e8ca68b7ac3", x"491ab1903c534557", x"072b76d1fb3c7af6", x"db8a1cc6702b2168", x"2dbf9209d79bce5e", x"73a59f86e3339cee");
            when 27347467 => data <= (x"bb87cc78d0c7905f", x"f2d1547b4b7b66e3", x"57c9dc1a4a67f849", x"0d3c9a07f20770b5", x"3c44e8692b8e6ed0", x"d3348ee60f03a8b1", x"efd59ca1baeda621", x"ccd9f730659f54a7");
            when 8367805 => data <= (x"2be0e95f9b796261", x"206580ac3200fbc8", x"8e7b0c8268fde827", x"53925442ec59f4bc", x"33ab6d7555edaf2e", x"b113c5c274e2e7bd", x"e3a33cc96a0ea8de", x"378b268559d5e9cd");
            when 3178282 => data <= (x"2e3dc021521b178b", x"f325c26a06aca5b0", x"4f22c09f40eacba8", x"b8590acb2d498373", x"b7706dbfc6776246", x"4478521f3db8b56f", x"bd8a6ca5a1a0590d", x"c918666a4ae6449c");
            when 23151119 => data <= (x"a5f3952feed079f2", x"367f18242034333e", x"00f21e66cdbb70ad", x"0be3627889ce399f", x"fa117aefec5a47ab", x"8ca871016f983614", x"4edc33341474bf47", x"376e0c7b585fba7e");
            when 18457561 => data <= (x"8fa9f01899174838", x"347ed9d499f90cb0", x"7eb789b98863382e", x"ac3d9df96712f2d3", x"4ff3f097eb554acf", x"1bfb90cb27a09443", x"81dd238fcbb8bd6c", x"664e394aa07170aa");
            when 11212634 => data <= (x"db76033b3a0e7166", x"4d1212e00c03942f", x"0bf0c1ee4f0636c7", x"7f198bd54f883572", x"513319719e1bf61e", x"309fcd1a64abd9ec", x"ffdee06122f9ffcf", x"5ffb804c4f40e2a8");
            when 7838809 => data <= (x"86a4e89430317a7b", x"64eb7c8e21b7c6f8", x"3fe756aaf015ba92", x"6b9c52a547ea6b8d", x"6880b4b1e6509374", x"ed3038a3d3da92b5", x"4fff3cbd6a115f46", x"99882f18c31b6f4f");
            when 8353712 => data <= (x"649b14e2a4634eb8", x"22bd9ab2c5a9f63e", x"ecc95d8dcf6b42f9", x"85aa916963a38924", x"7994d05ea65e4471", x"3a79bab6aa9a8956", x"b50a3cd14fa1941e", x"40cb8e59cbda09c3");
            when 28521751 => data <= (x"58343a5347e08984", x"b64fd924ef7f9adc", x"d1efc24a9744daa5", x"971663f1a04c80d9", x"070b983b51e0e450", x"82c65b17897c70b4", x"57ae6f39989eed27", x"4a038dcf917ddab3");
            when 10314611 => data <= (x"f7fcabb8c924cc60", x"afa3bab7e19ade85", x"11600b755fdb1c15", x"f4bfe8a27bb58f8b", x"1ba31dd6e7e6b0ad", x"97d895edf2d7bc06", x"25a61a13dc875bd3", x"2c4cb1bc8e33acd3");
            when 22730172 => data <= (x"02b4b95d88b7340d", x"01c9da85feb8c30c", x"c770627211aaa1ad", x"a0ae6d3fd44df270", x"5032764850ac91fb", x"fe2effa44993f549", x"e0e46e41d182e21a", x"49a3f0ab030fd062");
            when 2202477 => data <= (x"7eb4fe0438ea9f27", x"7fff63be29d9ecd9", x"2242138f18dd1314", x"126c1b0398d4727d", x"fc6563def72bc412", x"94bce87d5c2614c0", x"19d144fb6d0f0c03", x"d30c1dcdb61fb478");
            when 4207183 => data <= (x"8d94e26bd78b3fe1", x"8ee9483dbe33b04d", x"b63cd69aefc24185", x"da30090c667519fe", x"3d4b93b01de8da42", x"9b354dbab67572dc", x"1457309a51ff04b5", x"6e73c87336064bc6");
            when 7113232 => data <= (x"b43e04ce108923d2", x"42ef11628f409bcb", x"ae48de3b8fceed1a", x"802ed3ddc67fb5ee", x"0889437d6ce77967", x"5033eae072d92368", x"d2f84f760274fdd2", x"3bfa5186bc0e7f80");
            when 11504494 => data <= (x"60e62b4ca1dd501c", x"357045084eb1f43c", x"df13abfef6d2c5a6", x"622c44b3b72b08e9", x"c9d421a4a12a0664", x"bea7bb5ed883ad55", x"d2d46b28e79caaa8", x"b8b96dd120f2f9d0");
            when 7154719 => data <= (x"968c4c62739e4dbe", x"920d56a857ddd54a", x"2db58ac058a679c0", x"105aa51ed906c14a", x"63c88abfda02c17c", x"d48614c2750f52c5", x"bff95c4a5c768c41", x"70ca729a209598a4");
            when 16350482 => data <= (x"6a98b80a6d0df1f3", x"1054d7c29ca7043a", x"3184fe136a78bc9d", x"ab614f94ca45895c", x"4013d9a4a4dab922", x"8386b3492faf6ae8", x"0a3215b455529d46", x"97b586575fe4af01");
            when 8056795 => data <= (x"262c9462316a4599", x"66f515b923cb7b86", x"ebe9527343056b09", x"78242567c9572010", x"69293c88be817437", x"3434685773f4c79b", x"b4fdb28ccf99c05a", x"c4d5d19c273d0f37");
            when 16535362 => data <= (x"bf66c616fa8503b4", x"e3dfee28b19e932e", x"337576a579487f6a", x"62b7cea030a681b4", x"392b3c4e4f8c2d92", x"8fd669386b650a99", x"674825fa1a60de8a", x"92c25fbdcb57d7ea");
            when 3022038 => data <= (x"4d25a64613989627", x"851ded4279d10355", x"e98df1a9adc53a87", x"03310b898472e9f3", x"5a1f397afdd7ee5e", x"6a8aca1bfc817a8e", x"de5b87b89a907348", x"e1f5474964b30760");
            when 3570894 => data <= (x"f97f373a0948ac95", x"4e2f3a7d5f1ed4a3", x"a143952ff325f0f6", x"796b506070b0b8f6", x"7e7bd8aa93120a17", x"693062630f4887e5", x"711a633f22c90f49", x"7f035ed69f4c2f5e");
            when 5164523 => data <= (x"85043fd86aaba4b3", x"cbb46beff9aac747", x"5c2d1e69fcd3b20c", x"db0da681a7801df8", x"268d29e002e82c66", x"f54061e078b5fefe", x"73a361fc409d4ed2", x"57d123622fd7ac29");
            when 23534158 => data <= (x"20cc5857e1e41010", x"653786a9063eb87e", x"c5120714d031bf88", x"2d9b053ec906eaf9", x"e40caecd9cf23b9c", x"5823f8f1b32d7c82", x"12dbc7618fe17440", x"7502001d68920ab0");
            when 10315078 => data <= (x"c05eee7d4427dc39", x"56b2fd4f32cd7eb4", x"f6534d44afb336a4", x"dd8deb68ed5b02c9", x"ee8a7cbc45f7604a", x"c6f5c465a98dcc0c", x"c9647539b410e174", x"fcadfe0e40452424");
            when 12282831 => data <= (x"bcbace3595c0224b", x"2d1638aff01c1952", x"72f1fa13e16546ee", x"0a42b4695f542a71", x"f1ca957ca97fe218", x"b372fab5746eb23e", x"51e8bd9d21c9b6bf", x"66b8ab16872905c6");
            when 7511546 => data <= (x"1698414e8538a803", x"f13b7f9290de4f52", x"f36cf6b00518fe58", x"9d08a5d416c55fbd", x"7e6d1b11829fa1fd", x"47de0ce699645a48", x"a6791c3e0e066f13", x"44056fa82b463a36");
            when 9340002 => data <= (x"89e062a351e79bda", x"79f6abcef0cbdbb7", x"96ba63857dff2828", x"8ee2493804c611e1", x"83adf2f58809b907", x"8ad1aa99484f3bfa", x"054956015024f0f3", x"a494769e89f28f25");
            when 30455990 => data <= (x"352a25868cf4364d", x"73366f1dfa643ac8", x"cef12f056f604b57", x"f380c10e0a352919", x"57c72df25023174f", x"4be9d5c76a770a3d", x"30ef513f2d3460ba", x"1cef366040c7de61");
            when 33368606 => data <= (x"2378e21922064a42", x"6e56490b49c3b972", x"e4fd4fb701fcba46", x"98c0de43db811b03", x"992f34322d72cff7", x"08f775498bce6148", x"bab541294eae79bb", x"b4f3e3de8716060f");
            when 11100789 => data <= (x"73ae380f5354dd70", x"d227276f23542427", x"3d5b71412b4938a3", x"c3a20cfb140d2aba", x"10432ec57ea0cf23", x"5ef89efa8fce81b2", x"b328afdf0361fa72", x"7fb8405ee891d8ec");
            when 23658918 => data <= (x"0ffd287943a53081", x"9616ba3b494c277b", x"049259583840ffe7", x"c9059c4f556e1d20", x"9c4e75d1521af5e5", x"78217fdf29452c43", x"d612ca272764fdee", x"9bb638e0e7713c56");
            when 9890881 => data <= (x"1484d5e7f9fd98c3", x"342c67696580edf3", x"cbf3ec2c2dfdcc19", x"1f77c5df80b5bd0b", x"513cac489d56aaeb", x"935ee4b937e922bf", x"f429310edf3c7c93", x"e8e39fe47134750b");
            when 7155923 => data <= (x"1d10c5ffd0f05e0d", x"1cdd7a7afc7dadc8", x"59823eeab47f6125", x"dd8810bbe14bb6dc", x"aacef3fa44f4672c", x"b725dfc06d762511", x"2df9fc95f478f5f5", x"2f68dae76ca7893a");
            when 23540992 => data <= (x"8710cc3564c87fd3", x"1e2cc056f276f8f0", x"0cdef85ca1c6c330", x"c3895c59a134078d", x"2b09ef4588d3c729", x"d0a812986a7a562b", x"9a1e4a05366301aa", x"43fef9ba0510dea2");
            when 1563641 => data <= (x"d8dc1732fda17e68", x"d04f31f52cc0f866", x"78ae0150bd3d8476", x"de8c20b0043d7ae0", x"9af90be9750d8971", x"ccbc416fbd1fe21d", x"5a343ba2c891d6c2", x"96824c28eaa1a692");
            when 22300283 => data <= (x"1325c537404a5db0", x"443975dba99685fc", x"f2bc6a65d9bb0e96", x"ecd7541ae40cdbda", x"c42954f57a3bc673", x"5e38407d97386b48", x"c87150476b92e6bb", x"b96650df455be45a");
            when 23640043 => data <= (x"546e5fa1ac6be1ca", x"3640874d995e6957", x"45e368deb5b914c8", x"c0f3039efd9b1111", x"6f7179d2b6449dbf", x"2cea2cf2a30d8533", x"dc42aae3940c0574", x"408093a8da93227d");
            when 6550477 => data <= (x"4e2139f5510d3ac8", x"d7b64d1c91869474", x"bab1da01b71317b1", x"f431c41c41a1aaaa", x"7b792ff9b70baaa1", x"a36085d4a2f8bec8", x"403449e0dfb88569", x"e719b8d441ded1e5");
            when 10045915 => data <= (x"5c6726c7088bf55f", x"7ee6b5945b36d405", x"2ef28bf4334e4c93", x"ba3101d8d235f772", x"fdfbcccf8abae34a", x"893df87bf55a317e", x"b24a4799c22baae5", x"206e605c40b4af0c");
            when 17673448 => data <= (x"cfb4b8af768665e2", x"23aa6eb223bdd3fb", x"ab35c698276239da", x"14cd6de1f46063a1", x"445fb5d460cc432a", x"5e5bcfd461026479", x"3020aed9bd2ee0dc", x"04c5fd9e3d022aa7");
            when 24077360 => data <= (x"b7e001d67626c92a", x"97de302e9b293cdc", x"0d0c9bf710cd33ac", x"856d79b636b76673", x"b1a0348cbfd87d95", x"4da3f01139a144ee", x"bab98ce61f5a212b", x"aab55a969b2622ce");
            when 541761 => data <= (x"b879a3e381205cef", x"6cd2ede2ca86737a", x"c1d690d6bdeefa73", x"d6838895c7f33d87", x"6c871faeae753905", x"b84b75748e10296a", x"732d42ed43276e58", x"0b1531230d5e23a2");
            when 16124171 => data <= (x"f68c200d5ddf3eff", x"39fcfd4a623c0f75", x"1c391a32df0b1f21", x"6984bbd00d41944c", x"98cb7a1d58c679e2", x"30e198e3b5313983", x"24c52298cc2c93f0", x"261f4563d411a5c2");
            when 32338198 => data <= (x"a3aef25fdfb9a9c0", x"7924eda2bfadacc7", x"cce28971f4a9b7bf", x"17832f8c3ac91359", x"5a580a841bab511e", x"c6c2fbad553cf5cb", x"c14487ac81b54733", x"f16ac6db4c05a290");
            when 16017020 => data <= (x"ef18a1b25d6a9a2d", x"394f42784973dd50", x"967b3e90fc0934df", x"895de90ad1fb6d3f", x"566a77a16ee8b082", x"d3c4ea0c5e1e939b", x"c4fbd16aafe783d1", x"d7ca1900e66d98d9");
            when 14265143 => data <= (x"b9d87e87fb43ca5e", x"c4161fdcc37ca17d", x"caca6ab9ba3ce0e0", x"38e1250dbcebc985", x"dcbb5b2083420e02", x"e127ce91aa56e31e", x"8b0e99fdd681e188", x"d0d637721a89ad64");
            when 27931394 => data <= (x"70f9fede594c6d43", x"a23e32c63afe5cf2", x"a89e1b372349a93d", x"b590495336d30cce", x"1d27115be53ca9fc", x"41094acca58b2f4c", x"4bc26ccd44c6460e", x"69e071b69c141821");
            when 32195946 => data <= (x"efd232dd15efe23d", x"b68fce2eb504370d", x"6cf61537e9cb17ea", x"5b41b6c7d824fecb", x"1b3de267a1b41065", x"c8ed62a1e565b29c", x"9ddb08141adf6573", x"240fe723cf15603d");
            when 23988092 => data <= (x"f63bf3ce2efacf2b", x"bf81ac4e8ab81c4d", x"ac8c9cdf4df92cfc", x"2c1bca6d23d7e9d3", x"361772bb32ef7e88", x"3b0ce56f7ba3085e", x"a364d28fa9a39ec1", x"1cb1817a90cccb57");
            when 4345287 => data <= (x"4235ece20465ee5d", x"2505d8cfd9831246", x"53e1bdfb8ab00808", x"86da83870de8e829", x"6ca256d312745f7a", x"39c18be9dbb8c578", x"7a4fb5565ba26522", x"e53c3eef7090b729");
            when 19611906 => data <= (x"f490d29b49ba8866", x"101ce63c37dd27e7", x"df2da99edc9676ac", x"d314dcb9a9899812", x"587a2be7d40ae738", x"4c1acb74718d126e", x"b577d94fde7f4f17", x"f077474fa927177d");
            when 11035068 => data <= (x"3e754727608c9072", x"3fe953fc704112a4", x"85869c2400c2369b", x"276a1fe00155b17a", x"0bb5adb9c37c346e", x"926e2e3b226e3625", x"1daf8522d5cfbd6f", x"22de1c348f1754fe");
            when 24703571 => data <= (x"382ac204ac2cfa22", x"039638f704f05c22", x"8ea8a36725d45fda", x"04ddd554ebdb4ccd", x"b6eafbee2338f81a", x"6035d0c03ca9c135", x"dabca71994eb573f", x"4495400d6af20161");
            when 7205042 => data <= (x"3276f61a05318e0c", x"3ba301dd3ae123df", x"b21c2c7af201aa4c", x"f475a339a8972afe", x"911549956ba1616f", x"fb714261c152fbfe", x"b54231f24e763931", x"d0478905fa34f0fb");
            when 26449342 => data <= (x"3a07d59a535db877", x"6e4995d0f161a9f4", x"44c28adb31cac7d0", x"0fb5185dd4e89a47", x"708f4bac31658cde", x"4382c112e7da9d6a", x"0d8f095d7361f363", x"b9415d7b49f26265");
            when 13831141 => data <= (x"c2f3b2394725714c", x"395d35c109eb2b1e", x"c5e39afc8469d94b", x"e7fbd56b85761940", x"7ce49d6d91146926", x"3108507024162057", x"984400fbda0ca425", x"6e8b40dd067675a5");
            when 24319596 => data <= (x"8fc0fe01d7ff2e33", x"c064c218e6bb501b", x"2c1ba8af98f1e912", x"3f9defa04ef73724", x"725ed29b814d4967", x"2ee63664c5c61339", x"e9c9b136a8349d7a", x"8f7115625ab3706e");
            when 30461005 => data <= (x"6ffe60bc7bd61168", x"8232bc0175c4c090", x"312f457e3aa37a11", x"171027b6dad8ca5e", x"9fc22f391715f622", x"6228c4226a6d54de", x"8dbb84294659af5b", x"a8f876082f6ea05f");
            when 33335191 => data <= (x"0441a99339cbc161", x"13600464707782e3", x"f017622af8e8636c", x"bc81ed6c6ccf061e", x"3db75ce77e6f9869", x"a28f49e36fc8250f", x"099947307cec5058", x"040ad76fc69718db");
            when 3325672 => data <= (x"0d8d0ae9c6790404", x"5401e6db563b9c64", x"17978161034ef5fa", x"a57be2ee285b7762", x"0084c1c70f543221", x"d863e44bb7d93954", x"08ab1fe4d56a74e5", x"fd4e2376415ff49d");
            when 9152929 => data <= (x"43f2f9df90ff8e8a", x"89a55a4804fc1438", x"d1d546c2a706189c", x"a5f18dc296809ca7", x"649753c99dfc47d4", x"b1694f64994b5ada", x"413c6804f065bc45", x"43f34a250b6df81c");
            when 24352954 => data <= (x"d1b0c10c79447311", x"d235915d258f9b5a", x"5631492a20002302", x"e34450d658d20a4e", x"c293f938a4857c46", x"85a1ad011e561e55", x"1f8d4854f413779e", x"7f0e5a5c87ea8fa7");
            when 17080286 => data <= (x"f03cd40166934b37", x"95ac7fcb572d8286", x"9d1ebecb051f928e", x"b734cb06f8d6235d", x"86fb43c903d63b5b", x"33128515bf95d4d7", x"29aba910538794b4", x"9a445bdbfcceb487");
            when 6169028 => data <= (x"40b7b271ec17b57c", x"f0ce64aad7d28a4b", x"25848295c4f9f9b0", x"75689b8a1f8b46f4", x"9f6afc18e204ae9d", x"8bb092a9d4db6e61", x"8e2089577a5d47e7", x"bd4209dafe53ddfb");
            when 9433940 => data <= (x"ce360218953c9e19", x"e6f846974efb8af3", x"d4180764c7a75be7", x"d41ba7e64718dacf", x"8bfd13703df5fb3e", x"c4776149dc41d56e", x"754ff9a12ac7cb26", x"1420841216240b62");
            when 10825689 => data <= (x"c416d0a40dfe3416", x"5ab27ee1b1cad87d", x"4843cb94c59c188f", x"83ed855d6293cd0f", x"f5ea1171d4a926af", x"9e7bf1907e730b8d", x"50b749acf6cb0095", x"d9aee930e95c7cdf");
            when 16861339 => data <= (x"010b56bebc54a191", x"012c00fea981d046", x"f5e6e3609c849dcb", x"f08598db10e55a42", x"4bfcb23d66cd7091", x"1468f71963f92d9c", x"d976dfa5dbdaf2b3", x"88c3ebccf8982d7a");
            when 17017200 => data <= (x"830f39fcdb4668c5", x"a66d9f05c49e3233", x"36be35b41b5ec647", x"6401958f69e002f5", x"504e5d08df46917c", x"644ca9595ab608fe", x"e415a25f14b3fbca", x"074b91b7d1511f48");
            when 16567904 => data <= (x"d145c68024775f52", x"de99357e3e9ba5dd", x"ecd2a639041e5d6b", x"bee43d6c44cb6b71", x"0d882f1a5fbaad40", x"72158138c8e6597f", x"85eb798a2e5b8f6a", x"53bab2286fa208c0");
            when 9741045 => data <= (x"20a4cf63be275623", x"a686e4a33da644f1", x"133d8728d5f140f7", x"7a6aee78455d94d9", x"5911a33a6bb5de44", x"ed7b33420fa6ea94", x"617cf2db104189cb", x"ee5ad702314980ba");
            when 18896818 => data <= (x"d8616ac4d562600a", x"215da036ee8dc93b", x"bb9c087aae893464", x"bc7f01ea6bc9c31f", x"17d2fde30df4586d", x"0f2728aaed0fe742", x"2c35b7273a644100", x"242a8f42ecc7081d");
            when 32084762 => data <= (x"e52ff13b75eca57b", x"70c610042e430e0b", x"52291395e5bdfead", x"9a2dda40e90e0a13", x"ff96217872a8b21b", x"afa17dd49d8b49ce", x"e98936c5bf2954f8", x"e7b6a4194f22eb07");
            when 3673207 => data <= (x"0b331453acc24106", x"1fdff08086de2d2e", x"7cedc32e4fa316d0", x"ad6b952b61659c16", x"5aac93941ba975b3", x"63b172de78626ff6", x"79e02ba66fd1b964", x"91d9ad4b7533b2a1");
            when 33761126 => data <= (x"6cb6512e4ab1be81", x"f3607d8f1d47ec8a", x"d3650a3300f4687d", x"c87046c5ea43c290", x"4b71c7a44c5182f3", x"43908edac0fc4452", x"5e897fcda2b90f0e", x"a21a1c15d4d0f14c");
            when 20488887 => data <= (x"87359485a298f6da", x"adf70567baa7e0e2", x"8942ba297a552e99", x"cf3520484127920e", x"e3af6576d928fde5", x"d08fd114736b04e4", x"63b2cc4574b49343", x"8db53f28a255add9");
            when 23798251 => data <= (x"a85218d6c27936b3", x"c488f03ab09c774c", x"8fef7a8cdc3d410b", x"a030207d892bb53b", x"f9d0db1b23491369", x"d2ecddb7b3ce4d62", x"f009580bd6e4d0d2", x"e4fe30cadf271e7d");
            when 22253139 => data <= (x"529d1696693d8109", x"bd6568ce0371b3de", x"591b0f077981921c", x"fab91dd2a3f0741c", x"adcd1a871c875035", x"84581fc948a3899a", x"758995608813b34a", x"996273dddd6e4519");
            when 1783897 => data <= (x"6be6fbe4b7a2c2c7", x"b1d58708d64cd158", x"e01f80f02d5b854c", x"0b7e884eeb66f4d3", x"03c8184fc9287dcc", x"0676dcdd5aba4471", x"e8a33096e6255855", x"60e19f568948c6f2");
            when 20984125 => data <= (x"d55c94f554db2dd9", x"d339eedf7c917fee", x"ee8ca6471656fdc1", x"a92c313ac7310da4", x"6614bd5fbaf49fbb", x"6d015700a20edb08", x"a2b261a612da6c05", x"ade7f33470ad35b7");
            when 18201345 => data <= (x"6470a2010c826b1b", x"9e0c129e2af7e2fe", x"3d74f76d9b0cb9c0", x"4bab99da32f8973d", x"8cb55f3e3fcd9cf6", x"ddd593e0c817e1b0", x"657b8a7327fe8c01", x"3eea17628a3d4790");
            when 29125084 => data <= (x"046762df034c757b", x"dca7a1ab2d5dd6d3", x"63fa686c99c58121", x"a362909fc17e86a3", x"cc633aa6f0b093ba", x"b5df61033a47a50f", x"8da6560ef8e36248", x"4b142f54f6022d61");
            when 18894771 => data <= (x"572cb7b92027e998", x"e061a69fab56b08b", x"8205a8ddc666a364", x"4af3242a2b9a2012", x"47fc6aeb1aa2495d", x"b15bca33ae1f05aa", x"f4379c4885f6ce2a", x"410779d82ebdaf02");
            when 22564387 => data <= (x"96370b082df55d64", x"643608bb208e58a1", x"4d6e4691e7df5463", x"f34e13548ae1fb15", x"9c1e6368a7bdad1a", x"1859b58759334572", x"08f28c5dbad94eb5", x"d52d3aff5f7c0b65");
            when 29260908 => data <= (x"803eedc6930d2a3f", x"4f3b7e05f53aae22", x"e422fd5364112e5d", x"8ca53e4aa58330e6", x"46adc8f9b31aeb7a", x"041d824bfe985fd2", x"7ce6f12805bcaab7", x"229309679ef050aa");
            when 28151428 => data <= (x"528abd0aa310af27", x"c93cac0fa19e4846", x"cbd41ad57463cbc3", x"3b5c701536a8643d", x"03abddcf3f5611d4", x"8a44f90356633129", x"0d0650af29b7ea71", x"a3c7d11dba941f00");
            when 19692884 => data <= (x"7c6dab9f46340949", x"d58c0f10682dd835", x"6199419a9501ef1f", x"6027389dcaa2cec3", x"110a687e3228faf4", x"c679a69cfc2c9a2a", x"ffec109f80b91f35", x"d77cdadd4092910e");
            when 30200589 => data <= (x"41c337afa52e2772", x"19832ef9e37dbef0", x"d864d032d5ab433a", x"36cf22b583a02ffd", x"71be9fa877147b0b", x"dde09770bc8bc5b7", x"bf9b34f9c6379500", x"6a2be526241a09d6");
            when 2307768 => data <= (x"0149a611e21fd1b3", x"70ffc21a1a438c12", x"d8978fe1278268aa", x"f84eb949e452d464", x"96afb432f3df54b7", x"f1e4bef36c528f8c", x"0a41b2b8efaa7cb7", x"60eaaa6f58e1595e");
            when 5568727 => data <= (x"57dcae46216db6a9", x"5dc2eb9379be172f", x"0f9c52d8048feae3", x"c944c19d9ca08a49", x"2912ffb3e99b1a05", x"d76bf20f428efa77", x"b626db1761f3a282", x"8064fbf5f0ebac0b");
            when 11578640 => data <= (x"44b1512573c3ace8", x"3adf78f7dc0ff2d2", x"e0fd65782e1d9381", x"6912fea32ac4726e", x"6552e927e3cfb767", x"972f273d0d92dd3c", x"32f3add9595dc185", x"cce311e1d2cec364");
            when 19345291 => data <= (x"6b8e8864a51ddc2c", x"10f96256d1e0d02a", x"23fceb73fd2461a4", x"ba6252a673822253", x"7512b654998336be", x"75adba943825504e", x"af4f8d1b31e237d8", x"84c388d0f9d3d3c1");
            when 16572332 => data <= (x"2a53acb660605ddf", x"989aede2b88dfa27", x"94be4daafd5a7ad9", x"f5443f39e1a93c1d", x"f8ac07b3e149f4a8", x"554b2821532153c9", x"d5fc47b1f8ea3a65", x"fe96af1bd6c51152");
            when 4814073 => data <= (x"92e637bbd270a830", x"6d0f213de05b5352", x"f86c49d2c24b3f4a", x"dec6bc669ff74755", x"fea5bb729059a200", x"ca40d73f2eda6805", x"aead78add0b85be0", x"838c7b78f11ea331");
            when 32703919 => data <= (x"f9bacc0b988c423d", x"6f8b5f1272157aaa", x"2cfb5f2b079c8ad3", x"2ba1b25b27f43da7", x"042e03b01d43fed2", x"2cfb674372856cf2", x"2cef9c58bbb388c5", x"9f308137d10a6182");
            when 22523404 => data <= (x"b6969d590573ddc2", x"292191aa5d4301c6", x"01b0346b2a842a50", x"681ce6aabe7e83c7", x"fe80cfddee233f4a", x"5b54ee7bf7f6bc66", x"db2dd815b7733af1", x"14204ff9edc4929a");
            when 8902096 => data <= (x"25a4936654d6ad32", x"322b866780c64c96", x"a69e2f59e4a3a6b0", x"9b1ca78c45a7753f", x"72bce82b51bf0f17", x"23e803094ddb4f9a", x"5b49f628f0bdea1f", x"4540a8a63bf84ff6");
            when 16332155 => data <= (x"a9fa451b99c254a9", x"4cecfc3e4911c54d", x"875fca9283140e43", x"5f204963fe913a5a", x"50aa433fada97349", x"00c1cb47b252681e", x"cae8eeb1b06eca82", x"cd533d2bfa38d176");
            when 17786457 => data <= (x"a8af449e827b3f8b", x"6e6471cfb35979e3", x"7488063e70593e71", x"8634d78df3bd1ad4", x"d97e4048daec6efc", x"f0f7089915f4c9d8", x"6388fd14c6259f76", x"6e7efc5c71422ec4");
            when 20899240 => data <= (x"c9121f0686daadf1", x"6934854015ebbe3d", x"b8e00d8d983d0315", x"2bb56eec79c589f2", x"2c24d7dd320acdb2", x"8da2ce3c76d9bb32", x"2182d9bd4650fc39", x"64fff0648df0d9e0");
            when 11538048 => data <= (x"dc21b6dfccc43a76", x"6741be23da863c7f", x"8b511ee119c5ddb4", x"2dd8c081702fc388", x"b708bc6b0530bd7d", x"fb727c07aa740744", x"4d72409a15bdfe9a", x"67ac6efac965849a");
            when 21392278 => data <= (x"5579450e78186c52", x"9f8c5602802aee52", x"4b82b36936041cb0", x"011e9096239e496c", x"6632f8eec6c34938", x"1e2f64091f7e014a", x"aa6fdb3b5cc9254d", x"715d2c798aa21403");
            when 23712384 => data <= (x"685edfefca851149", x"1f5c4c3b899a3cb3", x"742ed3d79b419a1e", x"033cab4faea7d716", x"fe50f4f85e3e60cc", x"5ae074183913fe33", x"e917cc2b4181c5b7", x"e53156b3d03ce36f");
            when 11169961 => data <= (x"5d9048320536ef6d", x"9a60cb202e09bc1b", x"48d4e4f73fe93fa2", x"01c51d280aa6db29", x"bce1d5f05a9026a1", x"867f006bd5eb42b0", x"838e2c718002f1f6", x"f8fd6b570c943636");
            when 33341164 => data <= (x"6fab5cec85378ddd", x"d5e2aae47f8ad612", x"92ef7ffb159d3074", x"897f2728d081097c", x"b43fa99f71319b7c", x"92ac59f88a851301", x"c5c659becee35243", x"72f44554f709c802");
            when 24776569 => data <= (x"45c20bfa0ddf4284", x"65aba2a2f2d6b0bc", x"90de879091ed6436", x"c773d878ca211322", x"8efcc4252108fb79", x"b5c027e70f00b06c", x"0ebe8294074531d6", x"f2df6313f1ef23ed");
            when 3947974 => data <= (x"e25fe85bfd0437c8", x"3e1d2165676ec5e3", x"f44365b025852151", x"6ba06f6a62c8b0de", x"035382985d74f258", x"054c235d44868592", x"6bb8a9d47018c65f", x"3d7f2292215c7e26");
            when 25668082 => data <= (x"6d670d731c64e629", x"424b6a18f38e4b0c", x"26554c27b1393547", x"4799c3f8d2ad7890", x"910226b8f87e6ca8", x"0e14cc476487f9b1", x"5683dcb60582bc15", x"1739a69bef5d115a");
            when 27577125 => data <= (x"571a07199fefd565", x"f6f5c7594c7985f7", x"02219c1cb56634c1", x"85f6e8367e8b870b", x"578b9c05846d23b7", x"fee59ea67ac25aa0", x"0fe479eebbbb4488", x"95bfde78734ec047");
            when 24007351 => data <= (x"3d449bb8982c2696", x"439655a9921ad430", x"eb9427fd42e1e6e4", x"97d776536959f3f3", x"0905edcc39fd65af", x"b6f4c3b68d71f5ff", x"b4ab26b2313cd1eb", x"8de47b1a468c6661");
            when 33689117 => data <= (x"d9904093a361055a", x"970b3ea22f0c2bc2", x"2bb377bd373dd38f", x"3e09d1b12c59de8e", x"fae432fda148f02b", x"81937efd29f9ba50", x"df111137dd6a875d", x"f52d299a4c280c18");
            when 1033355 => data <= (x"c5d5c92e6688188c", x"3cca0ec18faec1d7", x"26b59420bec75204", x"3fe1aa149ff8d6f0", x"faf2379d0b230381", x"da7bee72bfb9593a", x"307ba6cbfdc720f9", x"835ac72ab9476e75");
            when 3039519 => data <= (x"05da17ed83230083", x"630dfcc7dc4e3b54", x"bd4594943e5835ba", x"38c55a4191c0e6da", x"adf3193bb83787f6", x"ecf7f7e27e5ec3e4", x"9083fde3ee99439a", x"38a47a834eca5575");
            when 16194435 => data <= (x"134df7beeaa99cbd", x"2d5f0cb6053e09c3", x"50db58f6651d5a99", x"ba8265e2e70e8845", x"bc3df59ae7123fbd", x"addf5a6a3a571450", x"a012dba212241cb2", x"486ec81b2b0ff518");
            when 13541333 => data <= (x"707b20c99f723cb7", x"ee78b597145c2b31", x"e4b0f96fa298c8cf", x"3b6ddae6f207705b", x"db40edef6e505b80", x"d59d573dfafcdd36", x"2c3c69bdae58ee91", x"6541b2f9d8509d51");
            when 28206344 => data <= (x"7d0fd4164be291a4", x"674de69277b0e5bd", x"db9b465db492d73f", x"9cad4b629bf5e110", x"d1f8b060e70eba28", x"4c318f90f4d7a730", x"02b659fb9ccc2dd6", x"33b51ae9bc1c5c98");
            when 26363167 => data <= (x"5d5657836e20733d", x"63af2de4140693a4", x"e57bb1ff50a88553", x"48801fc3cd248cfe", x"615c06460867f323", x"967be8b5d8eed85a", x"deed0eeaa130186b", x"cd51c7644cf93a53");
            when 3775887 => data <= (x"728965ab18ac2ccf", x"d54149eb1a251cf5", x"ff41404237d1e53f", x"fb2994d488d4d80c", x"c60c85e3cbca2e48", x"560bd316c6676e47", x"d29aa75bb2b5e1fc", x"920cf241047fdd7a");
            when 6744277 => data <= (x"49280d72559ab6b5", x"a12287e3089b4afd", x"defe242f99152c1d", x"f0be21ab0ddd1ec7", x"e5992ce8421ac002", x"c06241368e241d6a", x"bb47af9d00510a60", x"d85bcac015c51dfc");
            when 14438974 => data <= (x"0ade800a57f7d49e", x"3f81462339ea5a9c", x"e6e91dcd4d28a516", x"7b74f9d38aaddd7d", x"2bb6e6806a2a67c5", x"64c9f58b9b105a82", x"632f1a8193a7636a", x"08ada1a0afcc7ffb");
            when 10509611 => data <= (x"56626089e4ba093e", x"cf2dc42a94bfe8bb", x"35d117af18065209", x"93fbccfece035e74", x"98fa0190291601a0", x"613d8c916959467d", x"fd9bc7bde143da13", x"d4060a96c4db29f8");
            when 20530692 => data <= (x"457c0e4d19905873", x"884fcb38d31479df", x"5d6e370b05f7c2e2", x"cb19ed859c76bf4a", x"c5c838fef51eaaaa", x"ceaed4c36afe7159", x"ee42908078368825", x"255c9d2d4454c1a2");
            when 18478586 => data <= (x"b1dd80017cae5b7b", x"0d42ebda9c6f3e45", x"1fcc82347497ab8d", x"11667458c847f440", x"04379a1ba6f35e47", x"4d3c7cdb92c6b848", x"86cb0360930e5d37", x"560d0aeebdd947c5");
            when 12477585 => data <= (x"df7b0a77daabcfbb", x"76976b3ae63d4315", x"c4f99452cc4b7951", x"208ecf2fa1537fc5", x"044981632b27f8ff", x"288640f2c8cc2906", x"669618e11dff3667", x"d8c817174d75497e");
            when 30152692 => data <= (x"7861aeb2c5dfa6ab", x"90d13d87d8981c73", x"b74dde9c924415ab", x"80db7f1f29ed58b6", x"6322aa70356ed2d4", x"8356c8b202a81088", x"45f9f4b3d24e8b4d", x"ef6daf47a46f1740");
            when 5215552 => data <= (x"f4b87e61ac319cb5", x"c6704b03f2b3b415", x"7eba89b1e0e8bd6c", x"05243d92ebea0836", x"6ace8852fed739da", x"a78542265c0580a3", x"d98965916bd8dc2f", x"e5b8a88c2750c49b");
            when 26679246 => data <= (x"682601ff3057cb48", x"7c5bd56292921c9c", x"1c19ddaf6c482ad5", x"b3af5a6cb02fb5e7", x"00dc12bad7563f6c", x"c3e6f20932f7b1d2", x"4bedd1b9d9f79f3e", x"09b74293671f7342");
            when 1211030 => data <= (x"0680e438ce45786b", x"07bd5f559ef34e05", x"13b000976556fc25", x"70c097dcb54a5382", x"290495e849a0f22d", x"27bcbcf05012f9f4", x"f0e8b93bdd858e5f", x"aea74d7d1b7fe790");
            when 23290999 => data <= (x"d81e0277c65542b4", x"06e82b4b15e5a933", x"e9ed15a61c90376c", x"fdc8b0d287d29ef8", x"c6395237a24dc0cd", x"eafd83ee7900d8d6", x"d5dc7162302591ca", x"caf6ba7648f99ada");
            when 22258040 => data <= (x"e8de290b3a2b808d", x"224b696340e4a6ab", x"cbfd03ebacfed122", x"960e127f6672a5b6", x"7ab87a5d31e7140f", x"3e49bbca047d24ff", x"aeb0a937871b5c55", x"b896778eefb2e688");
            when 27822120 => data <= (x"43f7e5795ba2a2c2", x"8b1009508fabb38a", x"17eaf00174148452", x"3920e1be27101b81", x"6fbb8641f9f3798e", x"f78776a3e4c68023", x"f63e00474a348966", x"ddee8c42b6da8de0");
            when 17260223 => data <= (x"f4044a24f31eb03d", x"0399c65f85b8647a", x"4bb7e56015056485", x"369da348e2b08973", x"5ea551c99431cca5", x"a40c403bec0a19f0", x"91d429c3ad1a0064", x"777761ed4d5ef8c3");
            when 5531254 => data <= (x"197e48eb59a44c5c", x"d0068f0c5929f050", x"c798c03236fe9e7c", x"e923a806a97b0609", x"a50290855cb88b66", x"387ccea389f66233", x"026d3fc1ab0a6b7d", x"5ae545cafa035b4b");
            when 23632977 => data <= (x"502ddc33c0b6e052", x"689172cc668eb948", x"b812fa5b1573cd14", x"718af0028d8957c4", x"c43072f679617fb5", x"63dff45fc0849431", x"8604fd7abec4dfb4", x"8faf2e666f221d0c");
            when 24055954 => data <= (x"91793ab22c6a983e", x"8bab2c2621252eb0", x"87eef8e0fb58c077", x"724e847b0d18cea4", x"1ce6abc10d67a63b", x"f65713c7ffa823bd", x"e386f28ed9d3a7ca", x"d76b0bc74d592655");
            when 21213185 => data <= (x"42e4b9b50b47df70", x"19867c3c7d9c7713", x"fa0d5d11e9551928", x"be0fa76c6a47614c", x"3a0c9d939cfe153c", x"fd19516b9c7abe06", x"c5d0ac75fc2ecc76", x"72dd91dabe5f0337");
            when 32234938 => data <= (x"5970bc928335469b", x"6a920e72ee53989d", x"33682dc512cece81", x"92b617945ed267ce", x"7c6aeffcfba95274", x"cfe69f69262157ab", x"3d15d5a34953237f", x"814359137206c264");
            when 3203009 => data <= (x"f0ac82c871987477", x"1d7cefa63bc251ca", x"f24c8e54a20017e5", x"b41d2e07c2351acf", x"8f3f02f207f6789c", x"bafe1fd7053a716d", x"d8211411cbc79335", x"fae90f309c7d6e1f");
            when 1393229 => data <= (x"63607fcb2d17a718", x"071597e1787be03f", x"2e1d79f1634d2f60", x"0f6e0d8d10d7f047", x"d5004d13705f394c", x"4288bf7203408f00", x"8dc1a40d7ac46ec7", x"40e7e08840cee932");
            when 491631 => data <= (x"9d4885269872eef0", x"73d4ae653c503b06", x"191df7a2ddb28f45", x"ff700676f157d79c", x"ec647f599ad107d1", x"ccc062e0c4f0f213", x"cc754e8df2fe62f2", x"e0fbe32d5af1d8b3");
            when 23172516 => data <= (x"4562aa0eb898d6ae", x"8a8b174e216cef4c", x"40f78bcba391fc7d", x"22a9ecad7c23e923", x"183a32ed5c1a6f77", x"51f6d171e4f80b9b", x"54ec35fb0caeb8a4", x"241f1695ca8021a3");
            when 8195387 => data <= (x"f84a843df19a8dbe", x"c68ecf3d49ab54f1", x"65b418e0bb08e01a", x"68b8b457f04239d1", x"b8bec54bb23ca76d", x"43ca4c4ad57eb799", x"ce79c6d387e2954c", x"2eb6b82439d8c03b");
            when 20391289 => data <= (x"abba1c283820c14d", x"6bd5d3211ca6d6ac", x"a48c5fe021704ec7", x"5a37d68549d3e301", x"e4151ff25f869cf7", x"743947e31efe2600", x"e51e2eaf2aba028e", x"c639de4377c23404");
            when 26450176 => data <= (x"9bb0a28935ff56fb", x"c7d3fd04ef578b3c", x"92d3e137cd839f8e", x"796f9ecd8bec10b6", x"4e6988673a200b5a", x"800082752b1650c9", x"aca2234d0467da0e", x"a343c08a9b64bb0b");
            when 9311532 => data <= (x"8ab7f51ae2ac128a", x"ffba987165a91ae3", x"ef2c6d21b547182c", x"5ea574389969cdf9", x"f8f5f367fa876d32", x"db93d4c80b06a6e1", x"54646dad21b34b70", x"944e534c37fd52ef");
            when 26581490 => data <= (x"807f61f674a63538", x"ee64b609272256e5", x"a8713d7452bce6de", x"1a50f3a15209c715", x"cc990804c429a22b", x"31368f67b69825b4", x"162f88234354c33a", x"b1a7579c5b13c29d");
            when 10219841 => data <= (x"7b2422625ce26bb8", x"2e392a7c56c3fc79", x"05f3190b8e7b31e7", x"a8b596c757105102", x"dfc3ce36a4eaacba", x"03985f40cf696a7b", x"6231d95b7e090429", x"b275d809b30af00e");
            when 18347909 => data <= (x"027bf40cea143812", x"dfb510e9f30a498c", x"5247eaed79de63ec", x"726d8640216d123b", x"e09ffcb3ce2b77c4", x"5194bbf3cf5f9bc4", x"a7abc8e48ba0d903", x"bac5a48248330432");
            when 21990101 => data <= (x"4116746bc1b15773", x"e7fdbd9568d0e736", x"b1d2a9a0a5066580", x"6bdf22da09018e25", x"750ac08b4fe0faa0", x"118ee488527aaa70", x"433e1e4b8c9715a2", x"7acbbf07aebb53e6");
            when 18495228 => data <= (x"137f6ed1551b3b65", x"551f937c3569155a", x"9273cbe017d60a6a", x"89c065bdc64b0915", x"a194782781ab3fe6", x"1dbd5ed64b7c70b7", x"7330e09bbc76cd66", x"2fa431bc07a37682");
            when 20181319 => data <= (x"80eae2f69a83ebbb", x"a5d5ded593d41271", x"ca580bd5f72f6343", x"ab18e15622af9204", x"fc9b624182fc64d9", x"410bd964ecef7f13", x"b364ef4d5fa7e9ac", x"03bc1baff11ae327");
            when 30834793 => data <= (x"3b373abfc68263fe", x"21010c855e85bcae", x"969b60555e6aca43", x"29b0002bb8266e57", x"7cd4b29bb3c42f84", x"8933f8e9347592b1", x"9e630b6ec2d93905", x"9e4411a0f81fb3b9");
            when 27992791 => data <= (x"0c4e8d8f109f2523", x"40bd867246909a17", x"54262e530cf3bc72", x"9f8e938d4d06e651", x"74652098ff9d23c1", x"de95851caf79d40e", x"24957ac82a9425fb", x"339a4c2f396d8d7e");
            when 31493112 => data <= (x"e90cefe61a8cd050", x"7fe7cdbe4d416687", x"08efae5eeba34ffb", x"f722e329dd1a188a", x"65799c142cbe82db", x"b8d0b4f033ffe4b9", x"4266859b30348a43", x"2555932938b0752a");
            when 26950585 => data <= (x"48de9aeae8e9ef77", x"80ac75ab3de38a4e", x"dce6a07b2b9b2cf7", x"efc2d5df71d69092", x"7e3f0b597571c2f8", x"7da8cdddd877c92d", x"b1651aa8c4a57f20", x"6830f94ee34f2198");
            when 15671387 => data <= (x"32e00cfeabf9208c", x"9529a00e8961f087", x"acedaa55a518e867", x"129d1e74c248a6a9", x"04c4d53b370c7213", x"e6181decdc564674", x"b2842a666f08416c", x"a16a6732b8ebe876");
            when 22773511 => data <= (x"62450f0231f62fd2", x"d0243ac1cabf5b28", x"1652ffbe36f6d716", x"525d9b7594358b07", x"1a14c019e5a36f6b", x"1f1f37f82651aa77", x"71e21fc31e0d5917", x"b213ab2addeb0ac2");
            when 31236855 => data <= (x"039601004bf2a750", x"f7c3e5f7bb6ea943", x"17a3fe5342f3e863", x"5a1da98a6a1a0e1c", x"9b9843cb0861e913", x"391acad64ff33c16", x"cac16754685b19db", x"aa915bed4bbe88d1");
            when 27104663 => data <= (x"7143479131e65494", x"8fc03586f66ffa12", x"f5204fd74d90f9f8", x"ed0de1b51a4f889e", x"8a3aef30b37af588", x"862039d6940bc9ea", x"132f6b56573a9a07", x"6a82b72eaa2bba33");
            when 7037279 => data <= (x"4aec683b099943bd", x"a6647b65b2de3242", x"9c83349df34be6da", x"928070cbe15e2b03", x"e7b156026dd7e948", x"6d97a0432367faae", x"ff2f8317807de115", x"20b071046088f505");
            when 25707586 => data <= (x"4eb9078d1b147375", x"2c9610c46c7e862f", x"442111bfc94f77b2", x"a7acd258609c948f", x"83c92aa2f31a82ee", x"f4ed4beaa0b185e6", x"d6dee18ff560154c", x"3ed9187fca00ec1b");
            when 15841115 => data <= (x"b0adddc6271f178e", x"ee8c1f375d7bd19b", x"fe58eedb6ab520da", x"53738d9273d5a71c", x"87ab90e99ecfd6ec", x"25025ce26f662f7e", x"96e0e0f71d1a33a5", x"779b74953bcacf1b");
            when 1671087 => data <= (x"7914fd4f51168120", x"4e1dfdfbba909b59", x"d4cc20f3d6be2a58", x"7eb55d45f9c33ac6", x"4c37f4f3c91df23f", x"c2230d19c62b517d", x"00b588121c08e646", x"90791407a508ead9");
            when 20227539 => data <= (x"084de6d08043310d", x"e8c8b31ddc9f2228", x"b7d55f7a169750be", x"ab54d3c2f0109f8d", x"bc8b6333217b6bef", x"a103543f42119765", x"9b9bffa491876fbc", x"97f69e67aa0a05e6");
            when 14956042 => data <= (x"8ec03bf87ce9197b", x"cded754fb1fab61b", x"8066cad27a940119", x"2079ca705e44a910", x"453a30428f5294b9", x"ec0fb95e881d7da5", x"bbe4beee84f241d2", x"e85b1883ce523e6b");
            when 27807625 => data <= (x"7a731d4c26db589d", x"130c26bf773ed93f", x"2ea980285a6399eb", x"a8356578f4e792bb", x"e76003639d2c81bb", x"c4f14199366deb4f", x"07601e336bfaa11a", x"6581256947732ce3");
            when 14963719 => data <= (x"0a5cf7b6716ae231", x"2db074d60c090a02", x"19d76a471a61d126", x"56340326ef373bfa", x"f71d0f957537c2e7", x"6dda73660e557f07", x"62c60b2d000522e8", x"602c907c5402ef18");
            when 24903017 => data <= (x"7d0ef958f16700b2", x"7692f5f189738396", x"eaa0679fe5912500", x"4a2bbb2096205fe2", x"adbec6ba06bd9c6c", x"617161019f13028e", x"783ffed4f04b0252", x"d027dca1c3d94d1d");
            when 1349049 => data <= (x"91262a0e2d63051e", x"a7f9f3d3e756e92d", x"a2131fd73d05d1b9", x"32105e4587c6999f", x"efd9f63c5b499510", x"60048e688d8b0903", x"f4b9ac131233d55a", x"ce75091142c10fa9");
            when 10872854 => data <= (x"b0333cc0cdf65f57", x"560966241fffab98", x"53a11396984a0c7a", x"a78dff588e688445", x"b643881523a8f8ec", x"f1d4018e60be0b97", x"833c61755274e30c", x"c47d69dff55f514f");
            when 19864675 => data <= (x"177042ca3096e69c", x"de9aaddce0c30f6b", x"4c03e275e3941c08", x"6957be74326da635", x"e39e9600a0090317", x"8cd9663913bdf234", x"7bbe43643bca4de1", x"36e3f382a8f21d40");
            when 24710037 => data <= (x"c0937f56a1831703", x"9e668c317dd420a5", x"62f6eabaacb228b0", x"f72d23b755393fa7", x"200b89a33f9a086a", x"23ae81969e9098d3", x"fa5e737399ae560f", x"8ea4594af851e148");
            when 33805632 => data <= (x"dfc2e7397748f001", x"48c04056dc4c12fe", x"c8a4c6048e31f842", x"be08b777e500a4da", x"935bbd1343d84de0", x"037bf7ebb959f1a7", x"cdef1552a600b547", x"37476434b494e8cb");
            when 22044342 => data <= (x"384d63821b30fdaa", x"cb05c795f41ca30b", x"d1ae281ba571f2ac", x"5b9dd11709b36f51", x"e06f6e5990d07e84", x"62e0e4a219df58b4", x"52114e77fd3c2aa1", x"9160fabaf4ab8673");
            when 4907460 => data <= (x"761c6cb9d347d0d0", x"cd995a67853764fb", x"467bb6f5ca2ab3b9", x"8b75bc29d4bf5a2b", x"93fa6967d8e952cd", x"c3588faa559b6bc1", x"77fb856827f8c4ad", x"b9e7122ade642d2c");
            when 8710974 => data <= (x"119875a9aead219e", x"0bd8f8cec0d3dcd2", x"347686d2c99a50fd", x"549778e4f0600491", x"b3186e3a7a0ba438", x"31843cf19f33499b", x"6d1e383133818585", x"12a1120e2102dd38");
            when 3550981 => data <= (x"0ca3a7e9f67bd5fe", x"35acbed9ba628871", x"38023b55277b9070", x"0b428cefd3344a2b", x"43354b7118a86fe7", x"7e00de6239de17e8", x"4e9b87ce3dbf7810", x"ba6aeb9ea9f6b5d1");
            when 12145773 => data <= (x"2ad11577b62b3bb7", x"f54f15c6532ffec6", x"938a160e759dfd91", x"00d2af5f15a51cb2", x"d44c84967ec89d47", x"a20a7f0fb54f38ca", x"c45bfe87b61a4ff2", x"16aa34f8df5a5940");
            when 15701599 => data <= (x"c959829e63de9c2f", x"6634f67553d05783", x"c4af0d7a02d7f6f9", x"86a7d94493261fe1", x"5595a7bae87ef366", x"528b70b17f8055c4", x"f5e2b39ff31d7ea3", x"3f89fae0fe4c800e");
            when 33820583 => data <= (x"2ab27243278e3fc5", x"e1c669e05eeccc5e", x"338fc32a5fccee94", x"9e653e91a4dec77e", x"9531d8a0903525e3", x"184503605fa3a390", x"ef953d1d4812739b", x"7d90ffc6312da8e9");
            when 6845488 => data <= (x"f5c41d7608500b6e", x"9b6fa39f4578a544", x"46344269ab7eda25", x"f8b743cf8c59b07a", x"72d1db868af3f10d", x"c786ead7f7135509", x"5f31f2b49c7321c2", x"fc08c728703dbe46");
            when 15470528 => data <= (x"402f7041043c344d", x"21235e4822f3f778", x"182bd26153c191d8", x"3ee44d63205357a9", x"b8abdc3f2cd0ce36", x"22b0a258763dfddc", x"b1ec0140ef9b857d", x"8fd8ee97e689d5a3");
            when 12604483 => data <= (x"0c004ea8f843f26b", x"3c71dbd5bc486f5a", x"8bd06f69b32b74ce", x"421768241c74fcf8", x"a21b6b36e931107e", x"0442eabd15e45a85", x"adafde234e735274", x"3ed29892d2584335");
            when 1475068 => data <= (x"a110966627db6ba2", x"8ecca1f30e51136a", x"c358e153f4f1ab47", x"5e8ab2982ae8aeb9", x"ec26b668847faedb", x"77bbd7ee5db997d8", x"be7c0397c4524699", x"a4d28022691d9d41");
            when 20778729 => data <= (x"292c4dae5e195c85", x"39e6237ed67f5daa", x"640486d411a95835", x"0a6bd783df23146c", x"32f8b1c431ab9e02", x"0bed195214485d8e", x"cfb998514713b4eb", x"d0e133d0fc309730");
            when 22637981 => data <= (x"48a25bc3eb8dfbd8", x"5ee532bcc58e4225", x"44d4ebac997d3eb2", x"4358f954dda14dd2", x"fea480b1cf3d6e87", x"cd969328dde386e4", x"d0225ac011e59798", x"7bd65e2eed16389b");
            when 16187637 => data <= (x"d1e920f052ae245a", x"d57438540019421e", x"61b1dfac60383ff6", x"2fe538a19eff9b83", x"ee87c674d9cc561e", x"3763b4048f6ee781", x"dc7ba27f2f4e3096", x"328b1b2534ee77f3");
            when 1384750 => data <= (x"c84c8f24b3e9825d", x"2897dd4ea96048e5", x"464a45da6c230cef", x"0ba1553b2c83869a", x"29c88ee53ea76385", x"376551842415edb9", x"fba756fc5ed49b04", x"e468884c0bd1c531");
            when 30654203 => data <= (x"6fe7a73f019b3c49", x"8ad51294f6289dd9", x"eab71b6bd52702d9", x"5ef6fe4ede1b91f5", x"97e31d5bddee7417", x"f72998a7e3bd9760", x"302a77c244d76bf8", x"0a0a8497b06ff912");
            when 18339545 => data <= (x"e923607be5a67f99", x"930461442dab9a9d", x"a41c85ad94f4c2a4", x"37411d3b4c60c07b", x"f5754214ecc4d721", x"93d07e3ffabc33ba", x"1bad889a65d7423d", x"55c8dd5d4460a1a0");
            when 23582472 => data <= (x"9fa469def12ed919", x"23a013933ae8606c", x"b4b1c0dc8a824c98", x"cb3dec391f5dd795", x"951ab7b69ca44e8d", x"c0015eef610fd603", x"8e6b4aaa393d0560", x"3f2b232e9e05a1eb");
            when 29916534 => data <= (x"e21b1fac65e2f0f6", x"6b5e8ebb8a41ff61", x"00ab83b91f2b99b7", x"745a54ef641670bb", x"4548815cbbee95fc", x"4a79c3dbdc5c823d", x"0858b20282fedc4d", x"6a8b60be2bb4475b");
            when 32004528 => data <= (x"9200a2442ac63e82", x"685f9b3c0b1080d4", x"a98103e123d651af", x"061fd739ad2c7a2d", x"4e3bd8d71f79b653", x"b71125fc4cb5828c", x"5fb14122db22aca0", x"c53e4321548394db");
            when 22929815 => data <= (x"6fc5a10f197a7bae", x"8d39b880d2a8bdf6", x"5f34e143f2fbc485", x"cb107e86e4c9cc8c", x"0fe75c29c090570d", x"50f5c457c30362ff", x"0e46a08013df7180", x"ee1028240a87e416");
            when 8546995 => data <= (x"bd5d4bc0a9246236", x"27b934bbfce6e116", x"e7ff389b74b15e3a", x"0a047c5cfb91fadc", x"a34b63ce6e04c518", x"f813740960cfeeee", x"225b2e51362b7605", x"13e2155dde9f5033");
            when 26175532 => data <= (x"897a8b1f0b46fa0c", x"7a3d3d331d652ed7", x"fd134bafca0549eb", x"d75787e7e08c0929", x"58c4532196045273", x"b913fdd9ce6bf1a7", x"6333abc857874830", x"1762117b29cb1002");
            when 7482302 => data <= (x"53ba64607e7356d7", x"7780628d3d93e860", x"30afdfbafce12de5", x"ed8ce5bd17997fc3", x"fa0694c1a98e45a5", x"9422cb8b4cadbfd6", x"6cccf3dcf0a963fc", x"839f5ce3ccc8052e");
            when 27869475 => data <= (x"9e074d45653fa468", x"86d5847317d48530", x"1be02501c165b7d8", x"170397a536450c0c", x"1b1810ba71be5bfd", x"ae0ff3ac9fc6b3b9", x"9fcc618ea4f4b6d1", x"fd70d06f5d0279b1");
            when 27437380 => data <= (x"ec8ae266817ac2d3", x"ff92d2c0c69132fa", x"70a3fecce700b6ac", x"98f78bf6be4d4540", x"b2855f90c5f1730b", x"2727935f4ad22314", x"b3b8f839767b575c", x"9467f37cd824f7a4");
            when 27341630 => data <= (x"c58ddcc9d134200c", x"045b73b2cde52e64", x"0fb918552d0f8484", x"234e396f331f6c95", x"8257f2c36e5b1c87", x"6d44c1d0fb356817", x"171c7da75733a75b", x"6b7d42003b767b33");
            when 30247303 => data <= (x"bd37332542e66fb9", x"6a09f18d177a44f8", x"10a3fd865de880c3", x"a8dcf4dc5bf3e6e6", x"ca3a6dd3cbc4c5d3", x"b18b9781bdc8d45b", x"8fc2d07b213ffe99", x"2c46173e4a69c3d7");
            when 10541674 => data <= (x"3a864fe3c91ea59a", x"5da6b3d9d0779313", x"c3d28206ff5b7b9d", x"1c96c317b6115a2f", x"6f0a242091ed50d5", x"dc5466aff8a96677", x"d5cd26248809c53a", x"28090c5c36636279");
            when 17833121 => data <= (x"cd1c1e5681efdc23", x"23dd4425a9a39de1", x"c359e43e7d533011", x"cc6fd8596cd64cd5", x"1484a97625b2db92", x"2a92eb3c71c55dc6", x"d21f46008ad95ef3", x"f208e26ba001caa1");
            when 23700020 => data <= (x"c95a20d5a6719fef", x"246cc3bf38b5dca6", x"0db0fa11958767d6", x"55d711f978564f24", x"7702888ec2adfbcb", x"f301ead0ec8d9b00", x"ea906c21827f5be6", x"2c9c4dc62f8ef076");
            when 13004679 => data <= (x"87defba79d9034db", x"1f935f7b8bb1324c", x"fe8dacac49539790", x"48666f5c76276c8f", x"231d0d5b5d060892", x"fa16a0576051cfac", x"b0da5d92054003aa", x"914680e20c0c3e51");
            when 32359220 => data <= (x"796f421531337e14", x"c9ff747376f7712c", x"04466d30d2c9de32", x"c3ec52becba290e3", x"87c4e1650b79dc1e", x"b6aedcdb16e423ba", x"bb36ae9460999d0b", x"532c759446149eb8");
            when 24819508 => data <= (x"5c217646d49613bb", x"6254abbcc86b2822", x"7ed4165f1a7049c9", x"8a8a286cf2754c9f", x"3d9b525a89edbe52", x"1451f440cd5f7c0f", x"c21d6d6b65452bf8", x"0a5610669cc03dda");
            when 20288840 => data <= (x"3cb05dec8ed0f680", x"f04b6311638f9ac8", x"6f30955f0cd07267", x"15c276ce1140ba51", x"1622ce573a27c1d2", x"c1a9758da756abe3", x"1544f614a6e0c099", x"d348475930a255bc");
            when 12913296 => data <= (x"f0d53625fd69623b", x"c3d34e82a496fbbc", x"41d1ff5172dce5a1", x"fc2e85eb7b0c38a3", x"fbf1df8547eaa310", x"f49268ee1ca0293a", x"67250e5941c811d5", x"0f6eb449dbae9fb2");
            when 13763304 => data <= (x"d2f6c2ad5461fef8", x"edc7685d0a77e47b", x"87913779b55543c9", x"16cf01617569004a", x"a3e159adb9b28370", x"b4f45e0c56f13e95", x"a53227650640afa4", x"ddcd450e4be3e77b");
            when 1901175 => data <= (x"0a8860a7db2ba193", x"d1381730ea47f1d9", x"d9372978a069b010", x"ed58f9dedd339000", x"6a209c5aade4133b", x"4aeb0ae553e413bd", x"d04551ceac881f1e", x"5bd1e65aacb7fdb9");
            when 26459702 => data <= (x"2b218de5673a4d77", x"d6412c95017be1fd", x"43039bb5597887ca", x"79ac6038bab81d50", x"c97e0ffdbc02b694", x"4fc7042cd2b44986", x"5485df8931c5c174", x"388aa98ecaabe6c9");
            when 32709903 => data <= (x"7af8b0a11f34bb65", x"017b022d528febb2", x"4a1f322dd3c6bb42", x"4c5ce0353185dd39", x"2cf1b7924e0382d9", x"351060383f880a30", x"9a74e5d95d738e93", x"de9a50ff327bcad4");
            when 20397764 => data <= (x"4b59e025bc3dcf85", x"4a3b29bbd796f247", x"3aec5e7c06806739", x"3300681cb638f464", x"edceadf1d8bf31f6", x"78b62eeb254c7fcd", x"94506fda2a34b10d", x"fae51a94daf1bde6");
            when 24897142 => data <= (x"23ea2c1345c5a0e8", x"a0cfebc2efdb0924", x"b726d4d86b823464", x"14769b5bcfe46eb8", x"58e84964542ac28c", x"a665244f396b815c", x"7b95b2298b27a323", x"4fda3ae8d02cd85c");
            when 11338393 => data <= (x"f61268a3f5c6faae", x"533d74d03717a76d", x"fe30a9ba5de36c5d", x"d1f3edc7a22b3dbf", x"8c8fc50086649e51", x"76bb84d80065859a", x"9007acd2af466b37", x"552483ef265f9d1e");
            when 3790920 => data <= (x"bff9dc9aae89d0e6", x"61492d0bd4566d2b", x"63ce9dbec8c33b8d", x"3656ed44ded0d5bc", x"6da498441ba9a36e", x"7e53f6d050f7db95", x"144f91efe542b439", x"20444b03dc0e8c78");
            when 29938966 => data <= (x"98907606d8519c08", x"4fbfe71a3bbb5ea7", x"4cdbdd1185a79afc", x"600b65953a93ec4e", x"4baa1d6d1a2e4591", x"29013a0ec334d4ce", x"9be48a0c0ad2221c", x"85c7d520ee471504");
            when 17922746 => data <= (x"1f0d6e18c1a381c1", x"b2048176dd4a69a8", x"d5bff264539951d0", x"34c364b198585fc3", x"326187fad5f9db94", x"66eb0e08e788ba2b", x"40417d00d3ba78ce", x"e53baf8065b2dd74");
            when 6281761 => data <= (x"6b1dc7bbb658d44b", x"57718c7936a22257", x"44030b65934d26f6", x"f4c89981fa72e76f", x"377470fbf71cc195", x"4519d40b01e6d31f", x"ff2e09bd3d8edcd7", x"17fb56be552bca7b");
            when 22886824 => data <= (x"d4166634bbd2f33f", x"0aa80e108eaa81ad", x"18ef559fbe7c2280", x"b35c7b9999e2f9e1", x"d21dd4599d586800", x"e55ee8cf066ef77d", x"371e3371fb16ae0a", x"3fbd035abf6d43f6");
            when 15348718 => data <= (x"4614da4de0f5c3d8", x"e3617480c9037696", x"8035d2ada9dfccfa", x"35ddbbbbcc514052", x"5a6339f95abbd664", x"b01907848f70159c", x"3ecd69f5feedcc5d", x"416320b7063ec8e9");
            when 14403818 => data <= (x"432f4ab7f46fcbbd", x"b18e52a8679080ae", x"d5d6763bc2723c6d", x"7f059a59cd44c274", x"522c66efc206ed17", x"79ec5f32cf2c4a2d", x"65b03f3c2b3c11c5", x"8180e0ad0d4af34b");
            when 31062777 => data <= (x"31f33a9dc7af87e0", x"f0244feefe2eb904", x"8b9f754601fcdbc5", x"66f2f3edb41f100b", x"044091d08adb9632", x"52abc2abf0fdabff", x"fc49f11277280d4a", x"4e7cb4d19e990f73");
            when 12539859 => data <= (x"14b7cccc60499fff", x"074894e6833f622a", x"79a9458b8ac2fc1d", x"f8216c15a6c6cfa4", x"7f9871018b2b7ca0", x"df35cf03ed70f310", x"8c05a4193e5b27b1", x"0ce318f8e90d532a");
            when 28292253 => data <= (x"98165ee07bb8e37b", x"f5f04a1153eebb21", x"8da1bc7a660ff371", x"0c9016499aa4e849", x"9cd45a43a91d97e3", x"4b7540cf1cdcee96", x"67318b58a1fc3d7d", x"d838d7266a99673f");
            when 30377946 => data <= (x"b5d2ed85aeda8972", x"6190e32fc0d44214", x"d365b924b3e7c2ff", x"b19c90ce452f8c8b", x"e8d0e3b23577e51f", x"2af8a706e44926e4", x"346a3f555004b79b", x"7b611f1e12c67021");
            when 6034735 => data <= (x"cce66573b345d275", x"7b4e981311e4f436", x"bbf87a3513cddf37", x"31c2f888ef3dbeb1", x"5f504609c947cf44", x"6f5bb66ae8a3b7a3", x"62bfcf822a574b20", x"0f47377c74da0241");
            when 26492829 => data <= (x"f19a7eeec15d696c", x"77c2879def953611", x"74cb9cbd33102c80", x"0146f1994c5ea626", x"aeba73e51d5315b8", x"46cd772a8991774a", x"db479e1310b7a0cf", x"7b5403ff8a34b34e");
            when 26287882 => data <= (x"777a121d01063264", x"9382084a27a6e56a", x"f4aed2c63d545027", x"3d5a5325822db3f0", x"b816dc16420bef52", x"f55bcf1ee6d88180", x"3f43d0bbe7b448fc", x"4e46415265dbac03");
            when 575108 => data <= (x"ecfa8b1df4bcab1d", x"53531f36d7ce9c9c", x"d7a4c3d73defb505", x"fc9d64c5432c3cae", x"7143615507e8febd", x"423a7b868ae0321d", x"83a4ecbdc8fe2926", x"17e475990616e7b2");
            when 16305814 => data <= (x"6128e23b4bb8e8bc", x"cd33846b21571668", x"f55cf2ab6575ed8a", x"621d05c9610726cb", x"32170d19aa2dd003", x"3a402f5ebab25d33", x"a4876f84346f4951", x"ce95e074aba9d798");
            when 14409121 => data <= (x"00f8efca512f366c", x"27f5e5f39b2139f8", x"00f6c0335f17d359", x"91a139c3a10c9d02", x"e62b158ecb992951", x"16fb94aebde9fe79", x"12ad3f2790ca42c0", x"c0a383e2bb69c87d");
            when 17229237 => data <= (x"ecf6c52fe12de273", x"abbde186d1519844", x"539e95654f289bec", x"6b7dc42e711dceb1", x"ea16eb0a2667f256", x"1823816a9c9cc1f2", x"d1a5aa22089c8205", x"ca0cc4382a0296a7");
            when 25055002 => data <= (x"700649f8cb335585", x"557083bb42c03214", x"b441f61aeccba3f7", x"69f2431dbb97ec74", x"b497ac5ff85907c7", x"a8b9938daa2db851", x"60c4c3ac19f30565", x"f8b3f16266313e81");
            when 24461623 => data <= (x"e8e2ab6f58b04552", x"e9fc30e79e099c61", x"b95245750778e322", x"78d9c1dd2666cdba", x"5a965f2ffb99b891", x"59e37dcbb7f0ab2e", x"f7041d95d8474f39", x"6e34a9dcd7d1f75c");
            when 16353753 => data <= (x"34bf7ffabe7108d2", x"d44b4fb47d7c0aa8", x"5fb149c719894648", x"0ccad882ecdecc8b", x"ba4e000eb349393c", x"91fa30409eaa1e26", x"7f85e06979856cdc", x"6ad1edcc59dc6abd");
            when 28287533 => data <= (x"af7401e2e466f2f7", x"7427ea4a7b1b8959", x"12efb61c11ac8088", x"e6f4895eaa59461e", x"92a3a1dd9af47819", x"bc102ebd0e9345fc", x"8b190ef2314ad4f3", x"191e534768c5573c");
            when 29922945 => data <= (x"9b04953944d00bdb", x"57734b2414c37bbc", x"6a14b4c62c329a05", x"7a937f421087eb96", x"5d59dd2d67768cac", x"1cdfdc1568ff85ad", x"8f6b15383ec676ef", x"64e200a7823136b5");
            when 18808543 => data <= (x"a6a819ba0e92b5f2", x"387a32643ad7d50b", x"60ba1d78b9f4f9e8", x"c1678b4501c36fdf", x"56724d0803a1d0ad", x"cffa2ced2225505e", x"acd64ba656be3bba", x"c9f760f018a6f222");
            when 22365738 => data <= (x"a6dacc44143f998d", x"06f3a0f565db58cf", x"81ea4d76fb97dee5", x"1ab32d809e0c67ff", x"eace61af6a4c46a5", x"c374902669dd5bfe", x"b9b0a5fa0b1063f5", x"349baa477b25f1ac");
            when 6762954 => data <= (x"3a98c6122c678228", x"6761bd0007ca6020", x"86351bac44d9282a", x"2ec1c7e2d1bd0d09", x"8e45147aa2e70833", x"6da1315cf9da79dd", x"9a769cc228b3b1be", x"6fdf992e7d69a421");
            when 20437709 => data <= (x"81d9e48e71aee3f9", x"8a9127b976406387", x"1c04cdba4cfc37ca", x"af32bcec72009927", x"f61a0373a40eb456", x"cc6acc7df3d8ab39", x"e9bec7b9eb33da14", x"ade5d1311863658a");
            when 24112365 => data <= (x"64e53ab2b57bb316", x"519c2b96e7bf1ef2", x"d4024d359e327562", x"82e9dbc1e94112d8", x"363aa56df8c46814", x"a76cf6698aae6f52", x"dda6fddf5ce7b799", x"289707c1da235ad4");
            when 12374279 => data <= (x"4fe802a5279fe917", x"d505fe47086ea1b7", x"f78643f61c0ee395", x"e88c56efe1393206", x"dead442d8f344398", x"7b4013730eb380a1", x"c62ef1be766dabdb", x"4c3a0b614f4bbce8");
            when 9186100 => data <= (x"77fd4495af4a28d2", x"ca8a9ceb9e2e638d", x"822239f3590f0e5b", x"59130f9bde209b44", x"42460745f2ebdaac", x"824b5c603da2b83c", x"db2f5d225f39df70", x"30bc2d694c733125");
            when 9204604 => data <= (x"2ef25c76e143d82e", x"9659db1a10ac1a16", x"ee87f5a42baaba0f", x"9cd61b6e5daf154e", x"f69eeaac02ecb0a1", x"3eef789ef3f16572", x"39688cafbb1dea1a", x"b1ce2ad4110d73c1");
            when 23527629 => data <= (x"16150a584bc983d0", x"cb82ac1119e03435", x"abf5fe88fc7c1831", x"c47724886ce7762a", x"3b6f36c3fae40619", x"a277ca71d5fcba26", x"79fbd9916f3dc2ac", x"181de0b986c58100");
            when 4367696 => data <= (x"11d654a48044fd5d", x"5904640bfbb6e4c7", x"493b3d822fae4f12", x"58ea0fc09244eff7", x"97bdc7d7fa137ec1", x"00e4eb4eb4f9f6d7", x"7ea01f78463da756", x"79d88bfeb963280f");
            when 15612889 => data <= (x"61775c033b7005a9", x"0b4361d0d88ed289", x"e594148921b5eca3", x"0e15fcc5bf051a5d", x"59dc9872aa84dc8e", x"6c343f40442c63dc", x"f9b72f3f7eb0b848", x"a08e10c68aeef199");
            when 11048653 => data <= (x"f7eed610c1e0ed76", x"611a0e7fc0a4d7da", x"c3bb1eb4c42feb0c", x"984876ced2933dcb", x"969c3a937bf1fad4", x"4315422fefcebbe6", x"a335d6e83da7fe44", x"a92725cafb080e5a");
            when 25478434 => data <= (x"926881c255256ce3", x"1469a97c0b1cc1b7", x"37cf8dd7ab39e3d8", x"1eecd6658286a0ba", x"dd54762e3cf1223f", x"e453722cdc357a1e", x"b3449232fee3dc6f", x"25754ce1cc940358");
            when 8989074 => data <= (x"039e9048b055df24", x"aa84cbb756a6810a", x"107efe706edb54ce", x"5636422410781f1e", x"f5c2dc8823a62c8f", x"6c1ac1f0b8988a8c", x"91c448a73869296c", x"7a204b0519939b65");
            when 5647714 => data <= (x"e308c03c6b469f4d", x"eefd4d91f09bc3dc", x"0d4abc612bf52f77", x"92790b92c66eff03", x"752fbf476e2a8273", x"bc337010d8b00f65", x"3be3fc7620fa5d5a", x"8e32570fedcef9cd");
            when 10329235 => data <= (x"edb1c94084f4d78c", x"ce98240588bf208a", x"e953f7dcefe7be69", x"1d97c930c264ff07", x"e8c5dc08e7ee189e", x"93e49897f6cef648", x"c0997a76d0dc73b2", x"4f2ff6824089cd44");
            when 27621841 => data <= (x"cf6d946834c96a62", x"1596f77770a14bd9", x"bbb785295a232d8f", x"47405ac46e1a05cc", x"aa56c3103edb4d1e", x"0700e56db6cc42c9", x"c633e8b0c16f3d81", x"15676520113c4763");
            when 7169677 => data <= (x"900b5a05a8f4c990", x"051844a51b468e02", x"3c1f87c17c0b9070", x"cc6b9946714168e9", x"fb1c0dc18eb369a5", x"1b31fc5b7f11ffc9", x"4b8fc7521880288c", x"aa4d188b90a16abe");
            when 14898435 => data <= (x"a1ff8e86851c4f8f", x"482cd436a47cae7f", x"468a995c3b4ab984", x"39602ff572c16812", x"ac80e98464cf6388", x"d5b011e7890224ed", x"c1a7504233698704", x"87f074a926170a9c");
            when 3847737 => data <= (x"60306479356fda64", x"e7e516b0130d1e2a", x"e4b3b4e4d22dbf40", x"e4aef23a639ad5c7", x"855c01c5108479b8", x"b7723bc6ba2359aa", x"0e3a59eb83534927", x"ec5de595fb3a5d29");
            when 21430326 => data <= (x"9e7fbcb881e25280", x"4c3a0fe9621691bb", x"4f995456366969a2", x"5fff2ea259abeba5", x"6bc8ff4188870f92", x"b84b9df3e676e70e", x"d57ebef4324088e3", x"8176fb099de75bb4");
            when 11114919 => data <= (x"7e4c4d134f55d461", x"b317a503df5b443d", x"d20157dd4c208bf1", x"cbe9203dfd5e15e2", x"0e65b50e737fa178", x"77656c7f26b477ea", x"075a738351ecbad9", x"ac9e30e3a03bf85d");
            when 13225438 => data <= (x"4d940feceadf73f2", x"8c579d25f112a569", x"748aaf1c5710a44f", x"2d199972388f3b75", x"57957a17eaa88bec", x"22a9fee5fa85663e", x"267da63cc82cb20b", x"c8e6e2454d51fca7");
            when 31725353 => data <= (x"bd35ffbe9f1b20ea", x"d8593b8862372ea6", x"3d5423f049017653", x"d06301c1c80645a0", x"bc0e9e5ed66e8215", x"1d8e7c7b7928d63a", x"ea26f0bcdf958339", x"cddb56535548ac84");
            when 12837838 => data <= (x"ad3206cbd8211eac", x"ae41e79b34963980", x"01c0025fd8479a2f", x"0e19b4e6520aa969", x"bcd25e656312d297", x"f9d80b92a7b777ee", x"25740d9d531b9163", x"c75a534949cb977c");
            when 24369061 => data <= (x"04f12bbf96dd4a23", x"e5536a169c3af33a", x"2abcf8b5f35bf138", x"5c19dfa1f180050f", x"85e562223b920671", x"aa8700f041cb06a5", x"a7d76944c57aea37", x"b4aa5753caca5fed");
            when 14296268 => data <= (x"909681704d786fb7", x"62cdd9f881bc2ad8", x"843a4e89df888a23", x"a5e09753bcff1ebe", x"f45a1315f611fef2", x"bc92dfd26eee6041", x"291bfe614c7e118f", x"d8e9d4433f084943");
            when 27767326 => data <= (x"8f2d4d01e4079930", x"e18fb896975b5bad", x"9f00a1acbb307cb6", x"ef0a3ad9d40f31ad", x"5c14b1c56b6bd6d3", x"914c6c2532b4e082", x"a35814c49138ab77", x"4a32d9cfd92c052c");
            when 29258515 => data <= (x"2e436bc65aa61b2c", x"c7964d73830d2337", x"6d1816ad8dd08061", x"15e9bf9319d477d6", x"d266a48bfa1eb3ec", x"a631731d2f70335b", x"372c83efcc4c4f41", x"85f9807b93380c68");
            when 4246351 => data <= (x"ee122174451204e3", x"fff8954c38bb9450", x"d35ba83b6d23c236", x"96800471ba2e776c", x"cbe09c1881d248b6", x"0959d82ea3fab291", x"19e2a889c21687f3", x"e70202be6b0de550");
            when 22644624 => data <= (x"a9bffdbd80d1e707", x"df64391cbb9714c0", x"bf9e71651a7c04a4", x"ebba784f7a2672d1", x"92b34eccb630a073", x"80d9b3bd00a0b97d", x"107f06b308e6930a", x"2fa8be5dd4ed4043");
            when 3578286 => data <= (x"e2aeb6e276f5d1c2", x"1e2943d4c99b8007", x"de2de5bf49f2423b", x"2dd539ef79ac7630", x"8f10295551007faf", x"8ba3f7639c4f2048", x"5cbc99e77abfe165", x"452225fe82d00431");
            when 15785491 => data <= (x"c8ba6c109ac4d4b5", x"625c9dc3a9808b21", x"6991112f19363e2b", x"45e26b4e54c0e76f", x"c6009e8a41bfb262", x"4317613ee1bb97d9", x"90d1c17fcb4b4740", x"f57a67c2d2b98dc9");
            when 25916775 => data <= (x"5994672b74d9ad6d", x"175899d0997416c8", x"4300446464f079d8", x"5fe9d5f933cb6d55", x"d20ed4b313fa1903", x"8a400a5e117f0ace", x"88e36091c3f31050", x"da43b7a6c399194a");
            when 4939430 => data <= (x"2f2cbccf2a00ab3e", x"df54aef4ca9e3a3a", x"d330b6d792f23805", x"8478e134aed8d0b3", x"77bb924e6e71bf9c", x"9215c1f744eff828", x"0cb9e478b0031a3b", x"fb7a59f619aefa09");
            when 22766131 => data <= (x"a024b1f7e8d8e0e6", x"76ee1c9241f82b44", x"aa9db37e7675f4ec", x"0db1e6c067718be6", x"25bf07d5defdba70", x"0844dc7dbca742f5", x"b07f30f149955b35", x"5e513778e299c828");
            when 30055612 => data <= (x"d0c9e08170b5ad22", x"79fc970613c3ab01", x"df719b9b79563619", x"f4836d436247871b", x"40828c4b18bc2bcc", x"9c62ea032d4d0041", x"62c5d142020c31e3", x"2516a44522797620");
            when 8826674 => data <= (x"6526519a840fbf87", x"6be7aac2a6f7ef0e", x"b02521cbc7757e31", x"84bb03bd53186213", x"460da2c46853990c", x"443cf015b615520f", x"bb312d38901c56ea", x"dc4101ba86397693");
            when 19947986 => data <= (x"d40c4afcda7f10eb", x"89f94226f3e34a70", x"9264ba0135cc17dd", x"c351755ac346660f", x"d925d2c0d53a903d", x"2d1e8b763ca03de4", x"c7801fc8902e983e", x"463ae7fc20692fc7");
            when 9870254 => data <= (x"ed7a33aaf288d103", x"bbd50634368597a5", x"e35dbbaa26121aca", x"d4231ef59cafd308", x"4776544ef8a9db0f", x"6e90dc2b3413d56f", x"3a3c217ee1e0111a", x"c28bd8afd7f0d714");
            when 31412212 => data <= (x"2bb44bc884d61751", x"5d09c9aa2f8c8c12", x"c936cae426cbc0eb", x"99e7b4ea6a86078f", x"42f997858e50c33a", x"2ef2c11c145a43f1", x"58d6b1459eb99f23", x"d46f7ea74ee3d1fc");
            when 33242773 => data <= (x"23ab2f5360f66d31", x"b6374a75043a1217", x"56b81beadfebacf3", x"3682a081b8ef22eb", x"b3c8ebe9149ea7c9", x"c796be2c6a727393", x"41fe9ab8185726cd", x"1c76fe9d5187c50f");
            when 3813504 => data <= (x"05c77a0727590c09", x"7643e1a1f49e74d4", x"ae16309753c8e883", x"e886e1fc301016bb", x"9a72188c6284e794", x"59b23cb1de89198f", x"a04f66fd1adc1a93", x"247c1b92ba5fbe6a");
            when 7491907 => data <= (x"d5bf0c45d79db619", x"c41d7ab253a3209a", x"b8bed16a73b78233", x"2fc49051f669eb1a", x"8035e09af71a37da", x"8e720eec110658aa", x"d458184dc33a7079", x"6bf820c4e6474a5f");
            when 32890018 => data <= (x"2cc4ddb76126ee20", x"2033dca70a76bcab", x"8f53447d6cbc6f3c", x"4445f3f735031923", x"b2e72bb2847f2e06", x"79a58cf13f0f2eb4", x"0c36e75cfb431888", x"01e720c89674b314");
            when 10539382 => data <= (x"b4730932e7d26981", x"e5e01d02a228240a", x"7bf8e5ac2d1e0d4d", x"734c5f24f70454b4", x"199332463e8eea3c", x"bb9ef8a4e60ed619", x"271233fd7cc0e54e", x"f49a36b827ed5266");
            when 24037533 => data <= (x"124f13a78a49168f", x"32a6757cd9744541", x"edf1b9b42336ba3b", x"90a9f59e20bd009e", x"27730346e4f805a9", x"b1fbc4fe34f88389", x"08eedf98c7ced1c4", x"4755df487704d439");
            when 3892703 => data <= (x"b6503b5a94b3d054", x"22cc430c3493660a", x"89ff8c0957da4a04", x"6043464b1daa3dc9", x"4c79cf9d911c6b1b", x"dda00e6d5e517f1f", x"ee23fda7e9120d4c", x"e758bf26ce5c740a");
            when 21241135 => data <= (x"65e8b800fbd105bd", x"e014ec3246521a07", x"b745afa9e319616e", x"6a285bd4e721166e", x"28aa6b96ba120957", x"02af6c1776faff17", x"155f40fa83619021", x"033a177b96da0f90");
            when 13031347 => data <= (x"84297ff8f94837e7", x"b91c8ad7b21f2c4b", x"45b76ffa28d3eb6c", x"abd92f1e98e5d549", x"922433cd70361a0f", x"4a3af767292baef6", x"e12775b6d9781e70", x"cdf1f3e76e55fb17");
            when 19540590 => data <= (x"7ddb45c4921a2324", x"cb2a65811fea19b5", x"460b4de1bc371555", x"bc0d2dfcdac033cf", x"59b0e51207420419", x"2d80932d7bb3126c", x"1d069abcfcbd8f97", x"6786ba04ef9e4127");
            when 25816126 => data <= (x"c3392e7394283f6b", x"a7251e072741bb6f", x"ad135434f51ea40a", x"fa7f83fe08fa17a9", x"1ecdc16261729885", x"2548c566a968258c", x"89ac9a1737f6ebab", x"33ea6fb6e47f06cb");
            when 2681675 => data <= (x"048871481a7396bc", x"aebbf878b0393b27", x"5fa11b5e2c1af548", x"9681f44b5ab76373", x"f98e87483372b71a", x"99d2ade9aa4ad3d9", x"518467744788bceb", x"4dee3c53eea12907");
            when 24939086 => data <= (x"b318333c45033907", x"53c7688aefae620c", x"2ce38abdc551fc45", x"019c4d396cdadc78", x"bd50d52c09d6d0ef", x"52fc9cee49f2072d", x"27161547f96e367b", x"52c73d0a7f044b7f");
            when 19064048 => data <= (x"ab2aacb00e01f955", x"571097f7086367d2", x"551f2035fdc685a0", x"86e53e79fa702b5b", x"5ba01e22b9162394", x"bb7f3211dcff0f3f", x"1f3904d5e4322b83", x"39e766bd25bc0f1c");
            when 33069682 => data <= (x"bab87f2798720269", x"0d02d4c9ed2d11a7", x"cc10b58545e19226", x"83d04cf76aa6252d", x"9e0fdac6954319f5", x"dd383ba63d588417", x"6b1887a03780b6c2", x"4fe9d71dbe016c38");
            when 19261214 => data <= (x"a4363e99340ce284", x"d067f000f8a874c6", x"63b9a1bb311b5e3d", x"18ea438ab634f611", x"3a792157650f45b9", x"a1d4d71f38aaa80f", x"cc723aa6d5cd0c03", x"d7eb20d9e4b93682");
            when 10285180 => data <= (x"3c0dff5d4d1dd184", x"960e2b79b07c40bb", x"4a29d10b3ec19f3c", x"44acedc2abe368a9", x"38c7f5d60db2efaa", x"c09e2e2575870080", x"86a9445f151ea50c", x"a377334622a0469c");
            when 11538185 => data <= (x"408eefdb5d085951", x"09740be98a65fc74", x"a092170319660e81", x"94f05187d045dc7d", x"60017794f92ad5ca", x"dd4c031ba7c66e32", x"9045fa8a28d723a6", x"a2a874c560659be8");
            when 13103898 => data <= (x"959ebd69679d9739", x"634948fc45b7d93e", x"8ed14742b2e89373", x"fa2eca1535f9458f", x"1f13cf9806efffe9", x"c1794cbf2a5e033d", x"e1644ad45cccb46e", x"67416e1a3b6a5047");
            when 21645838 => data <= (x"6474fa2c2de106b7", x"aba0f07029c43f97", x"b06b0d5a78537b54", x"084855eedab83c81", x"a568c7b9c0d8f1e4", x"f253803e4a44b3bc", x"ed4613cd48c95b53", x"7ec10a5323d65a66");
            when 21655392 => data <= (x"ab968a0a48ed14af", x"329e52610f3fdf25", x"f920ada2ac007d56", x"5dcec62de6d02a0f", x"a570b38ae3baa898", x"60c036baa3ff10cd", x"fb99aa98fa39de81", x"ea020b28b8df69c7");
            when 15751265 => data <= (x"7f81f6912786a747", x"4a2c683ced433689", x"b6717b319d7f3b85", x"83fa6e2fd6074b0a", x"5b996792535c176b", x"cb2098d4e26e5945", x"8b73c3bf402872f9", x"9594cea350911e60");
            when 33067772 => data <= (x"501dab489485ca78", x"6fae43d189309d62", x"a4f94d5e7f226192", x"e44b19e2b22b3233", x"9ca5124f4ddc1c71", x"70ba6f475eac7c6f", x"5118dbc59d68f3bb", x"681757ca87300eb9");
            when 22398350 => data <= (x"165d221b755c4967", x"c15f6a1f33050ab4", x"5e92c9e21f8728fd", x"76409540f169b65d", x"c6fe63e5f14cfc84", x"1588e6d3eb2aeb5a", x"82999bb5b4a35d20", x"12f38826666a946b");
            when 22226138 => data <= (x"f6e03d108cb423c0", x"b8818f1c9b9b042f", x"9489e638af6fe0f8", x"33cdb7b59c02f06b", x"e759d716e2143777", x"84a4639e1674f984", x"377f41de3dbd8ac6", x"e648a4d44fc8126e");
            when 11763959 => data <= (x"b54721ce461e930f", x"a8ce9cff6f4db8ce", x"2cd96ad3d3215dba", x"7d0937f5eddedd19", x"5355c58ea172c8e5", x"68a99482c9119fa2", x"0d14b7a1d9fa5a57", x"5cf18a05b526e7f3");
            when 27257286 => data <= (x"16f01bfd544f3b95", x"ccd2a3eccca33109", x"f9a2b61092069a8a", x"33f060790303fd31", x"9e681c0046e59b19", x"689abd338d6d1935", x"c87e29a4425d73c9", x"8888aa09f0feb8c6");
            when 20347124 => data <= (x"21e6982f9f7744c8", x"aa68546f569e9d98", x"f148c04293bf8016", x"11036ec724d7d608", x"96bd6e5986b3983c", x"246bf9cfbc5acbec", x"2131e9229c474286", x"fa010630abc28234");
            when 3655589 => data <= (x"f57824455aff9126", x"0f85770310a441f9", x"84d49a688f0f9225", x"9df8373df3f968d2", x"994a00da8d0fb723", x"966eea9181e3a683", x"f53ff6d3c21f1428", x"599653a1f1232bbd");
            when 15537753 => data <= (x"70358513dff276ea", x"cdc22adea281065a", x"350042b0614bb978", x"0ee06bd35e3ff6bd", x"5b56e32069e73d4c", x"219e02298f907269", x"5312ad8b2e63d195", x"19414342c2a40372");
            when 25296315 => data <= (x"2d7208318438a1fc", x"4d326d74d20bae75", x"d13dae9578ab4c95", x"26e4dfcdfcaa918e", x"62137d6dd31cbee6", x"bc9caa904d679113", x"67c1ed95120566c1", x"aa4bd59a7769cfe9");
            when 22103895 => data <= (x"491587bef579a632", x"7567dd694c33e677", x"37d245cfaee1b5e7", x"2d60ef6914ae6836", x"4bf9d918773c4d1a", x"2b46adfe2924de30", x"a369eb1a5c5ac57c", x"2522894685809447");
            when 21538964 => data <= (x"4a499ae90cae0c48", x"5bc33d9564e8f3b3", x"7fe802bcd9d8dfa5", x"b0fcfb727d20dc96", x"b92e630846595a98", x"1cf78f082b3cf967", x"f86b79670e846cce", x"f08b1d071f2a9f78");
            when 4831058 => data <= (x"81e3ce281e4a693c", x"10b39b352961e169", x"9fff064b4b785d9b", x"519f7ec38ab827de", x"9a46861c15ab3220", x"a5e01a9ebba0059d", x"877a02702641813b", x"956777fc2f70c954");
            when 28987286 => data <= (x"d6739c0130e98605", x"46353a047bcc746f", x"7126f150d73b488f", x"e5e54d29edc6cb85", x"74b56953d40625c4", x"dfe2aff4daf3693e", x"56ab38664708a74c", x"533b9b2aa80357f9");
            when 5207160 => data <= (x"b4fc24110634cb68", x"a355cb770f9b2732", x"9ae1fd21a94ddda8", x"7c087f7ddf471704", x"37e0c0f5adb0c6bb", x"1dd587e5dbe2603a", x"24ee25f71abecf81", x"945f53919f0e1798");
            when 20668921 => data <= (x"8b7dfadc8e84c730", x"1d97d46cdf9a72ad", x"94e7cee4a34c0096", x"136eae1b398b08f0", x"19bf2e3075416f0a", x"9b23704fa31952d6", x"d21328675badc9ee", x"acf642837e51d81f");
            when 17232587 => data <= (x"74cb786a923460e6", x"73f0867c50d3bfaf", x"037f3d193bb13af1", x"8e04abf7b9884a4e", x"635dd99cc87cb09d", x"206c04f9cd5bc1c2", x"653dbeb371469163", x"c9b06f5b9d320915");
            when 21984535 => data <= (x"2774acbbc3343f43", x"3bd9e2a3b271228b", x"848f2be8fe9cb950", x"e6783d601e1fe1d4", x"72abf557bf8bc52c", x"d34acd847257ee24", x"c8b9320a8440aea8", x"2551110435d18bd3");
            when 8926706 => data <= (x"9e24c7292dc631bd", x"e4ab7b33c2e6c6ab", x"b16ff763e6de41fd", x"06669c35f351115d", x"f65be7abbb5aa791", x"babdb27b96611e30", x"d7ebcd92ff0f7a91", x"38bda20a323d0141");
            when 24643334 => data <= (x"535c0ae6fc9ca3b4", x"9b4aac9408e4b788", x"b87482201e0e5ad7", x"cc38a79be456adaa", x"3f88aef70ef4115e", x"c7bddf54410c8e8d", x"2afb059e62ef03b7", x"325db84da4ca42b7");
            when 14491155 => data <= (x"b0a0f47004607066", x"ee5e2f0a1cdd6d82", x"7b16c339cf9b280e", x"ad27f32a2768cc7f", x"9c1c5a8014da3c84", x"a3baa03f5d206314", x"c798fa191dde45cf", x"1432e9387e284df3");
            when 1750127 => data <= (x"683f6bf9c5023dbb", x"a04a109e14d669c4", x"c4ee6691dd1e0a3b", x"9fff9c20707745a8", x"dcb768198a9c47d5", x"37358b0cf0e5647b", x"e97e2c847e39934e", x"6b4c629b0942399c");
            when 31110770 => data <= (x"d09c264dbd07cb95", x"df3902a5f706a7ba", x"ce2d772f40833adb", x"4807d649a7b4b408", x"b01de62e59862783", x"920fd6a339657c9d", x"7fbe3006d83414e8", x"a0b61aac9ebcab3c");
            when 23636630 => data <= (x"3cd52f5b72275c45", x"37ed932e7106c2de", x"527bdb46c5cddd55", x"f06619c8df51ba50", x"ff47fab38a0c21a8", x"66d422496576e023", x"e4e766588e90708a", x"21d81d5f1d6c8142");
            when 21461607 => data <= (x"d8596c54472bda8f", x"a2a8b06fd2f30521", x"e4862baba90bc1ab", x"29ade51801dec422", x"c4174955de92e079", x"d86f54d5a44b3edf", x"fee6f0671a4df9dc", x"5ce82716d7da6d22");
            when 5912238 => data <= (x"94b2edfc25526f45", x"97d97cd7e636cbf0", x"c68ca03073fafc27", x"e11f9f0b241c7d3a", x"83a9c352bef7d912", x"affa2344a44a5408", x"fa76279532a782c7", x"8fd93fdf0a3595e4");
            when 25979983 => data <= (x"4011db6556b8a782", x"6904a3f20e697c7a", x"f3e8fd1f62274255", x"ef3f9cc7b3d26d8f", x"b2abd837aaabdec4", x"93d41722b74ea77a", x"20bb69c72b0d3d64", x"a44b64fcf7c34cc1");
            when 17933671 => data <= (x"503c6d763d08b7e7", x"574f5431180ae039", x"cf14702064e52998", x"064281e4cb94fe6b", x"268ffc60e200ddc9", x"a804aae12caac805", x"6c124ff37d1c5beb", x"2b1a9b55139d67c7");
            when 1104278 => data <= (x"bb7d68757d93d8fc", x"88f50e774473fa5f", x"59bd1c7456b3b985", x"07fbc6f1f925eb97", x"f8b2350ab65e5e83", x"d919d7934b8302c4", x"e014a5519dcaf472", x"8172f1a85b609b5b");
            when 824793 => data <= (x"1842326f976c196c", x"23675c6c6c5c24be", x"9661d75dfa67174c", x"a75516edb487da46", x"edc2252698b98916", x"f00e23720e91a470", x"b7ec76af5fccd3b4", x"58a895222f7a7ece");
            when 20825707 => data <= (x"cbbb38375b77ca67", x"15c0d02b4e82acc4", x"205f5c6041615e1d", x"3fc338048541047a", x"12ae5f0e039ed333", x"76327b0bace14715", x"4d8acad44081d9ee", x"de8623ce2055a2fc");
            when 7816438 => data <= (x"fcdf927ee214c75f", x"375fa4caba569bed", x"1e71fbe97c650493", x"bc2bae8f77cbaffb", x"27e39d5b41e445be", x"e6653aec22ae1efc", x"779982eaca2aecb6", x"8962bc67b7ad9fbc");
            when 2479370 => data <= (x"810016bf7d999cf6", x"5e419aa6df05285f", x"be115dfdd8bda82c", x"d9fa32953ddaccd7", x"0ac1cecfade71949", x"629c88dd7ade5566", x"0db0ee3697fe9109", x"2ee7369f23f48cc2");
            when 11715045 => data <= (x"7a21aa207c068a51", x"283b82531bf037be", x"3a60df36058e8c73", x"aa2fd3fec27f55b3", x"fd2aff8991284012", x"e9f1fd8747c613bc", x"a12b83323ca83242", x"755460f2470d589c");
            when 2525394 => data <= (x"2e7f81cf84acfab0", x"3b7dec61bdead8ec", x"39a5f2beb095734e", x"f4a6b3168e324d24", x"a1c922fc97704679", x"d613196574fff6e8", x"489eb35c1aa172f8", x"92ad49df454c2bbd");
            when 17720489 => data <= (x"68d30aff458552b3", x"bbe67560c6de975e", x"1f7c209a56c43df5", x"9db76267cf260149", x"caa6116d3712c5bc", x"c1ae5ba859bd7d31", x"672a52fb08042146", x"2129399285eaee28");
            when 33447162 => data <= (x"63325b1fd8292470", x"f58fe05cfef27650", x"b5c161a42a081239", x"c1a520250bf4e09d", x"9386209ea986e28d", x"1fab7211d1efa9cc", x"f4430d55236d0154", x"2a8c070fb9dc4db5");
            when 13392197 => data <= (x"dd29c6a81b889fc9", x"274b200736be94e6", x"d09a859246e9b03b", x"c9ef292fd9424cbe", x"65a6f80fde07e997", x"156f4ee57fd0bdad", x"3742ca7ea60351a3", x"62ee93b489ee0df3");
            when 13641333 => data <= (x"457e57ef3d3bfa3c", x"5da600514855edc7", x"1c8b89df9207f7c9", x"b326b2bc16f5b41c", x"23c506f9d10c5da1", x"10227419f91adf6a", x"eebc39e8f666fb88", x"43e4f7c2ec195d9f");
            when 25901530 => data <= (x"5081e2526772ecb8", x"7d0291e2e1b1381d", x"2b59f801dedc9205", x"9f3a83e75b4c611e", x"98b90d74e4b52405", x"b2bb2931b43d9153", x"9bd763f4e72aa415", x"e0d326cde7154fb3");
            when 3321633 => data <= (x"7315504f99057f61", x"82d9df95d77d3966", x"c0279445b14e62cc", x"3d9107e5de083a55", x"b549d02bb0a1dca9", x"0645fd92c7692b79", x"e0ed9e65722b11ae", x"40a6923e3fde887a");
            when 4846415 => data <= (x"5fda8372f310e9b0", x"18ec5abb5f43ec4d", x"4a649242a639a94e", x"ac9f7acf4d6d4ac1", x"65dd131f97c909bf", x"1f47d73a5b0c573f", x"73385819fdec6967", x"c4f17ad380616b8a");
            when 21164778 => data <= (x"235ebc0d3f2d9d14", x"8e54e645fb272834", x"dd0b867a404a527f", x"c8f854b79cef76d1", x"4381279d590a9531", x"da8ebc3317e0b528", x"1cb4c0e4ef1f77dc", x"efbab39793b7de91");
            when 12533866 => data <= (x"48e18a6bb30dd4ac", x"461e688ac969c7e2", x"798cc9f9e52d48b5", x"b691623ae610a04b", x"d1975357c47cb772", x"070d8285d827602d", x"5656b4683776eaef", x"794164822fbc8e82");
            when 7413823 => data <= (x"3b57ebac3eff16c2", x"93b48a63184b0599", x"0a0a283751b36969", x"3ed63ee64e67f200", x"46341150ad8d2287", x"253b98ed5ae277ca", x"e4407c34c26ee30f", x"f9361aba8a4249ea");
            when 10134630 => data <= (x"c0ca12c3daa7d751", x"6725ec8e27504c5c", x"9ccd6101f6231a25", x"dcf4c2a193e71b06", x"43d1610219b3236a", x"21e8ab67478074af", x"591fc414a791b172", x"46707a6fcf8b8d07");
            when 25641175 => data <= (x"2bda2f3db9f25d6e", x"a4bdaef1732ea280", x"cdf83565e308dbed", x"7ac7b3e6bb69ead4", x"31870103800f6758", x"ce3b98ec68e29063", x"ca7b6c5a3537dfdd", x"f1801c93bfa6ddb2");
            when 30076428 => data <= (x"4446cfe8a1d1a43e", x"1d953f6791f97741", x"bf5bf4596d7f6735", x"92c9c61f324f1d1c", x"188a8925d78b5e03", x"fd6c8aa28f67ad68", x"6c92889f28edc795", x"561a3387e695a7a4");
            when 2704217 => data <= (x"81c37198a5668e1a", x"4502ff5326e8f6b9", x"5b3f38e1721dca80", x"688d85a9eb717f8b", x"1300bbbb1ab45f46", x"574e6a65c5767c46", x"ddb647a9e5a14eec", x"91cf9c149b79a1c3");
            when 23384472 => data <= (x"06c9b42d74e9de69", x"fe115b330fb51dc6", x"27c79ce553841477", x"5bec73da8a79b501", x"633eaf9eb34bc41e", x"e266af8f833c2bc9", x"297031ba699dfbef", x"b3223d160997b792");
            when 25421838 => data <= (x"b56409dfd4b6a3c4", x"ebf2e1e029ac9baf", x"3f2af39e6f9102cc", x"59b92d145d8a845e", x"d8de5e61403c5920", x"b4e0f35fee927463", x"e33a13f38b8eb196", x"549dfc3dbc5f10f5");
            when 24859968 => data <= (x"2cb5b4a2a44d8be0", x"4441fa07b18f88b1", x"5e17002963dd0220", x"83828d952c2c3dea", x"cfe8ee46668b23cc", x"75e187814cd2a8ec", x"0f93b930ec5f064c", x"76cb74083c3f27b3");
            when 24947971 => data <= (x"b0e71fecdb9e294a", x"aa6c75a56eaa5e8c", x"a6c49edcde4cc673", x"228c33940deb1c52", x"c753414ee6d322bf", x"6e79dba65ecfc4b4", x"0f712f03fb776bb1", x"6ded59b0923061ea");
            when 24160332 => data <= (x"c53f2740b4491077", x"98e1aedda9ba0b2b", x"b36d8b439b1552b1", x"eb87da4cf164a8ee", x"b05eff676d5704a3", x"09f6e08f25af6026", x"0ee56fb09a491dab", x"23aad8ccb289d97f");
            when 15190824 => data <= (x"c259c47e2cd88efc", x"4a2db153258e1d79", x"b16cd6cfc7a9e87f", x"59d2d63ef64ec12e", x"6c66ec0dc8a28713", x"625d0219eb1eb022", x"3be41181c7dd0c4d", x"0b53550f8065d48b");
            when 31546125 => data <= (x"d8b3648c1d2fd0f8", x"5ea3bb37ba3ca724", x"90ca23f1b91fbaa4", x"9ef7c3c8a34eb63b", x"e0032cb4b622c1b7", x"9dd6b61f60584f64", x"d3906e1a02a5ea88", x"972e63a737efbd1d");
            when 26432377 => data <= (x"54fe308b25661773", x"42732d7f2cf0ea2a", x"45fcc618a3ca2529", x"f8f6f691d29be7d2", x"a2501ef5722afe2c", x"f7ff90cc6a2ba03c", x"6a0bb344c8adb213", x"04c496a772ef2b41");
            when 26799611 => data <= (x"beaf28a335847c29", x"775d16e851f9bb26", x"0d9fa16afa5bf147", x"66742bd4be7caa47", x"cb657568d58f635b", x"fb0679cb33b7b39a", x"4fa9583952347afc", x"a7c89766d9cef1d9");
            when 12994284 => data <= (x"bbc8038d3076ebaf", x"dc036fc731ffc27e", x"82f11e6098bf02c5", x"1a42e98becd919ec", x"3ca9bfd26a269ad1", x"113b9e2459a5a5a6", x"54180dfb29ed2ecc", x"dbc2003185728353");
            when 19326927 => data <= (x"875a877636024dd4", x"dcb4e296b7903052", x"dc07d503db0a4cb9", x"e2444e028444c88a", x"82f709df93799622", x"81eadcfb23bfef89", x"e39a4e967e40cacc", x"25a23c0c70ff3e63");
            when 27998357 => data <= (x"27d0bb4359c3a684", x"904a8911ae4f2293", x"a6bf26be050179a0", x"57063706399aff66", x"94be4d6ca31352a1", x"651c1fa2e3432d70", x"379ba1623fe67623", x"0f6b2f83775fd354");
            when 10782279 => data <= (x"d841458d04d4d75f", x"3a170404886b6f23", x"94f994741a802309", x"d78fe9474e53d0e2", x"ce2fcffc041aba6f", x"81ad909b93343be4", x"49bd8a84f777cebc", x"857f66a25a3e8500");
            when 22537647 => data <= (x"a3d73bb37d35979d", x"1116e5f9d83ddb5e", x"0efb1645ba051eed", x"c903553e1c1b9721", x"0471addc6f3196b2", x"8b9aa19762a259d9", x"099cec7e75d43419", x"1fd112da5517cbf3");
            when 33449484 => data <= (x"e0d07e1819ad7266", x"91f617bf4b41c7b6", x"bd1460b620dc3d7e", x"8edd7747572781ec", x"2ea158f9ab643983", x"84fdfaec37baf12d", x"f2b1c6f6abc83884", x"dafad8055e12072d");
            when 1828070 => data <= (x"00f4e0a97269dedd", x"4579f822e82257db", x"35f173ee286b60ec", x"16652f48a156484f", x"2b0149267b98cc83", x"fc013f5202c38d55", x"1e4662d20f484725", x"bfd488552ce1e8b1");
            when 32436063 => data <= (x"65af712a209c8673", x"5c5dc708772bcf3b", x"817708ff46eeef40", x"22dfe9a8b0f87aee", x"12571199bd9dec03", x"be68bf9250b27aee", x"de7dbea696d0f524", x"09bdb9b898dde068");
            when 32712666 => data <= (x"2ac16cf8a69ac726", x"c37c4d3cafc3ab21", x"6918a208af247501", x"bc070c28b87e77be", x"c7a3a02ac02c6246", x"62e66656f59b06d6", x"92a74bc63257961e", x"bd26140edbafe976");
            when 19532094 => data <= (x"74384879112bd9de", x"7e4620c63ca86af9", x"db916a63b1429a46", x"5093282bfe7353f0", x"fe62910f3faac9a6", x"768e63fb5afbbd81", x"8b1c7f2c06208805", x"cf04574033918685");
            when 21494092 => data <= (x"190cec89d5a2f6a2", x"9ce9f282f26f5cd3", x"073fa92bf6e64b4c", x"db7edb4000f6eaea", x"8c774d2ac6c12bc2", x"f2e07440c6dfbe1d", x"f174e50f06a8f633", x"b197d69e886d4ddd");
            when 17789486 => data <= (x"3043c2cb380a2594", x"b128254e7da99550", x"56c9996261daeda5", x"0c6dee572fe03fc4", x"ed7cc428243551e7", x"78ee70734588b7a0", x"4a83aa088f507862", x"c663a3ef6b1f0de7");
            when 23509448 => data <= (x"a04157c944e43bec", x"8f72ac8dd0bff162", x"5b5ebacfe2f9468e", x"df11a42634bc1014", x"6e4ebbdacb29bb7b", x"3723d3d2dd5c7ea8", x"5dfb8ec88a8c084a", x"e61f644141472d57");
            when 7413007 => data <= (x"3b0926e7ed81c60d", x"82d84f49c4e97758", x"3ab63d2f99671379", x"bdc6115e7806538b", x"68abee7628ecf48d", x"bf033f8f50de21d3", x"ac9b1830068430b6", x"2895565cce942174");
            when 4565696 => data <= (x"f0a39a023f27018c", x"eea388b33d027015", x"8edae3489ed26461", x"f3063e417b9d3868", x"64f742b4af4f356e", x"96920fd35b1a2e9b", x"0665bc5ad5871112", x"16b2f43135426e8a");
            when 3738946 => data <= (x"9335a7f3df05ee1b", x"bbe537344a7811de", x"a5e94c5c96d15f7f", x"e39b4f591bdc43f5", x"f0c507a36417a7f7", x"7cb6c0914a52ca75", x"8923907c1711cbe6", x"07c29a7a31407229");
            when 25950875 => data <= (x"65ca59f3cc4aaada", x"f66d5af61a54bcae", x"656d00a56cf36c9d", x"1aa4c5e78a7500ab", x"b686b37b1762ebee", x"096212a53a22415c", x"d914b895db3fcc9a", x"ce90f56621ad55b7");
            when 22169555 => data <= (x"15df6c76db22f6a1", x"d6044c753fab4bb5", x"7c9009da4d36a334", x"db5999ac30633ae2", x"1dd31477fb65b4cc", x"86d4ba1b06091d89", x"3f0f4de03846e737", x"6151ac92304fddfb");
            when 28906888 => data <= (x"644c3e5f442961f2", x"106053114b990eab", x"78691f3bb78296f5", x"fb0f44b7298d4653", x"c29967580130e514", x"fd3659d14c991dc3", x"b88803dee51b8d7c", x"0c7c626687e022be");
            when 8380755 => data <= (x"e63b7f5e3987819d", x"0a62c59bb43ccaae", x"3429ce653e8044ac", x"76bf9a4974d6d21b", x"19a557337e277624", x"660a06219ca71fde", x"76afda0aedfc61aa", x"ef7cb10a3450cc7a");
            when 860995 => data <= (x"51389bf2a5abbca4", x"428af5be2d30144c", x"4ea170bbf893edc9", x"11c16025ff289f60", x"b7b1e8ba0922fec2", x"8664eed93cd03006", x"dccaf76a15299de4", x"0d618ffa83e0dfbe");
            when 12336861 => data <= (x"f27fcfdb81f82e3a", x"e876582eaaa34404", x"7a936f5a489a130b", x"fa3f914719a185c3", x"b8df5e539faea8f0", x"9055f5f7885dafe3", x"8adbf552e91b6bfa", x"9c7ea03c69bc936f");
            when 17768197 => data <= (x"a55eb9fefa8d4f7a", x"9080a90aef75d3b2", x"72f8d7d1fc8a3ca8", x"7a4db403286fabaa", x"c5a42112374d9093", x"8a3fbd3de72b583f", x"3d955207f47903d7", x"90ee22fb34fa1c58");
            when 12799331 => data <= (x"a2601c993fc7ca64", x"56300aaddf945491", x"a3ffb140c744af3a", x"74d9f81e3ce0055d", x"a95387e0ab7cf600", x"f44ee0610c66efbe", x"4248985f2c56cff3", x"05d1e1b3f5d48b39");
            when 4320638 => data <= (x"4a82acc1f40fb040", x"928d70398eb3b53a", x"55ddee8657828667", x"639c50c0ac119ef3", x"5f46ea98f84ae9da", x"e79611114e9ebb60", x"326ba978f4577a81", x"bf7541d1b5084a97");
            when 24982375 => data <= (x"ff8cde10788a7539", x"5d474fe577d001e2", x"ca98f61f8b7772af", x"386d989d284d086e", x"4543d6e5e95b9d58", x"3136d89846876986", x"16fd3521be5b69dc", x"ef060126212956f5");
            when 33803974 => data <= (x"4c688c640e72a0ff", x"41a9799738d9457c", x"05e025fda99fdde7", x"e22ddbe4b5c1868c", x"29d8f353514e59a1", x"8ba135a93dfc9f2c", x"8ba6780ed2f83f6c", x"c3a21e1edac2c71f");
            when 14135599 => data <= (x"2ca34ae01ebb3785", x"6c94e2b24c70bbc7", x"44c19da38bb8efe7", x"462edaf8e41bc3aa", x"19a325a1409b04ee", x"5c01ef92b5b42fad", x"8a7d85d24dce43f6", x"b541dd1fbb00fd02");
            when 28206933 => data <= (x"2b9a3f5e82d1a275", x"506d01679f8cfa6c", x"91263c7bbff4ddba", x"7d36d4522aaef664", x"b4e28bd0e5574a00", x"8f81ee05b36b131f", x"5b7da9b27c94ae69", x"a491d0cbed986382");
            when 21125905 => data <= (x"a5bfc8a804c42577", x"1479fe63c9fc5689", x"207e1a055b1340f7", x"e59eba844adba475", x"850493c682601dc0", x"30e677336f611ca5", x"ecb8c29bb60552cc", x"7cefc99099a7159b");
            when 28146091 => data <= (x"50dc7edc852c3965", x"d11de9b947e9d2c6", x"800c4f2ef08ba0a2", x"e2bab6d8fd22b59e", x"b1ef57929b84ef1d", x"b2db1049053988a2", x"0fa0e8c32af44d77", x"a55e9621c347ed60");
            when 3760243 => data <= (x"5843e8d0e03a9b70", x"bf6e3e88ebdb01df", x"19c621ff2c3be3d1", x"6f3554ab85aee758", x"4058d1688ffc7458", x"1ac9de93b70f0eca", x"a623a9ab79aecb1f", x"247edbc2b784445e");
            when 843862 => data <= (x"613f0a1a11870aa0", x"91197d639011183e", x"8beebc41ee133517", x"cd1cc0c03988ecbc", x"8374cfd6e3247bf7", x"40bcaa9cf673305f", x"4a3fddb0f820e9cc", x"cc57d876b6a02834");
            when 18770908 => data <= (x"f8c7a8f673b2c384", x"acd6b22c03f2cef2", x"95e4c689804adfbb", x"39e323009cd73d02", x"d0f53e8d2628a50f", x"85b1d90cae8023f7", x"1604e80186f12c0b", x"9f74b9f329cd2a75");
            when 16809913 => data <= (x"01b960a9089b0fde", x"d734ee281a38a458", x"702ef7b2e3580071", x"31e1951d0db9bbba", x"a921dde68ebd0004", x"e8feb6ba4a64a594", x"0f8a3b7997a78ab2", x"26fe8355249660e3");
            when 32223154 => data <= (x"530230301acdbcc2", x"6c64a11feb08dbb5", x"e199d7e177b0a225", x"04d38da110734a71", x"3c64ff4a053e01b1", x"36e3f2b8182e8093", x"13311e124445e82d", x"4b64b9a3b2474b4f");
            when 25807375 => data <= (x"0f49382d8198e37e", x"0feb13a47d254c6c", x"cf61e178d68d35e1", x"01d031e76ebacdf7", x"ac1f1186b5a0a3a0", x"e0b7256142b7f85c", x"bf1f1348493d6f4e", x"17f97522c1a029f7");
            when 19912292 => data <= (x"7a24c47c1da8f099", x"f26878546afbb350", x"5e09f53bb72d7f2b", x"d38118365961549d", x"9b74eedbf10774e4", x"23663a4208b98325", x"de2c089a39086580", x"9b15cae7efc6654b");
            when 19389050 => data <= (x"0c404519194063e3", x"cd1f9503d6af4d9c", x"ce2854558614f03c", x"d00af7bd5179b376", x"2d507aa0b2ca7982", x"2f63c697e9cc9bc5", x"c24e32ed93a18d4f", x"342d2f46ab992f24");
            when 5022286 => data <= (x"4bae77b4273c5084", x"fc6e0ab46974c349", x"4d1e41d5c1ccce25", x"ae0f5a5481063d66", x"b4521f181b68f992", x"5b7d722f4eac59f8", x"de33fba05423165d", x"7f33bd4d0401fd23");
            when 27821897 => data <= (x"d4803ef77dc9cae9", x"8b5ae15f4549589b", x"4c02ba7811d78606", x"0d663e2299a6fb3d", x"2e9a57afc8da78ca", x"437f2b8f35422f97", x"78d6e767d45d6570", x"a9c0154f0c5cd6a1");
            when 1669909 => data <= (x"5818abdcd7cf36c3", x"3afba5bc9301efe8", x"96ea89055cdab33e", x"b07e41bd3e60a217", x"c1b51d8bd105442c", x"c374520abe2eceb3", x"76dfa1c7261027fa", x"ad2e81504d867bf6");
            when 3128983 => data <= (x"ef675f7234cb2f70", x"d6092d8436ae3c45", x"b170fb61422a0043", x"259e59a991c1db61", x"50daac7185d17a2f", x"d0ede21dedbd4a4c", x"ec640b0fcabf7276", x"4dd91d726777555d");
            when 28603404 => data <= (x"6c7378beb8f2c40f", x"41daec03bfc0c645", x"106c8403f6e6769c", x"7bdc10bc839b613f", x"4c51c1351f86cd2a", x"3d73054e88286f18", x"16537b5e6eb55bf4", x"08c194e0bc3b6272");
            when 21513866 => data <= (x"12f4d146f49dd51f", x"0b492014ae6f37f7", x"af250362de538aac", x"863cb459ce39ad28", x"c80a632b2e32e326", x"1a64308a06795356", x"43d163dc2dd3a019", x"8deed1ec9643a242");
            when 10388516 => data <= (x"b1036e7c219d6549", x"42070947764ae68a", x"e13de88f9e84747a", x"2fc99b6f9e523f8a", x"e05b58d80a41dc69", x"b3300f4df4e26660", x"d73dd7cceab09165", x"c05981669cd61887");
            when 21106518 => data <= (x"623d4a9b5671ae13", x"0a2b11d020aeea20", x"9ec6d4364dc8b9a4", x"cbdaccece0b89f49", x"ebf2dcec5e1f89a9", x"3b235d89949f3f97", x"1e2f7d4d592a351e", x"21f7193b6c9d4894");
            when 21451586 => data <= (x"d5cf584c82a1c90a", x"5084950a82991e4a", x"8073aefd9fb97293", x"5a4538a5ae7249ef", x"ae2e37aca606c4d6", x"383d1f44196d635a", x"9bccfd931c43098a", x"513a7ce2f31c6801");
            when 33299809 => data <= (x"2ebbe91b795eefb3", x"b6e01f2ff617d358", x"fc15cdc4befa7be7", x"228c259b1de6f500", x"2e897c2ea9c4fda5", x"7a6228fb7ff40204", x"8b42ab258bdef478", x"80aa08c2d59f5420");
            when 14966460 => data <= (x"d58b7f27ea88e02b", x"e660a3bce6b748cd", x"16b5ce3e9a7409a1", x"9ff4aee0c05ecba8", x"afe8993ce7770692", x"f826b024aea3a231", x"48731e399d96fc49", x"160f1b388eed59e6");
            when 13793033 => data <= (x"dee510dd6859e74c", x"aac3164137ca4199", x"448e2cbec8b40daf", x"72700bdd6a6960f8", x"97375e824871d39f", x"2b2f54aa557fa575", x"8a8319dd66fffb95", x"b52fd33c404fd5ec");
            when 14198551 => data <= (x"6a3eb18182d0077d", x"92a8442e68b9c05c", x"7f1f4c92ff1ef68b", x"eee1ca6a6464005b", x"e5a94723cf5a0200", x"e3e469f2a376796f", x"f64a80a50d09eb37", x"e2b67712dfa74470");
            when 7392452 => data <= (x"db2d7d86a3527f70", x"6ce1f93a1d935a35", x"649503d3f1b67c63", x"2c9c37a6deddba5e", x"1401641f4d8d2130", x"128d5a0246f0cc0f", x"9b1a587c8cab1981", x"3657d8098445c771");
            when 17015005 => data <= (x"ba16bebfc218d82f", x"2a48403f3a292df7", x"aa0240a6b44aa9b2", x"f97025c0ded2996e", x"b47dfc257bd27c64", x"54574ea950ccf5c0", x"b1f8a68562f52471", x"34f1ca16017c1cc1");
            when 30107885 => data <= (x"a3a16ab971f1c744", x"e7c4500493e4879b", x"cfb94d9c6f34733e", x"07fb5c83bfea3dbf", x"d90ce67e55b8aa73", x"6c63e041513754e4", x"359b24bf33ed42c4", x"0369acdc61283edc");
            when 26975727 => data <= (x"020e299d4f48fdef", x"54d2a5b99bfba64a", x"fefd472dfebbf2c9", x"e97537854c04796f", x"bf3eff26c56fa675", x"4520d262847b1edd", x"9ca1e9241f65e53e", x"5c16416fe5a0be37");
            when 3373175 => data <= (x"5e427cbcc02a4a2e", x"e0cb07bb8a0185a6", x"658c013565d9478e", x"ecf7bac545e3bbc7", x"871bf3a0916846e6", x"e9ada722eb53ef57", x"994cf4662d44c187", x"fd58e822446bcc58");
            when 15625558 => data <= (x"27f84d3b8d998aaa", x"d7c89988dd173502", x"9193a89efa04cd8e", x"723d67549a0104fb", x"b004b9bcffe7d2b6", x"9d274372019061b0", x"27d66bbbd45df7f3", x"af787442c8315891");
            when 28640588 => data <= (x"52e5f7857acaf25e", x"64af2f1b900ccef3", x"003e0d44a9acf96b", x"7275607c3e23628d", x"c468303cbe0b1edb", x"60ecc35269cfad74", x"c5a4eee7133a4e58", x"6dff76d3e225c9d7");
            when 17347552 => data <= (x"9fd46513c17de46b", x"14062ccbe1c8d858", x"0ea7f1746e41dedc", x"b0a10138a0485cc2", x"3c75f9f0952640ad", x"ca1d39d7247a0d6f", x"036c8a16fd4d25b4", x"1aac01c18d8e9767");
            when 6858898 => data <= (x"7856e621be5ce9c0", x"53ff3ea7d9eddba6", x"50b7b766b3e27eae", x"0c29f53467aa0554", x"f7f36d5130338b34", x"62a42c1da35b02fd", x"cfead897bcbc770a", x"bab9b37ccbc66383");
            when 5998058 => data <= (x"4251ae8fb1484708", x"fca5d0e64dfe7621", x"2e29f445c536bd8d", x"aa13ab36d4f18267", x"a584beb8b24eb238", x"d25808c09448758c", x"5ccb1933107f8bf3", x"2807057ac3949270");
            when 23362099 => data <= (x"c069c217e18d041e", x"eead71200eaf65a0", x"513bf9b62b96f7d1", x"485e2985ec0198f4", x"5e8fa6644d06a9e7", x"d1f815652471b3ea", x"de2df4fdd20ae6e4", x"a93d0f1c3cb7e6ff");
            when 17010727 => data <= (x"65e77ca84be7a63d", x"8febb56d242df8a7", x"3591b8ecbb444faa", x"5235c232bf2daba1", x"b2b1ad52b125fd90", x"cfa38835862c634d", x"bce890d18b25c873", x"5f726a7ee2da237a");
            when 16473948 => data <= (x"4432fae79d05c929", x"f62e3b2909ffd2f5", x"ced9534c3da64e66", x"8d46de9c50d0b288", x"5a45606a8d970f99", x"747ac5dc504939be", x"af2e783ee821e7fa", x"90b862c618391379");
            when 13223668 => data <= (x"c39e60970637955d", x"b95e62d2376cb2cc", x"9bc3be74322a9217", x"886ab42d23c7e06b", x"621b4a7ecf7ece67", x"210b84f2255bb86e", x"cb2c548858a7e3ce", x"7be187f71efef6c9");
            when 14624763 => data <= (x"6ab1c8f401027e8c", x"9ed89524b5457163", x"0f18221d4dbf166d", x"a04e4e741dfd661e", x"2408b68a140b721d", x"0c84de6e282e581b", x"3079e5735db56ee6", x"83b8528e8a0d9df2");
            when 1671700 => data <= (x"547173d284e5709a", x"04b6e6155a8c104a", x"1854c42f957965cf", x"c1c6a2785ca98a82", x"fdfe37f4e1234c8f", x"faeb2bcda05cbc7e", x"ae4f223babd51328", x"e11b1f8a4921fbcf");
            when 9164789 => data <= (x"e54d4ff0649171e3", x"ff4c015b1c0685bb", x"c56a8e684b9c1357", x"ae3eaa3e6c0f4a70", x"5445dfabf309bb1c", x"b24dbb8cb51c8b9e", x"635c1f3ec8248c92", x"4b51c713299bb496");
            when 27192868 => data <= (x"6a2dae8fa3f61c51", x"8390c140762b7441", x"36a19766d8882bc9", x"135644b65ab19afd", x"4319e0d51d782c25", x"cc95e08df22961f2", x"8c27d15ca2c2ff26", x"1b38c9f2f8b85201");
            when 26453353 => data <= (x"d63ac9694066599f", x"46af2aef8d4cc03d", x"f45fd18b6e90e815", x"7077e12c4446cddf", x"9011d9fdc34c4be0", x"5043c7a0626c310c", x"83b6b8d0373a3769", x"b4e391c05ccdd7e5");
            when 959162 => data <= (x"12870376decc39c1", x"cb252146cbf8a2bf", x"c9b551f842694557", x"8d511c629c3588fb", x"14a94defaf3a7a7c", x"d4f74b81f5f76ec6", x"f82dbc64aba3d79c", x"9fa099ac3b790570");
            when 5499136 => data <= (x"a073001d5ff39050", x"4539f2976f020891", x"7c3232cd85e8660c", x"0cfec89e35366191", x"97d54ebfc2b06ba0", x"fc5ae518e5fcc847", x"13b25d920fc945ca", x"436226478362d0be");
            when 29818518 => data <= (x"80ebd9f2939e8ebc", x"837b2db14766cbdd", x"a0fabcb4b35a09c8", x"8f6bd70ab4a7cbdd", x"b97cacdf38d632f2", x"0e419f741b887b34", x"a927e25c27e6957c", x"691e9172b8605ce7");
            when 24547016 => data <= (x"260a57ce11e42e78", x"e51a22bbdc45023b", x"315a68d7cb40c556", x"7a71a32d55b01d26", x"3ab654b8ab58aba6", x"80b2a925df0a2411", x"0583738e65ff1195", x"f479bc8ee09fa8bd");
            when 17943855 => data <= (x"c560eefb221260f2", x"12aae835d0721605", x"8e2c324d3f55e1cd", x"67f144809151d1f4", x"2d5ed9fbffc97ad7", x"c7d9f2cb8e0824bf", x"0eeab387a01172ff", x"dcb6432e7fd3993f");
            when 16138690 => data <= (x"48ad53784a6a4835", x"aa3b50c8bab326a2", x"b3f9b6cfff342c06", x"d4b0cbd99a1eb6e6", x"6864f8f222f27e4a", x"cc13f05b23b09818", x"fff7fa643e5fcdd5", x"348662f1d187b796");
            when 32161295 => data <= (x"63333f32c1bd4989", x"563e8402798661c4", x"fd56991d1b289b00", x"ff4cbd548ae80243", x"ec89595d675ffb9f", x"4a89cada74c21e3e", x"47e5678c484ef099", x"de5783dd9ed90520");
            when 18817815 => data <= (x"b89ca049f78fe825", x"ff2d81f7c40354ad", x"02087f811552ac1a", x"461c321e774b7a7e", x"00a62f27b8b47709", x"371ae5ab35036e9b", x"81ba852878f68229", x"e97426bdfe6a0272");
            when 22299544 => data <= (x"6ed214e3723327ee", x"b9c73092f3e006c7", x"99cccbc88a777177", x"eaa06e8d1ec4a59a", x"9a3dd7b8c8390144", x"ecb2a52fbde87d91", x"1a4f3da7618368fb", x"cc09d9b39cca805a");
            when 32980416 => data <= (x"bb5b174c7f7e52b3", x"6fe9f04fe8deed14", x"56172b9f3b27a439", x"37f0e0a682774e23", x"870fa95f9484c9bd", x"7b461f33928d1f19", x"eda2639c397a8e45", x"bc0999eff2357659");
            when 29206928 => data <= (x"b645cbb11a230a74", x"9e93891135863b9e", x"8fbd7d35f53199f4", x"e29ded2dd7e25118", x"53f30fb4e35fdff5", x"c2689c6e55262ca4", x"ba075ec1ea4d77a6", x"47d3ee2ad26725b5");
            when 12188599 => data <= (x"a0426f0ed02bebc2", x"6fd64b1699482924", x"fd3c59f8f86612cd", x"e8c37c29eb88bde5", x"30c2421a79bc8e92", x"2e092e3ede902a2c", x"a28ec1fe3a1aca47", x"500e9cc5e3c4dc5e");
            when 8007281 => data <= (x"0ea511b4c106850f", x"c2f2332a519e961e", x"6ee356de41bc94c2", x"ebd818056f6186c5", x"318b6c0bc9a34083", x"6b780bba3f0052fc", x"6ef6c9bac6fc5044", x"e9b2f3491d08b636");
            when 28398261 => data <= (x"d870b4fdf3d0d0c5", x"0e8b2cd02e52353d", x"f1476d80d7f5d4d2", x"0c83d1a1f8cb4cf2", x"a5fe1acfb7d81bcb", x"4f32eff74448d687", x"19125c0cca4fd562", x"84675dbf0f2ec83f");
            when 7920313 => data <= (x"b748548eb8e690f6", x"e8690df76286472f", x"9aea83334c074f70", x"a7a806721cf37d04", x"480d82b20b3fc7d8", x"7c2c55903ea2887c", x"9f8002e5e62c04ce", x"81c5e269df4d1d25");
            when 10109237 => data <= (x"45b85905908d8c10", x"f7c945e297f6cf69", x"aedd2530b1e185f4", x"21bf1c93a19f2634", x"ceec2a6fa4c5fcbc", x"1f38c31c07242854", x"f9ace9a5855d922f", x"1cdf64de86a3385a");
            when 8814945 => data <= (x"cc2452c130a44643", x"f0e46c390ed96fff", x"1a757294bd512e27", x"5027f1e0467b4c1d", x"1e57292349e36749", x"072f02ae9dce6a2d", x"04265625006562df", x"db621aaa1201b06c");
            when 19223783 => data <= (x"b5fb734badceebdd", x"5d73b0010226172e", x"b42d2f9da0a4a672", x"2759ad347bac228d", x"1c652854110ad57e", x"3b72b95651376d49", x"042c9328e9920a15", x"1c787985c8fb1bf3");
            when 14852642 => data <= (x"8ba5ce0c914e058e", x"1ae3418cc7943b8d", x"5bd36a542007d244", x"167b55f85f2b4d26", x"078837f6f6d94a26", x"ea830dba25f62cdb", x"9fc5525a363a1000", x"2edd28e36f609909");
            when 4605111 => data <= (x"f8e6bb6010a7b2fc", x"b4629bbf4fb5bfb1", x"726d16e0344f8651", x"6778f24debfc4880", x"2bb663a75015fb7f", x"c555248aedfa04ed", x"e2881d802f336648", x"ad961d5454e82a77");
            when 32774959 => data <= (x"00d04663a10aeeef", x"6d8d315891e0c218", x"7b675eec0eeabd61", x"59b72abe353f710e", x"b755e5262756ce6f", x"d9a3b4bf0ae3a6b1", x"17b1a1f047a82773", x"e8d368297de45a1c");
            when 8705083 => data <= (x"a47075a8ea877774", x"809db4f2562e1777", x"9d8af14f899c0eff", x"69d9939686c7d56b", x"e1dc42cc7aada4bd", x"ea13ccc0a05f3a8d", x"2c0a4f800ac7d749", x"5e726e71afa9e69f");
            when 29751642 => data <= (x"7fa106ae0a51a6f3", x"2a1af0e6f65d8d64", x"6ea92283fe5aaf03", x"c2b8d2d0c1424168", x"42dc9e0b47f6639a", x"dbe781aca1819470", x"d4bc2c4176e9db26", x"938ef72d9e28e607");
            when 26441805 => data <= (x"12613d8566c3c90c", x"a8bcb60bffb7edc1", x"bba8af7413552dbd", x"06c7df1e66e65337", x"9cb6e1cbad6b2661", x"6eb087756b5c79c1", x"dc1639460ec1af65", x"8476db3aa4f02bbc");
            when 20196911 => data <= (x"c725f134ba23503f", x"5b1c3f3f46e0d3fa", x"5dc74e115694da8c", x"7a29ad4c2ef48c79", x"7f515f436a57486d", x"0d1a7d9edabffc2c", x"88121141c0facd5f", x"d8340de9febd0087");
            when 4660772 => data <= (x"4b6a434b1a8f4537", x"86ce5ad4b809bea4", x"829d6601411e6a50", x"2b5ba5215860c352", x"bdd1d091e6eafe7a", x"b6b70afe7385c204", x"ce5eaaaead2edb6e", x"702f273b9e0217f5");
            when 26108152 => data <= (x"f8db40c7bba38ae2", x"d40db7c1677e5d9c", x"0f7eb2d7989d9f88", x"b43e1cdbc2158e21", x"6c74c1d125e7893b", x"5e859ebd0bdbc4fc", x"b662831da39fd439", x"e89622d447991fe3");
            when 2342760 => data <= (x"7ab6c5534c332c86", x"3edea54442abad8a", x"20d63f4fe7b33c5d", x"298828c290cb3639", x"d4ca454b4175c76b", x"09aef3e836c612c5", x"159ab87e1652283a", x"78b392e32e3bea7a");
            when 4501156 => data <= (x"d9eaba9d5b9ce117", x"8635bedfe7c8fbeb", x"36e7afdcd560d015", x"40839e18a2bac3fa", x"17b505aa100550da", x"47a4df0b5bb8f236", x"1f2cc630c83eca5f", x"3f8d7c473e8d2b52");
            when 26259315 => data <= (x"98f8d683849f1224", x"667b6ec7a4125088", x"ba99b85668fcc614", x"e9f2923f01cd0ffd", x"85b0d63112e441c0", x"6f81cfb23ba146ef", x"d5f3e94f46c7b2b0", x"cf36d76e8413a7c6");
            when 29110268 => data <= (x"c7681f48280829da", x"315621fecbdca752", x"9cfa1672efb2f4f4", x"2c49ff79650c8550", x"9d4f39ab72c18109", x"d2497b5b16d5df98", x"18441376ef59c5c9", x"dd6dda1e97751fde");
            when 28621878 => data <= (x"72318e28d22a599b", x"5263c58cb13380a7", x"eebc76a7dbf1eb24", x"f20cfa6110c6265d", x"90c481d017d9c64a", x"e2287ec32716a1d8", x"c1b4378ce1d838e0", x"39bcce9beded9de5");
            when 33543991 => data <= (x"08308c8f05155a26", x"044363d770ff2bfc", x"9266dcf412ee2fd2", x"097915b6e71bc034", x"27d54d84121a420e", x"c03177ccbb6751e7", x"70115065338149e5", x"05a9e657cd78d747");
            when 28391224 => data <= (x"618c262a38eaa2ff", x"dde11e94b4dea079", x"6d3f8164f47d05b9", x"5cbb05b114164c85", x"958ba0711eb4e60c", x"b3e27268d90b3ec8", x"bec51629e2f535f2", x"4f3e07dc707036b9");
            when 14463831 => data <= (x"48c2d955c9123aa1", x"a7d0463e1603a49c", x"8e264a621ef614c6", x"ec61dcb5116f7127", x"dbe61ae3f815bf75", x"6b6a083b4f9d59a3", x"0205ec074f72b363", x"3e4acdf7dfb7cdd9");
            when 8087431 => data <= (x"a6e3096142bc20c2", x"6fe4c57d745e0cee", x"d52977b9e23063b3", x"fc01219b52cdbfb3", x"7a2f2e7f6259f8ca", x"e5d1447d6275cc0f", x"bb139a6eed0288ce", x"a3405fe7a4507eb6");
            when 13801540 => data <= (x"2d1ecc0cc70515a5", x"9bb68f1c5790652c", x"43e51f0c531784d8", x"a100e57d61228beb", x"0e76b906cb421b7a", x"0ad00e52a39bb948", x"69139b3380a243e1", x"50a839a852bfa781");
            when 26981518 => data <= (x"04b658f0e72d5a3d", x"ba18f746f2d38d1f", x"466af1f795d75b43", x"d39ad851b8a36f60", x"a746aff4f60c392e", x"c7b562214da5a88a", x"115674b290f2177f", x"b8613b2565d24924");
            when 9475660 => data <= (x"d0c316b80134ce1b", x"db91376b071c3cb5", x"ff0008203065097a", x"d6f7a3bd24630482", x"6bfdc2917aec1adc", x"93673a44fb59735a", x"549b0a1fa64c934f", x"0a4f89df66c5b115");
            when 9608471 => data <= (x"8f7744755baafdfc", x"8a89c95fe935c567", x"59e3523a273bb88e", x"1ea664ed93ab179e", x"effc13e9e72a0df4", x"4a2b3503e0bbdedb", x"17714ac11735f5c2", x"325e1ed8e230e97d");
            when 17883727 => data <= (x"307f9e6455c7e2c8", x"a14b38b642b729cd", x"6106b6605c3bc48c", x"cc617f5e260fc932", x"d6497c01f433633f", x"05dd83b25afc0cdc", x"6078b2a4532242d9", x"f31a6dce5e29c6b3");
            when 12698726 => data <= (x"bd5b1ab853cb78a7", x"814a2154fe660d95", x"b7f486015eaab17d", x"a3525aa2d0b7b2ff", x"94e1ccd130bdc3d4", x"c20f3ba2f16a276f", x"8d1b759750f12280", x"6d5145915e0e4b94");
            when 7283706 => data <= (x"a3a9a0bc1e6419b1", x"be64fd5a5c9872c6", x"2292fd48f3d83b3c", x"435d3ee7eb3c016b", x"16ec5c76f9b19665", x"30970d7e3786ce32", x"77cc47f0d6ba2e0f", x"ad93f2bc90decf56");
            when 22205742 => data <= (x"c7290c7f87b1a7af", x"e3b740a153f414ab", x"08a7294a754d44fa", x"4b6debed247847d5", x"448b2e3ac1e040ee", x"67f73849610a3d11", x"5421a35800335c85", x"defc68b222ddbc54");
            when 31730623 => data <= (x"636a43de946d8267", x"998afd233a22074f", x"8adaffc5f5147b38", x"3168a0a1f9fcf9f6", x"3369386aabfee0a2", x"def4634750ad6509", x"4fa0166630e52c0a", x"8b019da8ddd27d4c");
            when 33809569 => data <= (x"5f539068d77856e9", x"1c81076f5d9bf8bc", x"8ca2e950a8d3a991", x"7a3e36382241f932", x"ed52d107458027e4", x"8b335a14ee881450", x"e6f9c4da27911fb7", x"f95eb9a0c41d6ebf");
            when 18317786 => data <= (x"e49d217de7a475ff", x"614826062ef7c631", x"61b00f71231d01a7", x"051bc59dc9188e2b", x"3b709fb62d726184", x"91149e580395e27c", x"316ada52e918dace", x"26edcd6d301b98b0");
            when 31683546 => data <= (x"bd2f4f7a24c93f86", x"484a55a6270cef83", x"6d30ebe5dcb20c03", x"08563a1c7dd53dbb", x"fd8f39d84e56ed3f", x"21f1a98120de1c05", x"7a48e5f24efa7ee4", x"adab555b15b6d798");
            when 17050890 => data <= (x"2ee403daa0c867b4", x"2ef51d0cd4a2f675", x"d0bb5cedac80cce2", x"b9abff0a06b22f3a", x"f3810a26e16e3411", x"969ba6cd1109766f", x"4dc491ba8217851f", x"878703928aa21446");
            when 25962377 => data <= (x"e9fa4c6b955cb4ee", x"225372c5eb823de7", x"3c5fd90985eb69fe", x"5346d428cf5a2e08", x"2c3391c4c13a9b83", x"ab779ca5b91f7c7a", x"fa695f2fd4f9275a", x"8d31ed83a1210c8e");
            when 28784024 => data <= (x"4f1f3ccf1dcbe191", x"1c693a83b1c9f678", x"df3e5a3e400292de", x"ff6fabbcc5ee739c", x"26385ff8dda578ce", x"d6a23affbe85e090", x"c5eb1e6c3cb89c1a", x"aeb7ad01d44d3508");
            when 659982 => data <= (x"408aa656a2a25b5f", x"700c87be1fd329d1", x"71a9e0fc80d4c7b7", x"b106cb296f070e90", x"ef26f798282384c8", x"d44f0dfb9bf2f453", x"865c13a2d4e37782", x"f057621e83472770");
            when 22299682 => data <= (x"12d4827a27851aa3", x"289650eb1d3e6de2", x"c86d360b9a0c99ca", x"f1574fdbff41584e", x"7fa9784e91409453", x"2bb32e6a2b4c67f7", x"bd32a2f501e02138", x"07f970350c198c65");
            when 9359131 => data <= (x"cdc509f7afb1e51f", x"1bbf0c541a775f9a", x"d16cb65298fe67bc", x"b07d3a3f1532adb5", x"eaa544264177d2c8", x"2c72dbe6059fe572", x"0e4116f14ca27885", x"4bd36f226620ac29");
            when 20288574 => data <= (x"2d840f609eebf527", x"97e9b62e7530bb94", x"4317d186095f2bdd", x"6c23485812cdab3a", x"ea4285d128b65428", x"e3509514051fa1f9", x"e919ed5fdbcac367", x"681fe39d1f16d993");
            when 19274502 => data <= (x"90a1803dd28ff7e6", x"17b8c1f27a72a34b", x"889504d7c7256fa3", x"c0218a386294abdf", x"06003be6de959768", x"8d70eb99a29db980", x"237ce670ed141124", x"2f6fd24658902906");
            when 27956131 => data <= (x"6408d333ed63c192", x"a6441ea4ab104213", x"ad2c5c9ccc909946", x"22a5b84f6386ef3a", x"60fab24c008fbf5b", x"fabed04233d7c2f1", x"c7e47f5fea5f3d37", x"e4b2f46fe60045e1");
            when 19917690 => data <= (x"a99e64d74ca10610", x"cfef160244e6db23", x"717d96ca6c413e8b", x"c531d0d00223d3ff", x"f6732d66134f8c3b", x"f62ba64313348a72", x"30771596be6705cb", x"a1d5d39a927d9fbb");
            when 7649168 => data <= (x"1f39e29d3bd6300c", x"cf673085a35b60a6", x"948430e898a103d3", x"51a4693fd7b7f476", x"1f64cfc8968d8492", x"fe72e8a9331da8de", x"59d7b806d0b74d13", x"d5a282727bca8f29");
            when 24228907 => data <= (x"c456d4b7598c2d0e", x"d420b68d147f7c4b", x"e78f5cb746547575", x"00ff746c49f63acf", x"b2ecdf6e3fa952c5", x"737306752201bee5", x"4c4ccbda7409e0dd", x"9721395405d82e9d");
            when 29440936 => data <= (x"338069585d54ffa2", x"924da13f8519b44c", x"a4eae719b290136a", x"5c99f0d3d3cf73ed", x"2d418b6f88c89fb9", x"955a64dacf60a3b5", x"8201131f18ff7094", x"4bc689f62b291e87");
            when 28208364 => data <= (x"a0de3407917a5707", x"7da80466d8f2b91d", x"0dd40b21e1b9c117", x"6fbf9184bb2031a0", x"3bed2b007af9b66b", x"71b50da6a417a8f6", x"1263ec56a8b0309d", x"da912484b909b8ab");
            when 15642612 => data <= (x"c86b9c4fa5386fb4", x"ec30c1ef0484ee36", x"7a085d3b5e1550ea", x"fae41512c1327326", x"f6a99962d40d2a04", x"213672254e0fad23", x"89a45cc9c333e3bc", x"1049081462300abb");
            when 16651603 => data <= (x"c559eb988514410a", x"4ecbc20a2d089f43", x"47a3d4e6aaa43809", x"1ad1630f823e30eb", x"bb398cece96a6257", x"87d4f3423df95aa7", x"43eb3dbbdb4b97c2", x"f64aec69ab9fc0f1");
            when 24197556 => data <= (x"f4d957d6a9c4892d", x"3381189214c09438", x"260c9872bff74c7b", x"959c905ab5427ec8", x"1fd75c06d1dbeb17", x"c1f744d85f6bf02d", x"1a490a64a351aee3", x"4202c28fec8897e4");
            when 10812433 => data <= (x"99ede2b86851bc14", x"67b6f6a26b457c40", x"c5f8469ee22b81cb", x"0cfac5658a698ce3", x"10f0c0a7ce740a54", x"f46586b670fd71f6", x"03629d2b4a07e101", x"c98e09cb9bc8fc75");
            when 17768361 => data <= (x"c5ad8414fe72df9f", x"d148ebbd74e9cab7", x"4a4ad4f8cf3b2359", x"77e8736ef48a41d7", x"e4d08b98b9faa0f8", x"486fd2949f2ac5cc", x"fe86e3013c9d1f82", x"00eae9369382ae96");
            when 27514438 => data <= (x"39a1e9e5af8786a0", x"6aba873d28c3492e", x"86940800ccd17c37", x"bb173ed1342d9df7", x"8cd3f470d14a0cfa", x"08326d43799d7035", x"6ec7ef72d71cbbca", x"33e7a2a4e8cc8b1b");
            when 31872597 => data <= (x"a521a81a5f2f10c1", x"990f13537c282cf4", x"45fb4e62dea5aacd", x"5c41767bac8a7ee5", x"751d1d4705721695", x"46a6ae170ba9c910", x"a1bc9b3d104ec06e", x"b4fc40318ac18abf");
            when 20781722 => data <= (x"f26c9d2d7fef1836", x"ae83a32891fb0153", x"0942a2e797641504", x"8e44cc4a62ac8371", x"0aae3b9e0a0647a4", x"595fcd84227b1870", x"011d08b2ed10a10a", x"d9ca0bf143f8a576");
            when 20584917 => data <= (x"e4cbf95d205742b3", x"b908ab6030257519", x"1f4a6a1ec345400b", x"534147b67a8a554a", x"d0d37c7aa61404bc", x"4b4564eb0c8e0a51", x"730664e58132b3b4", x"a7f75d3b8c97efa5");
            when 31725117 => data <= (x"2dc26587c147661d", x"a5694c5ce245e49c", x"7acf5252d761bcde", x"2a285bf02ae53a23", x"737bf95b05b99c00", x"bca34b8a7c1c8305", x"ecfa68bfa7533c11", x"a87046c00207ed90");
            when 30595517 => data <= (x"ba06ad53a9614b6c", x"6954d41c4f2e331c", x"a3db9cf1f13bd961", x"5fd2f773084e2424", x"c1188eaf517f7410", x"d87bdfc2bf5fbf7d", x"ae93870351272fff", x"963005d0893456ba");
            when 22232938 => data <= (x"5998238610230034", x"d3a28482e37a4423", x"7baf0fe94e386059", x"5297bc6ac51e8ca1", x"07f18fdf0ecfbc63", x"e089295b8b862db3", x"75f3705048d693ad", x"936e2d78083e068e");
            when 27463834 => data <= (x"d5e68cc7a91e6a74", x"eda91fc22a7dc7e1", x"51e3e9450cf81a61", x"6a8b942ce9794707", x"1958eb69eb1702a8", x"e34fe1a0159ba2cf", x"9fd0efd3e2086cf1", x"9e78c78943812ea9");
            when 31976780 => data <= (x"711904dfb5aba2b7", x"56f12a516384005c", x"1ddcc1edc9dbadb9", x"f92148db038c541b", x"99cca46c7742f9f1", x"4aeb10cf15d9f75a", x"f89e8daf8c14dadd", x"0bf717d042dca6f5");
            when 6070557 => data <= (x"48b5e500ceb479e3", x"6477e051338be659", x"bd0c8c8a931137ea", x"16ca7f5141adeee2", x"3fe855eb3bfa86d6", x"01834a49d9ffde5c", x"e6d5c661f248936d", x"3429bf57a70b43fd");
            when 13875695 => data <= (x"ae621509d4ac583f", x"b29d37176fae908e", x"07f906e6c10682bf", x"b648239ce98db4ff", x"8d94117c807b554e", x"897b5a36ddc935c1", x"0ff132193191aa69", x"e764d5279c10de75");
            when 32361887 => data <= (x"07ad6c4125d5a026", x"bbc8c0293a15ff4b", x"9bb3d302edb3d1ae", x"fe42a6764b25c24c", x"7e04e14025695043", x"0fc6ef3a27d080df", x"f35e98217085a5fd", x"43547965c9f69b13");
            when 24589400 => data <= (x"521d56dffb5b36b6", x"53a15979f79dbce9", x"c27192acdfa1b43e", x"7a3290cd20706f72", x"a4836992137ed81e", x"f1e6e1cfd144f462", x"f001c4335ab0fd4f", x"8289e1e236beb4e8");
            when 23344006 => data <= (x"fc25a24a7b3fabf5", x"5ceba025d6d4740f", x"ed04adaedcf20f02", x"85773010d98c2fab", x"4a091f9a388f790c", x"b240ca36d091d1b2", x"1945c80fe30ab10f", x"ded019a711300823");
            when 9739809 => data <= (x"d9dac0aabaa56986", x"2d64d992114cf919", x"8d8791682226e419", x"1a7aaebce9de8cff", x"e49d9b2780143786", x"e17e59ef643b8b32", x"f65d2ccb3a1de53c", x"646cb814a7e966a3");
            when 9894051 => data <= (x"52de2d561cb23358", x"2bade83ec73ee951", x"794f9ba14bada760", x"71347fa1d6915bf7", x"806978cf9183dfd4", x"b2ab6101a480afdb", x"cddb69d7dda09ff2", x"42bd4acaec63eed8");
            when 5503840 => data <= (x"4049f69bf6583fb4", x"a163d5fec461b865", x"52069d6ecbcde8fd", x"eb7801dfdf881d68", x"d9335cef41461c94", x"3c1d472a041723db", x"b27aca91ee9e31b7", x"c1ae26105d400d77");
            when 25928172 => data <= (x"655c432d6007da42", x"b764f2e940e0310f", x"21a9f42122bd08a5", x"66ac4c07a63f3925", x"23663ab6d41af659", x"68ac320aec2d0d12", x"b2f586e7392eeb3d", x"090a517e486dcda7");
            when 27226298 => data <= (x"3152f75a511c0f71", x"3a9fc74d3d4b8b6e", x"3e5267cb9787ec27", x"fd69af3d352d0a36", x"bff9cf8c65e4339c", x"add46b2e3e018e2b", x"9b218a9e69799892", x"e7b51c18c30b35a4");
            when 16147548 => data <= (x"f25f1af0cd87fc73", x"593c6133c3fda1c0", x"37b11170be7c2436", x"fc8f2f25974ad7af", x"9832ecacdde7f40a", x"626be5ea847e899f", x"e797a39f4536b3ec", x"fc19aa93e66fd729");
            when 25110956 => data <= (x"0f00da31dfe5b952", x"a7bbeec9255c9ab6", x"f7386a326c277f50", x"0fd5cefe1bdafc29", x"21fe11303b8b2590", x"9b78b2171311aa11", x"908a4722ad0ca2bb", x"2cb4d1481c9430f6");
            when 25634821 => data <= (x"1c66780ac1185a12", x"78533ccdc9d59db1", x"465298f88700430b", x"64072e31dd10b8f7", x"d0ea58b878be33de", x"ced9792c18642f74", x"ef2061d3b229f275", x"9fee4b045e5e88c2");
            when 16843119 => data <= (x"bdbb7d35c1a0e2a8", x"d9f7cb250a64a7f3", x"6c5edd458bfc5bc3", x"690bd0fa99f13e3c", x"9f343d0906c94ade", x"77f98e6194cbbf3a", x"431d67b1b92490a9", x"71864be5fb4a56b1");
            when 3552300 => data <= (x"8727df8d198b8d7d", x"967247a29e8e1435", x"faa90c17e5ffe1d7", x"e8fc7c764e9d3fa6", x"a5a283afdd3595da", x"f4bf47d4050aab7b", x"991172ccd2bc3499", x"4dd08f05b7a3506c");
            when 28264202 => data <= (x"5f674d7646d2f94b", x"d695769f242ce2fe", x"73b3cc2ec9e92f31", x"5d2bc684078ff6bb", x"af8692f46df63b06", x"c91a3a2791ce757f", x"162e46727dae815d", x"93a18598da17b35e");
            when 13978921 => data <= (x"f04488c45a62ccf8", x"b21669516e4bd424", x"445b6221413d7c82", x"7aeb7f026f8fde20", x"197a25035881fd62", x"28deb122037b1a81", x"ae740a0bf2121c46", x"6502432583f39ccb");
            when 32923345 => data <= (x"323e390c3f556057", x"aee33eb414f44970", x"ec703274797738a5", x"e4695981ba14d04f", x"60727c85103bebb0", x"57b259e932d47006", x"ca802432aec4d9b9", x"ada08ae3c81e9471");
            when 746239 => data <= (x"0354d092850f208e", x"f52bc6c88eaa7365", x"10ea3b7da976de91", x"8e8f5077e2015541", x"0f850b3a2727b8dc", x"e73ba93f22155ded", x"091e7331c8e98708", x"9b8f2a59e401817a");
            when 2946172 => data <= (x"d019ce5e92562f22", x"4d6ac90ea203b2af", x"939d3593aac6467c", x"6e9fb915b1b42352", x"081c4d2f24e222ae", x"dbf5f9d2045a27de", x"1437f3089bb08bd2", x"bbd34829b7dcf888");
            when 30938558 => data <= (x"a9e4516a543d1476", x"2cad13b677456fd8", x"0d2264a9dafc65ae", x"1e54d2c0f3a477cf", x"c0c83404f40b90d7", x"ef318658eecbf5b9", x"3b36e73b0e29571c", x"330ffbb58494cb97");
            when 2439238 => data <= (x"640f063557d4fad3", x"1d458d0d4b2f6067", x"ff49f59a9852fcc9", x"a11c0afaba6b024f", x"ca8148eca58d1e66", x"15b81c6d1a08be2d", x"08acf2a13e4f08ca", x"1d3d6939f1135bfd");
            when 20713578 => data <= (x"10b68af7dc20ae32", x"32bc8b9ee7ab6e9d", x"db1c2b7179ed9db4", x"7ed05d95d3fe4903", x"7f8b04585ada09b0", x"77a81518b3c4d2d3", x"73d686715a0143c5", x"e118d7d38ffd578d");
            when 24142136 => data <= (x"10b8cc8f5f8a5901", x"3d6541193cde97a7", x"1e3fc4267a6d3e56", x"b330ebe0ffb20590", x"3cc6739f30fca64d", x"7acf4d1e5b34883d", x"b4989095b0e52e68", x"a08edd7d803ca7a0");
            when 26236597 => data <= (x"2543a2d3a3a51dce", x"27b917dc85b98e7c", x"99084ebfb085e785", x"c3921bc174e17646", x"85f92fc7acb30c89", x"ec3240638c252709", x"5dc5981e343a54c9", x"d20ee966a7adfe14");
            when 6431463 => data <= (x"df0b5e711394498c", x"4f1cdcfb78e9a02a", x"f201b326589e7f2c", x"0f54494bcc8b9b52", x"006fcb193f315b80", x"e6ccd987713c05c7", x"5e0789b8df214f11", x"ad39a2b5ec34af6c");
            when 16850619 => data <= (x"155d6dbe7b4e99ff", x"d1f2c79b23721f32", x"3ab4604caa0f9463", x"7df5e491e27d566f", x"3be42adeddcde12e", x"d59398361f808890", x"ed4a2d5e8cd94e37", x"45339358e37d46ce");
            when 29078327 => data <= (x"b3000400b46bb63c", x"a533a5df3752e751", x"6a1d730b4fc5ea47", x"08c65f6ee91183c8", x"272b58fe9caec7dc", x"293d1419905ed184", x"7e46a327db9b9002", x"55a0814de2b045bb");
            when 17099260 => data <= (x"8f898f854c4dfea0", x"cc18c5512ee44c7a", x"b3e29584011b8ffb", x"98743ad992da69db", x"c6a18aea940c5984", x"4daa9b3cd19ea09a", x"458007dd8749c699", x"f730c9e9f954af74");
            when 26473552 => data <= (x"364c87b02a400075", x"0bc512b42f58ede0", x"454f51b447bec648", x"ed205ca7f4d2915f", x"d7fafac39c54e3e6", x"57e02756eb148e33", x"cedd2e3d6af8c47e", x"0c9f2231bc2eeb27");
            when 2378431 => data <= (x"fda0ddab5e1c2bff", x"aae862bf9a9bad3d", x"17bfea8a2d34779d", x"072678433a5207c4", x"c31f200587024b76", x"8bb9707e99d524e4", x"c722231c4becd224", x"98509eedea15f4d1");
            when 12558753 => data <= (x"e825b086db5a7bf7", x"4c30ed0abc41d0a2", x"fbff34675b2b9168", x"298c52a89471c537", x"acf67d849e3281cc", x"c257c38811ece202", x"457f6fea0ab497d1", x"3cacca8233747e4e");
            when 27364939 => data <= (x"5a6ccc32d90e4156", x"5af337affa6c701f", x"f31998cece6f99cf", x"0c3fa3b9bac3bf46", x"fd906dc9d6673f89", x"b4c36a9a0b27dc26", x"50e759877ac8cc06", x"8c63f42969e628c1");
            when 31134730 => data <= (x"d407e044447be1e8", x"7ed70e461de004f9", x"b7c5409c33368a60", x"9783acf4a5b720b8", x"4c50f2847ff1ad10", x"982afcffd1795d61", x"2c0ff55a7f587831", x"c3c2ad148e48bd4c");
            when 21909594 => data <= (x"befac50e30054e45", x"fa206742d706e22f", x"3ae8772af930e8cd", x"f12b5828f5f7487a", x"8f7ba3ad2d0a6647", x"4f8e34f0407a87c4", x"ddd9a6be4b0c02d3", x"904e6d593e360239");
            when 5053998 => data <= (x"2742683a57058bd9", x"af25d7028c9b73f4", x"bd67dcb2a359b55d", x"d5d436bf4c748340", x"56a741a21db5b3f9", x"6cde6512d6338461", x"2980cefe96b3e890", x"1b2cf549d8fa88fb");
            when 936801 => data <= (x"e8edeedc93923cc6", x"b99a8dc9d8613934", x"754ab6a8be3f03dc", x"830631ab95b369ce", x"bab103432971fd4f", x"6e4291399a867a15", x"ff89b4475f2aae29", x"482fb7359b385932");
            when 29569363 => data <= (x"296363c479745cc4", x"197a3790910802de", x"30b3f67fb5d03d1c", x"a45e0976e825fe92", x"36de5e62d619bc39", x"09a61317f2940c46", x"ab30d3d0ab065787", x"f4030b939ca2435b");
            when 12048599 => data <= (x"647b365d90314b64", x"8515d8a0f5ef57e7", x"5ed92172c8f2a84d", x"06927290e4912c89", x"20057e5a0d50c0e0", x"566ae253e3a49288", x"c30db6cf11dc6a5a", x"5f23a4bce749749e");
            when 16989246 => data <= (x"6f602a7465a93c11", x"7866ce6279eac83d", x"34f8ba218ba80783", x"5aae0d86b3cf7e21", x"5505f8430541d78f", x"eed4b644b0ffe7ff", x"6b5c48522d52d80d", x"d35006c0be579cdb");
            when 23465654 => data <= (x"5dc80a5c1a80dde0", x"cc94190c4be10401", x"8f592a29e752377e", x"6160402a370c1e8b", x"20ae23ab64bb3a17", x"7b3bbd268d4126a5", x"7ef33cb317227869", x"61816047a17a6552");
            when 3136434 => data <= (x"5cdff2e0f5d34787", x"361f8d007bfab3d1", x"e8a1f83345bc543d", x"c8e89983c36c07d3", x"16a3e285b8385a5d", x"aa14150179d027aa", x"40c5b1f9d0d64959", x"0ff4184a15b51887");
            when 14574888 => data <= (x"d4c2a6d778ecc37f", x"a0ab2d058ff64b7f", x"a2f1ba24080172b3", x"3119ce55b36a6fe3", x"d716229d010fb1d7", x"3d00f5525778a36b", x"4b53576ddcc552a7", x"44653f75f0bd05b3");
            when 33119935 => data <= (x"39fd84a70467e3c4", x"0e3a09c3c0a19d85", x"febc8d4a6e524c63", x"7004fe696d03362e", x"7e1f0cafb5107e0d", x"d8cffafbdef9bc40", x"cc9c585295b4b040", x"8f6cf40699fbec1b");
            when 30682177 => data <= (x"e20fa47d86f96731", x"572667fb47e5ccca", x"db1d1af6bcc82269", x"059845f07894b927", x"ec6d9b3d777c00e4", x"62c08757f29e3e3e", x"36cb8b70a0f39c9a", x"614fd184fa6cb9f7");
            when 19283838 => data <= (x"3f990d888494ea76", x"8c3777509f65b9db", x"66944c3d5f87a485", x"96d4a8dc99a53d9e", x"3c71a8fdbada0eb0", x"1941e2bf3c45a608", x"f9158eef39a7125a", x"1dfbcb531aa70b0e");
            when 20295958 => data <= (x"2ab649798c9a0bc0", x"029551da10af0e2a", x"29007b35a0085c6e", x"b55e5ec576f4819a", x"2d622785791d4a8b", x"0bb56ccb4fc2e772", x"37223e50ed5fdcc8", x"a561ec9d38991950");
            when 23898546 => data <= (x"fa3c2df3afb19e83", x"d68f0dcee644d636", x"bed7c7bed4147950", x"d1d3daff8a8da3bb", x"52abb77f6adc711f", x"662cc0971a01beac", x"f58d60602ff6a238", x"114e115c187780d9");
            when 26341465 => data <= (x"841adfe0f61e6dc7", x"662de6708d0022b1", x"9ce61189ec86cc81", x"68719b4d94802075", x"000cae0849b24596", x"a62db7c13db52140", x"48f624ed5f4941de", x"49d5f460ab47bf50");
            when 24540855 => data <= (x"bdc173acb385c44f", x"ee12b97c1b4bae0b", x"144f96f498e27f16", x"1adb9c935acea85f", x"aa3470148372d356", x"0a0a56294dfdcd89", x"c4ca74ccb2d5ac9e", x"d9915e6a66e27bc2");
            when 10264773 => data <= (x"5fae27ff45e2cc1f", x"dd0ca9af53fb6d88", x"fbbcafe3cbe89cde", x"e563e1fc01771a48", x"80b6c3ce6cc7dd02", x"d5a7a2c77dfc94ef", x"0fee7fbf8c846ac7", x"97a94249c5ba17c7");
            when 20655189 => data <= (x"3ce3ab30ecb5ba59", x"e2462e31c3c52e62", x"a5af6f649290f575", x"31028000f21b2714", x"72ca24a6a120ffb8", x"c072d3706b2754c9", x"6336cd25832cac2e", x"398c416ceb2da70c");
            when 10387405 => data <= (x"1eaa072cc46958fd", x"58c9e9eaafa9f866", x"4f96f810f5b8bd73", x"7f0221d8741a1f75", x"46b9f267435315bc", x"470aae3543e0e822", x"a676ea7db41e1f2b", x"3ffaa1f4651263e6");
            when 8177232 => data <= (x"421b2ea4142c8d1e", x"04c6e32818301434", x"a29783a316029111", x"b43e34f190a08338", x"ca97a23c3ccaf43a", x"b6ee450f2dd787b1", x"7988ccdd24ec572b", x"e2c739c3863d0f79");
            when 25393309 => data <= (x"50490ca56a3fe3a2", x"7f00522696a1ce92", x"b27e4357123f190b", x"59139f1256658d42", x"75ab880817d06257", x"d1f18e1a39e2d0e2", x"29642ed31f679e15", x"e89ed43efbf8546a");
            when 3019178 => data <= (x"32370ede788fa7c8", x"b19ceae8a292aed9", x"a94d0d1640cc43b8", x"e971e554af620b13", x"df64f0ed06922884", x"b307b3abe1dccffc", x"5ad73e3317c9aabd", x"8366d3947dacc803");
            when 30347550 => data <= (x"f741e6b7b700e237", x"58cff888484832f7", x"ce05ec4f2d065d22", x"1bd4cc631a51eca9", x"f13796c05cbe523b", x"ddfe667950045e16", x"6b2f32cc1fb52d4c", x"bd9f0d8f0288f2ee");
            when 9672925 => data <= (x"e42154abf3519cc7", x"a3751d58df80c09e", x"ee2077b0aab1b199", x"fbe24322af582a0d", x"2a08c12a0a261589", x"ed6b83df8f8d9364", x"f8d25e2a8c1332ce", x"530db5d9238f5a2d");
            when 17799505 => data <= (x"1259ee59d5ecb068", x"5353753fd0c94ef3", x"fccbecc55fb65cbf", x"8766d17bdde35abd", x"68790c13b1c86f61", x"71e82219608d3fd7", x"f2f82e65a092e1cb", x"8489a1d6bb44dd59");
            when 22826667 => data <= (x"17e4578cfbf454f2", x"cfc1c038138de2d7", x"f719b94f384e319b", x"2df1b357cbab991a", x"04bedfa8d3df5366", x"247928c4051b6b5a", x"d616d2ea3c6b8903", x"99850355dd5b5208");
            when 10843315 => data <= (x"b36993d7bbe62c74", x"462e596b1153d063", x"a678f74c24b4be36", x"c81ee817b5275b1f", x"40424153e809035b", x"b73ba965036fad1e", x"7cadd61345669161", x"a77de1fb9eb668ca");
            when 3128616 => data <= (x"bb8086f1414c01cd", x"735eb9b7987bc538", x"27685577ff4d37e1", x"796d33f983494860", x"b45d37e747780593", x"eaf0689cdf4cc84e", x"8f78a9da8365a948", x"d75d5bad84bc18d6");
            when 3301665 => data <= (x"cfdfd823a0e414dd", x"6b7977ff9ef166e3", x"5e693f7a03ac9619", x"eb27edd3e0b83bd2", x"80dbe6a85a006755", x"0627ecb61d2eaea3", x"0272c2b04f28354d", x"c43b08201a8a64ce");
            when 12791864 => data <= (x"7aeac08d298c63f1", x"4c66e7b351795538", x"437bbc5fa0310564", x"2ddfcd27f2078cbe", x"e8dd60e2d587bb46", x"f9f8135acb46658c", x"ff4b3f220f9cafa2", x"be688a2c94371afd");
            when 25643761 => data <= (x"e767d3083f81443e", x"12eabbb5ac86ad1b", x"7dcc25bdaf63635d", x"3f2ac6f42dfc734f", x"8aad3e0f4d7a0c71", x"419e1135cb2a65a9", x"857d36867786c571", x"7de42c30481e3585");
            when 27484656 => data <= (x"21e9c5a581a03817", x"fa48fe2ef2c29edc", x"ea57ceda26c3f114", x"2a4f86dec609c2b8", x"3de4d2f9a229dd93", x"4cbd1420ff293f1e", x"6a62d04f1f306d26", x"4ea72d06f8f98a9b");
            when 28778780 => data <= (x"4cf7ad75e74fc30c", x"c5aa1829c0396170", x"07eb163d7b8a1309", x"6e62d4c7b9b488c8", x"e3758f6792fabfd6", x"a0e4ff0b722b3d5e", x"08b1a97591e37cc0", x"01b8e0ce4c1e51e7");
            when 10060533 => data <= (x"5b85791bdf6fe1dc", x"ca1afd3669bd18c0", x"bb94fbed6f79a7a3", x"d722999016b8d3eb", x"4544ed0b0807ac18", x"1a729bab2d5ea9fe", x"8b3e15e45618fe83", x"7543c35515987fa0");
            when 12380203 => data <= (x"01ae7d1c34fcc297", x"268b0e49c8eeba24", x"704235792295e8c3", x"cece655f9f2b5960", x"93a7969e541ad9dc", x"1aa8d5a7f9f97e3d", x"55b9968d8486b426", x"b6aff3119aa3bd60");
            when 6970743 => data <= (x"df9e2c215ea598d5", x"6de36879b37e5d07", x"a34500a699a85166", x"809ca0e277bde0b2", x"9fe7d398191e2144", x"50895f9fc3e8e4d6", x"86c4ced0a755e57f", x"4401740d7a7c890e");
            when 27549158 => data <= (x"39101ca1b2421129", x"db4cbf8bdbd76773", x"b71200e6371d4f81", x"308910090d92d037", x"1552584a3f07437f", x"9ba34fb19bb57272", x"c0317fa4c1dc2ce9", x"5a5525ce0a52e060");
            when 16593016 => data <= (x"fe36b13c33992572", x"be99d5fabdb86ea5", x"1cdf6e099903e55d", x"373949aae6cd8f08", x"ce557e886ea841d2", x"abcab8cef11a5f92", x"5be5938ba6dcba07", x"b58b31a91da2bcf5");
            when 26603862 => data <= (x"4f9593725e777571", x"c45021e174f1d485", x"ad043e2cf27539df", x"2b339fdcb88be401", x"e09d73e9aa8bed7a", x"2b96fae30240aac2", x"357d4c8b5df38e63", x"229d43f4b798a66f");
            when 10511473 => data <= (x"37cfac66c5573d49", x"e8d31997c400dd2e", x"0734f9275d42aeca", x"4bf13de03bd2b42b", x"07945dc84db34e62", x"ebe623c7998efc08", x"25060dc5b257931d", x"0e80067c0b635459");
            when 387890 => data <= (x"b1fad63b91eeefd3", x"1e707edc12d95f50", x"a4856675c44897b0", x"61a4b5d3f8bbafd6", x"1bda3acffee4719d", x"25f88b840573e05a", x"058d492f4c5d8d7b", x"fe896220c59ff933");
            when 26773677 => data <= (x"3e88ed9711e7c756", x"64efa66e6eccfa63", x"21c47c276acee2df", x"c2ae3963e3e0ac9a", x"69341f31de498a03", x"4c6475cb20518d10", x"6d375b790524ee1a", x"d8acb46d04a0f840");
            when 33056277 => data <= (x"97f07c96ba945a1e", x"13217bacd9cf2420", x"3350b24caf9ea5fd", x"77d1bff38b846af3", x"36452b669ed00c2d", x"654b63991b9c444e", x"f0a1ff2280d79ff4", x"4d13d3bcabd2c65c");
            when 26417692 => data <= (x"b0c3ce084e9f1a39", x"8091bfbc54a034d8", x"d91cf36da480a11a", x"ffa4f7c6adf698b7", x"81e86cb3515d754e", x"3019ac73e8b3e423", x"1e301b76669da88b", x"1f1d50dab72fa08e");
            when 861924 => data <= (x"4e745e8fcf83d9dd", x"aa87c4905b9a0cff", x"1f1eadec1914f014", x"acfdcf6ba88eaf1d", x"c25bba429e8714ad", x"b76abcdd4b92978d", x"afa80eebfc1835b6", x"78b40ac91af159d0");
            when 1801626 => data <= (x"23a25bb96095767c", x"800481272d7cda35", x"86f43471f7f466fb", x"cbec044aa54886e7", x"804db4e1e9fa032b", x"919d9d6a4ee187a8", x"2cc821e19d7a2560", x"6c8a46acf883aaad");
            when 32653448 => data <= (x"213f3f6622015af6", x"ca27c0ee34a26cbc", x"c37aa1f3e25cb5d4", x"5da61a0cae746322", x"6ed6d7a69482df00", x"dc6afc75c76de043", x"8b528fa1ace72299", x"7d11e170f2dfe6c0");
            when 22461614 => data <= (x"3d5a89c8ccae7533", x"9900a3cf3f0fd494", x"c823a08fa3a59993", x"2178ad8555f52345", x"8f1a079dbd3ec159", x"b79cbfc856cc32d8", x"8e8ba76de893cc19", x"5aff32558598c0bc");
            when 17231476 => data <= (x"67d95f1ec9d51d54", x"267e70e4b7c28e0f", x"265eab1c00b28d44", x"b295eaa9ed7f2ec4", x"504248ff4cdda5ea", x"5f93fb0572000153", x"ba2d6fb4df9ba6bb", x"bde7163b4e4c7c86");
            when 29110133 => data <= (x"c339e1b9ea362e46", x"f38ab2da03543874", x"f90837fb3037f89e", x"ef7e3bd63eff0afa", x"823d588fdcd8b7c3", x"be6d78f43111acae", x"2085a517af454480", x"2eb68ebe51ae04d6");
            when 17324759 => data <= (x"a93a8b39a7e77f89", x"2cd47227fe408673", x"3d7844a72214dde9", x"c41abef1f3801473", x"a517544b7a8af6ed", x"b4e1c91fbd8e3812", x"431191918d2abe8d", x"870d8b3ea2e1e866");
            when 31431768 => data <= (x"1b4c4692ceeb15b8", x"f3fd2aa4ef4342d3", x"fbe72fb4df84d47c", x"f487cc864f970d34", x"d8c2dbf3328f0e68", x"02438a23e6253b69", x"4355a02a64667be9", x"1fd328ba6a7ec54f");
            when 20810542 => data <= (x"1b5ce827719fd2af", x"295ad88025714691", x"1036e0577d610796", x"6b1cccc3d9fd31e8", x"020a1b544d9dfb6e", x"54b0f1387792d11e", x"3c8c274528b184f0", x"51885f58e719a165");
            when 26894979 => data <= (x"2257c4f271462802", x"08fd6623bd7fcbe2", x"415f9af9f3018547", x"6e0581258a0b0c1b", x"48236aada61d1e30", x"cad7e44fa72300bf", x"01260209bd1d0aef", x"f244f01dcd35d092");
            when 10379129 => data <= (x"609dec2df0911c6d", x"930bdda109443c0d", x"76d9ac4b4eabbc97", x"e5664f49541f8c87", x"c779738339a4c5aa", x"76e766af40604a39", x"54f63f64fc30dd0e", x"ebf15258e59c73e9");
            when 15927050 => data <= (x"856e44895191d8f0", x"bbfa5ba6e70fa833", x"c6f39ed6099c3565", x"81bd58356e3c4cdf", x"028a438c665878aa", x"6e4c3df9509a9336", x"82a5b5658a6875bf", x"df0d6b4c6fd73355");
            when 6233169 => data <= (x"d6f0bfd4db94b4f7", x"a365f3654a4380d3", x"ed7b2896f97e756c", x"6bad632af8bbdb55", x"18d075a1e1115fa9", x"f2991c3461bf9154", x"7fb6fcc5a06de919", x"8180560b1790814c");
            when 29198783 => data <= (x"5936b9859f7826d4", x"417dffe7fb621de8", x"42418c696e634880", x"25c959ee6b0d6ae7", x"81fb764c986c3dc0", x"b5c08e7fdd7b0d18", x"ea3c132a2ff5ec3d", x"a801a39fa6390312");
            when 10899282 => data <= (x"d6b3d05f2a95f271", x"bb8afaaed9019bd5", x"dae3c111906e0e34", x"7ded53b9a109ce88", x"9b35d1896a563d00", x"893d8f749ad16daa", x"2570c73522cabee3", x"915e5a21937ae92b");
            when 26674764 => data <= (x"f82d20faa1598319", x"0b5cf08ac9cba87c", x"4b392681f91be522", x"80e338afbe0833e6", x"f9a27c4fcbc6f81a", x"0263b801656d7c7c", x"9198d6cbe6ab5407", x"671bc8cf2e7a3334");
            when 14158124 => data <= (x"3bac5d8b2f4f72c6", x"15f1634868b442ae", x"392f0c0462a060f8", x"585634797541029b", x"83c0bb55390fa6b9", x"1249b12c070e1767", x"dc9dc1662e2e073b", x"c9b750a620068c1c");
            when 18249957 => data <= (x"2a158a6d02b17ab2", x"7b0ba43e0a2fcab3", x"cb1de9498c9a9249", x"ece4a1d915211458", x"5bc97fce5caeb98f", x"eb16bc00b5ed0b54", x"b4efd0a4c52a8850", x"9a35e36619bc35db");
            when 33581737 => data <= (x"6cb9863acd39e7b6", x"3a7f73130e61055f", x"679ba59a406b6faf", x"0c5a6655b52dbeaa", x"783a4a35574acdcd", x"c7e97369f3ea574e", x"902bff6c29b3efd9", x"f6ee49c50eda7466");
            when 17633606 => data <= (x"b09c1c6c935d4ffb", x"8a405eb4d021d0d4", x"323f553529741d1c", x"5481f91201970b2b", x"392fcdddcd8851f5", x"58ac8300e1027c1c", x"3a79d3d60d69d73e", x"792bf7ce85311107");
            when 12431125 => data <= (x"3b01b70e2db750d4", x"a97f3d5ea9904a29", x"c0f5597c6bba94ff", x"76a060b59b69a21b", x"652be6e11f8ebd11", x"d09be886677d664c", x"00112a4ab3611b3e", x"354ac5c6559cb97c");
            when 6488482 => data <= (x"19d4c7c0d4e94b2a", x"8ec35ff67d0951fb", x"05b8e74eb9711695", x"1e650fddd5707715", x"cb59941c6eb4e9ea", x"cb9da5dcfefa0bda", x"1bf30ad38f0b12bd", x"5a538c2724f9bb14");
            when 6491146 => data <= (x"52efc10fe31be2cc", x"f91a5aa727d26c7a", x"5d01928ffcf21f6e", x"21bd2b47688d855f", x"7197b0c8787ed834", x"a33b0fe7692912d3", x"7d195fe7615de67f", x"c19dfaf60874f8c1");
            when 4423953 => data <= (x"b236859eb9fc5fa2", x"af35cb613121a3de", x"61fe4bc4537e09ee", x"a2b5ff803349b4d9", x"17568f06afc56216", x"af0e76a03984beb9", x"0e545149e70b11a6", x"9f13663d24ef79f6");
            when 32258188 => data <= (x"c8e0244609dd37ea", x"41556972eccd6ba2", x"b7362da0ce8a67bd", x"c2f818bbc77cf803", x"527082bcdd0cb28f", x"5414133d80520497", x"e5b7431749ba85b2", x"1af9ae1c7e1127c0");
            when 21639998 => data <= (x"4623527b66a84c64", x"ad29483e3de721ba", x"f01df0632f141893", x"d9cc3c00e158fe49", x"ae3a94c2435ba6b4", x"cee9eb27cd5251c6", x"6807e9babb40d11a", x"e62b9b51721fbc0a");
            when 1374942 => data <= (x"d9194206afc01e77", x"672bbc79f31829e4", x"d3920a36d9d76ca8", x"062d2e3d72c11e8b", x"794dc185bd3aebdc", x"af6686c33de45267", x"1eed69597198864c", x"4548ed614d854ae5");
            when 2270530 => data <= (x"ee6f3e20977c15bb", x"2472d3fa254a0153", x"dfe3e8abf2206d36", x"f8ed0d7fe45e38e8", x"3bbd0e2841fa0f32", x"7dd1d16a6233e8a4", x"d6248763ef8ba45e", x"77627a17807aba37");
            when 23161797 => data <= (x"93280bfc1ce85afc", x"d1c205e44278f2d4", x"31492403680e212a", x"e2ef3dec669454ac", x"f0fbc7e2fa182cea", x"1a8b03397838ca44", x"eb78cd45f2ba17cb", x"3b2e61179383c1b6");
            when 25673804 => data <= (x"1371b459a89fa539", x"225fb84fb6e545ba", x"2b87195d31b91521", x"6ab39ed048628ebe", x"2caca969acd0bc9f", x"f73a2b7ff869a2fe", x"0d258c249c64f6d6", x"5eb02476a1576d22");
            when 33300752 => data <= (x"e7ec99c21042b50d", x"c0d77f0de10912d6", x"37a79e7620da095f", x"ce90121750a9668f", x"bb0df4351c3ccd89", x"175b2d7a108beec2", x"f171f44106147a41", x"4a662f9864aa1d07");
            when 21778707 => data <= (x"679cb5ee057948d8", x"fdf00f8aa08f750e", x"7c2646dd5eaeb97b", x"9b78b7d87b16425d", x"f32811a70ace621b", x"ba04471afa9d47c3", x"10712c2433933afd", x"49d00e4e98e3f7f5");
            when 33026727 => data <= (x"c223fc786c20f344", x"4124fc2916623565", x"c69bf3f36c2941ca", x"63df14db2ad1fb33", x"5ff88b6e1be881ff", x"c6818346523045b6", x"bd465bf8a0653b28", x"3c2e0a795239aac1");
            when 23184039 => data <= (x"8c9bd6c8b6f2bedc", x"e213519bce1cb1d5", x"10bb2789e12f1e43", x"47d3663b2e7988ac", x"0d26b8adb8e9dd72", x"c651b098637b1b98", x"5134980443b4aa96", x"d8fe40dde29879f3");
            when 32230157 => data <= (x"4ad025085f273479", x"6833d3ea665909ac", x"0952a58f246e4615", x"7457b89ae6e4409a", x"2c170ad9376dba47", x"4f8ddab802c180a7", x"1cdc2bfe4537f802", x"7662514defc72560");
            when 28352394 => data <= (x"ebf67664d38eca74", x"b06022b79a315e70", x"2562123ad7d37e31", x"71683b6beb8bcc15", x"5943b95aae57f902", x"f1503e47b7bc9d14", x"d0941020b6917ceb", x"7bda16eb86f65f5a");
            when 14249015 => data <= (x"f659741df96048cf", x"aa9a6442ba7f27db", x"8dc1d318eff1b5c5", x"2ec49600b88a78c1", x"98f3f8b411f627f0", x"54b5393fffb9e68e", x"a39dc692bda520d5", x"3bca4b5c859d40c8");
            when 16904412 => data <= (x"82c81cbb8f24d8ba", x"34822e5703352e25", x"8fd2777e8c5db12a", x"e0ffe860276cff08", x"d9c1bab858c7438a", x"d847820ff6a13b9b", x"4006ad314c9df642", x"f8c03eaee28bcb79");
            when 14512265 => data <= (x"725547d18035204a", x"c0ce121f8bbbd320", x"62d0117302d457b0", x"acdae7c79b197802", x"0f37bcd597c6e2bf", x"058ce5eed91b4bd3", x"01fbb9922fcfc419", x"87140d43890eaf8e");
            when 33605917 => data <= (x"c513d16ff037c3bb", x"dde3d366ae4d7c61", x"6b8a6d16be90e2a1", x"b4fd3d2de4c9d595", x"67fed32376003fbf", x"9310174f8bc668fe", x"374d3774a6ab821a", x"5c76675855822c8b");
            when 33171573 => data <= (x"1f2624f45d87319e", x"544c7352664e0ebc", x"1768118fd574290f", x"ead1f6cb30f6601e", x"3a0a9d67349980d9", x"a6eb070f35f02cd0", x"0800186859229421", x"e464a8fb08f5ae3f");
            when 3413573 => data <= (x"78a3f1240a4f9037", x"2f24b9b36c2e70bb", x"e7d98eba212ad7fc", x"3ead9232368e4635", x"0da4323334d1f5ff", x"636969e825f1ca7a", x"0ce2a84e01af58e8", x"2ccde23222ff1e8e");
            when 5995041 => data <= (x"349bc4e24f0d88ae", x"7900058ebb4b5851", x"8b712a52e3b3e6a7", x"69696b115d4d454e", x"93b41681954259e7", x"1a41dfe56ca5de0f", x"f8c09997a5fdb1b5", x"6b167805b261dc60");
            when 11056611 => data <= (x"d9194a03923db52e", x"52cad98f49950bc2", x"901fdd6a8688fcaa", x"826eff81ef9cde5e", x"657b5a3e8b687156", x"20dff5abbc21f85f", x"f8cba7d63ed9aff9", x"55743a5fa9bacf87");
            when 22631556 => data <= (x"4ee21f7a75513066", x"f5db62735be1c675", x"7c2360fb9b313abc", x"55cd03df69d2d72f", x"ef569f5ae82e37ba", x"892e75142d3c01ab", x"8cfb71bced20fa7a", x"95128dcf67e714ce");
            when 26070873 => data <= (x"fe2833fff2df6b82", x"bedee769db5fd30c", x"bf8b8f4153037ddc", x"36d7af76879c785a", x"1c9c9f1c59cde7df", x"2e80abb3131391e5", x"fef59b905e85491a", x"3e9b51abbedf72c8");
            when 26617135 => data <= (x"88baf78a76f6300f", x"849cd592b9a4fad1", x"492f06dea4ed2d55", x"c35e3e3eecc5f8f0", x"aa57912b335c6319", x"1114bb10fba6ac20", x"8c4b666f25091527", x"8bc52b051115f800");
            when 32743867 => data <= (x"837415246e846c01", x"88b2dc89eba3f448", x"fbe9dc4bd536e856", x"e18a3cc58fbe0a88", x"ca61edf4192500f5", x"7efa8411e1c95d9f", x"a7262301e85f8333", x"a2a03b704a406669");
            when 28475442 => data <= (x"8a16ae9694c3e1ad", x"1ae18caf51cbe7ce", x"0b901023782be913", x"5427990c9bd4f9e3", x"2b11eff14ce91283", x"ae3fdeef8346a373", x"48b8c204be2c3e65", x"80e42c12adcc9ec2");
            when 20573754 => data <= (x"f8f8c6589dacf70e", x"d4c1d3f76e7b1d52", x"d9c25ee7d4c543d4", x"478654f2ea92d377", x"5348100f7ea86c49", x"5e334d7b2e99a64f", x"36d1e2ddfc29b0dd", x"0a9a77fea244bd8a");
            when 14904440 => data <= (x"f73f28510abf939f", x"2bdc13f8abefd381", x"c49c43167b34878f", x"63f45d6ec5364e83", x"9008f682bea1985e", x"da401450df60dd67", x"ed20391352e43227", x"8e9b711134c5c7a1");
            when 7443429 => data <= (x"af20c8aa23c6408d", x"9ca866feb10be117", x"262d23583a72ca87", x"94c3cce9e80d8fdb", x"051661f2396b72fc", x"21c1ab4fd6a6480c", x"57f3c3394f17c6b5", x"d80d8bb8272bfec4");
            when 10386635 => data <= (x"2e9f4e837617f293", x"b937748b454a108c", x"6618a817f3d87772", x"dcd8ba1fb80c4f52", x"8c0356249b5df8d9", x"08b33f77749ab28d", x"76a2ce756524c5a3", x"907c53ec15ffc08d");
            when 22716516 => data <= (x"807c558e4a190c6d", x"f73ea9249ccc018d", x"02af5a4fb95fc81b", x"67aa844061641a43", x"f411f1e39c652b8c", x"db3913fffd1648ac", x"8bb94db097320c16", x"44327425e81e4949");
            when 14153265 => data <= (x"6b8fa4731241f58d", x"bc663071e4667665", x"29be2c0dbac90e36", x"5606f298994ddf6a", x"bd4bab38b1b4a402", x"b4a7a8b21ac878ac", x"6a50d2f13130e9f8", x"ca3ffdcf472d0d77");
            when 27113122 => data <= (x"04e7269f8bc2c224", x"5c87ac5edd1dd173", x"7ed7e728f4f11ccc", x"ce839a6e0ccb0049", x"7a32208b24660a2a", x"f5b6558f0f796363", x"06614b60e18dceb5", x"05da8f5ed08e905c");
            when 9409008 => data <= (x"ed897274f8131654", x"23b8c15bd3f0f11a", x"bc088435c534f9da", x"811f551c27fec7bd", x"605b9eb0245ee300", x"23de44864e041a83", x"a33a633fe9910894", x"4f1109c3ce09a440");
            when 23946531 => data <= (x"5283af89ca4bb182", x"2ce7288f0ad82850", x"3d2456adf074fc38", x"eecf69a59d64dc6b", x"26542b507490403e", x"193df2a7fbb35181", x"f7b9534aefeb9e97", x"2ed76d90b7e56533");
            when 4067172 => data <= (x"7852cbfbcb11b01e", x"8c5e23048dff0f26", x"43d4e6c062e19482", x"9d50c2b99faa62f1", x"9287cc3189641088", x"01853db76d46fbdf", x"607d22279ef5e564", x"1f8aa488f4c951cf");
            when 5869250 => data <= (x"9019bb6f88a38d71", x"79c0a76b26601c1c", x"8a76530fe735406e", x"44f15461349b60af", x"496bbbcbf4c8b4ae", x"9e87cb60dbdad30e", x"25d2abe6e9c616ce", x"ba92f243dee41fb0");
            when 18992122 => data <= (x"1b2594be38749993", x"51cf42e2bbae7e5a", x"80944396a6345159", x"3b56c7e37fccddb2", x"2d8c6cf2d924ee94", x"e1df13101aaad356", x"ab788fc6a6b0d8f5", x"6d8cb65ca91a966c");
            when 28033910 => data <= (x"9dc4d19c16fd1ac9", x"df16cd484218f790", x"acc0747ca5d2ab45", x"a0bb4803acbbeb4e", x"5f83000b871c0d83", x"07bb69570e8c264d", x"63b62df4cd547905", x"802340339052c098");
            when 25691625 => data <= (x"80b1a61155e18640", x"d59a34f3aae86776", x"e23a1fe154088bc1", x"9f1e4b943c2e162c", x"7025117c54f8dd8e", x"8256973223f36595", x"d28fcb3a839eedce", x"27906dbc401adfc1");
            when 2264065 => data <= (x"5ac739f1f1ad12db", x"4e60415062c5f781", x"218037ce61f345f5", x"4e7a7c491995d1f6", x"00bed10997bc75e4", x"4e4ed391590001bd", x"e8180e0f3377a31a", x"e88bfc324d3b4ae9");
            when 8817708 => data <= (x"78f011713ce1e03b", x"6d8748746ee73ff9", x"07c099c34c3bca7c", x"802b2a61958f6758", x"d3dc43a8b11930db", x"adf91479a9617c19", x"7fb46f07cc47e012", x"5a7d05e5fbd86a5d");
            when 20647307 => data <= (x"78dfd8cde60527f6", x"62bc3a57cabf6c06", x"5bcdb3ff6171df45", x"2382c46add63ab63", x"9a4f94a37cc9e70f", x"cbe0ff6fdda650a3", x"64dd7f7f95fe110f", x"a7cd78146dabaca3");
            when 29670125 => data <= (x"1f1cdeb9f35a35e9", x"9bfd0126d0660130", x"4f1afc6974500500", x"36c0691447898daf", x"4ff75c4c390bb093", x"6e6044f29d36db58", x"a33c1dea34eb399d", x"40c0b3b7893d29bb");
            when 32402773 => data <= (x"3c2c79c7fac99df5", x"da6d457c43ee8249", x"ac64ed81a532e308", x"122500d67c539a07", x"66fc8f4dfb0b7994", x"f386b4d589771bd4", x"d466e7db77db2ba8", x"e18b25bd1e834ce1");
            when 31591125 => data <= (x"a74041ce1b65c623", x"4dd30c39dc154e85", x"ab58f8afa67b6c41", x"4820e64fdd85a136", x"3b77ce2b75a56e6a", x"074f3c5cb4e65360", x"ec18632dd1a7efb8", x"e54405d9589b9697");
            when 1405216 => data <= (x"c0b90cb5d12641a1", x"e1c94e613dc456fb", x"ccd65760b380f743", x"ea039517ba7673f7", x"34c6e1dd8ed2b325", x"09fe29252cb57fcb", x"aa0bf9e9a0a7062b", x"67105e0cd1b0dd2b");
            when 3860767 => data <= (x"afa979d25a82b715", x"6634a196a0b8e49e", x"eb010fb933114975", x"a186edafc24b2de6", x"cc1ffec68da4cbd1", x"b94d1ae45faa7708", x"48da4f087881e789", x"f11abcc8c5cafcf5");
            when 17971430 => data <= (x"3d87dfd041f2755f", x"12805983bf01d33d", x"06957a1d7a303350", x"282dc33137024cb5", x"33ca66c02b121b3f", x"a6944fc4de54be33", x"6c78cfc1855487d2", x"2fd813b71aef42c7");
            when 20772180 => data <= (x"2bdf7425ae21b945", x"7b05e811ef349ff4", x"4f8cf4bcd32ac400", x"71bddc381f56e22f", x"e884cb333eb56f1f", x"1e7d1ea3351ca618", x"a1e2eb3d52f16e2c", x"ff85c26b46b1d7ab");
            when 15765930 => data <= (x"c875a83d05694710", x"8216700bde3ac6d3", x"cf31d58e8b558ec8", x"4ffbea8a2ab1ef97", x"7dd83c1773571f16", x"6f6fdf93b6ea1810", x"3be8a4751411e530", x"89e8c3ebbeb4ad28");
            when 32161461 => data <= (x"8d5d8174e1cbd684", x"d82ba2da169339a3", x"b4187514caa4535a", x"2f18eac214b457c5", x"4f2e388b577c9b44", x"98a0e74e0dff9fff", x"cea778990096713d", x"ff0f7b38af1c10cd");
            when 8914276 => data <= (x"562a233f03e1b299", x"2e6402f455791896", x"f8da1588c02592e1", x"6ba0dd85f445d7f9", x"96d8f493f53d479a", x"ee4ec38abb4e39ba", x"2173e2b2026d823c", x"0b8d84afea61e721");
            when 15133951 => data <= (x"4a132e54396cbf4a", x"efa773e279664228", x"52488fa65d8e4c85", x"0f4088b5bd36868e", x"11ed0bf38bfef04d", x"674c2ee2f1ccdb70", x"da9013fa8a7ce8f5", x"7d6a778c3ea6c3e3");
            when 5089346 => data <= (x"eb40b131add362ce", x"a68de9a2c85f7cc0", x"c7d49ff7446c0a4f", x"cc9d2d353e307cf3", x"bc8381213f201c9e", x"6ddca202d765bb34", x"67f0e425660cae95", x"7c4ac35219fa7298");
            when 28089941 => data <= (x"d8c870681916b34d", x"1322520f63a4e683", x"5a1c8d504ed48607", x"25da022f1515dd46", x"2c37aac023326501", x"ae84b7855cd1ddbb", x"c754fd14d36ba8bf", x"e8f4a3c8f55be7ba");
            when 1519611 => data <= (x"14a1ba6d0a36f61e", x"eefbfd8bb38850bf", x"44c6cab6cab3919e", x"77201ad929a953a4", x"2b3ae72bd65abbb5", x"59b7070d27e12a3e", x"3bfe6efc7bed4881", x"08ef081f36738c6e");
            when 28453882 => data <= (x"5bf272c36ae70b42", x"93874d926d22d4a8", x"f3cdd6766a7768c6", x"7cce22d2647f6e71", x"9e79ac83de309237", x"5ce0a0ea2e726546", x"ef2045620d74b8f8", x"2e59289ace82e049");
            when 23229718 => data <= (x"389048bc5a4b3669", x"c183a8c67a429927", x"d7d4aecd6820a6ae", x"37cb2d220137637e", x"038238b7e67a16d1", x"d49b05909fc446a7", x"ad78509a181b12f8", x"98eb602bf62a51c2");
            when 19234845 => data <= (x"c704f46861e6a889", x"2fb94dfa02a5e3f7", x"aa5cb6542bc9866a", x"681ec26df404c3ff", x"129eeef83eaedb9e", x"35e85b54a5e8f207", x"729b65dd742261f1", x"eb94117875c0eb4d");
            when 16368873 => data <= (x"0a0023616fe56ba7", x"fc32391a62452040", x"24ea196b65f23d7c", x"39f85747ac199f6c", x"50fd28f3cbe02e07", x"3a3efa870f07a8eb", x"e8c66b394556af9f", x"6f0263e5ba732308");
            when 18067312 => data <= (x"b4cdf2b6fe3c99b2", x"77086d692ca3dc49", x"7cc43511635f280b", x"c4e8a9c406947e95", x"9fe05a5e3e5818af", x"22ef7d9a81416a9b", x"6e97c7e5f916ab7f", x"751077c6a30937e7");
            when 14149998 => data <= (x"b2d678bcbe3f0aa8", x"ebfbe754ad244d7c", x"e3a604ed1602d67f", x"b7992768e9b8d5f0", x"653d203d6afee875", x"ab41ee20610a3342", x"4b57ad3b6302b275", x"4935ae7eeb7b89cd");
            when 28438137 => data <= (x"008993b81f45851d", x"723ab541b89d7c99", x"5247f8fc18481cd9", x"ac460100046ea2f5", x"d65f655e133d875a", x"7899b4c0ac693e44", x"92daabad0ef6ee95", x"c5eec442055a59e5");
            when 30497197 => data <= (x"9c07ed62e174328d", x"4843ff51facb639e", x"07e38acacdef3a61", x"142da16071cbd4c9", x"d943eb93e75fd4c7", x"91613b29df2c5428", x"f9f00fedbf95b97d", x"513262f0b1dd8927");
            when 30649193 => data <= (x"6ee88fa500906237", x"df9d19ef207b5af8", x"5154dc17a87a3726", x"95cc033bed8bdbe6", x"e3d005174a6f4679", x"1b0e1fe3c62865b1", x"c2541a97ca5d7952", x"a3109eea772ec3e9");
            when 7573699 => data <= (x"148f9a205943b54c", x"e1a2f2a6146dcf18", x"3ae54f8dd5e42c2a", x"3c2d4756eacb1121", x"4ea1f16e0b0d5d76", x"116da1d28c8acbef", x"df5f64c436d67f99", x"ab86426861160bb9");
            when 712440 => data <= (x"bebed1473fe166bd", x"2f4f5ceb46334ac3", x"8ce5a426e04f3e8e", x"d0680748ab16cc59", x"62670c5099b3c72d", x"433d0b5f047a9031", x"6b88529fd8a7e73a", x"5be719f26fdb6d89");
            when 933679 => data <= (x"4c23604412b4a07c", x"a9ddd6c307de20dd", x"1adb1862a2c69b62", x"a2fae3e9a0bcbc07", x"b546f27793ad666f", x"14ad6b1640909f9b", x"6f024b7fb66587ec", x"5dd3d85d3d4b6595");
            when 29620037 => data <= (x"8e6f907f1a209d43", x"1b1cb985341164fc", x"7f6fe42eb8009b48", x"adea345a7dda66ac", x"80f65ae4f0b72170", x"506e0f8a7dbb665a", x"2f148e377c5b481f", x"d8afecc92d6228f4");
            when 8275158 => data <= (x"61737495bc2ce30e", x"722473b7273ffbe5", x"4fd305565bf09910", x"690a389af0bf2740", x"03438fa4680dcf3c", x"88ca5a86619527d4", x"6701a63f205547db", x"54e66892f972615e");
            when 20841053 => data <= (x"0cb9a64000a83fdf", x"72e1f7125084cbda", x"519e6bee7543a841", x"8ddc87410c1fd23d", x"7d9065948611ef70", x"f95aef5507ffb274", x"5c973b4f94e77111", x"3a671c9f493990a5");
            when 33853873 => data <= (x"d7ba03c84cdc8084", x"0f8c6dca0a1a7bf8", x"172b8344ff9c2cf9", x"dca85fb387670a0c", x"1b47efd8e2c350f6", x"18e02cdac8a0b2a1", x"4c6bacbee1085768", x"65db0631d10b2862");
            when 16248549 => data <= (x"0838cd9f9f8b2ed2", x"ee2da6e0c528c8d1", x"b3bf146801286196", x"ce929bbb9b088ed4", x"1ff5bca496483280", x"2df8fc9f0a4d2540", x"30dbbd35fb03f4a9", x"23aca716d5b118f3");
            when 19624824 => data <= (x"668ad35edab20ba2", x"19db137cdd2afd68", x"9af391aca6ce3978", x"51354836f3c39361", x"a0fd15039eb95649", x"41f15c95f9d78659", x"8953042de4e06d19", x"b2d941dd6376f52c");
            when 30052904 => data <= (x"48b166e6152d7304", x"df47d94084e2c39c", x"e9d8ccec6ad0d3d7", x"996ac1582ab9ff85", x"553370a45b68f893", x"961e5242267404a3", x"5c9711f8a77a7ad6", x"fce0ad6dbc64df54");
            when 30867180 => data <= (x"584d8cdfed39eddc", x"5d682634b695b243", x"97a39353ad9866ef", x"564495e6374a3655", x"4b95196c66f7cd9c", x"d5f6315b9378a904", x"aafa13e6896168af", x"3369ef68dd2919e6");
            when 17769196 => data <= (x"3b886d79778ba096", x"77adfd7de736f1ff", x"5438748f0ed83f70", x"4641b415ea25820d", x"cdf5432f788de2ad", x"ba76f92e23d46a73", x"09edfbef97ddb903", x"38826d00f2028d76");
            when 17925097 => data <= (x"704c626d6eb13772", x"b4309c919d02a814", x"b690cd8cd2363616", x"5111c674c2f8f078", x"189ea36e167853b5", x"f8ca1c92ce1d5654", x"812df2c8a59fc3f1", x"dbff985e7da71991");
            when 33704530 => data <= (x"ead2aea122f4bb07", x"ae0044564de490b1", x"af13ad70bb64c56a", x"c01e2cbdfd5911aa", x"3f5190189c9522d4", x"01918750ce0b3df0", x"54e53fb8f01352d8", x"3e4a7f7b3f4e9b27");
            when 14037142 => data <= (x"df02748a52897e83", x"05f5237ec4788e3f", x"cb46c0f4ba4001db", x"889f40640219aa0c", x"3dbb76dec6929bef", x"78ee3ec293803c7c", x"945b202663789dee", x"47bf8c77518d13ac");
            when 12710548 => data <= (x"01e6707dc72b2266", x"d35064c82a118e1d", x"793143f86bfd43a2", x"47f0d0609bf5fe0d", x"6171af9f3495e309", x"d23eade171c77e59", x"c2ff5eade5db7ed0", x"94216de28dd00de6");
            when 23604352 => data <= (x"d55ed2a66ab3f6e8", x"570d1049b454b03a", x"d7ddc2d26f0d66dc", x"695c1cdadecb3ef0", x"a8041b5a87c3921c", x"4e043b7b4d75dce7", x"d52af54e526cfdf4", x"6b2c74131e58c635");
            when 11591471 => data <= (x"2ff11aafa7219a59", x"7abbcc5861d6e879", x"be51cf360e18a242", x"3888a5fc4d243f8f", x"9a88bbe268fc9c4c", x"25dfc398367089b6", x"71bc925bbf0c2bcd", x"a941c34aa69dc765");
            when 30528834 => data <= (x"9d67872cb7ece3d1", x"76b28bcf2facbf46", x"a3c5f4f66b65293b", x"e886b912985fa26c", x"e37380becbfa8e5c", x"216a6bccca056d54", x"8cd3263107e505fb", x"41e9ba8182c7bd31");
            when 14113903 => data <= (x"badf028ed285c455", x"25ac0af27eccb164", x"a15c8ac29fd07a0a", x"72e1d1813756a9c8", x"26d983a4b7be3723", x"9405cddcd1423ac1", x"95bea368a151ee62", x"88ef241f513f6d50");
            when 32995872 => data <= (x"2cccd8f542e7473e", x"5e7971cd42c49f5c", x"cdef823911d0ffad", x"b079fe08ca466081", x"775502a3d07af146", x"2e88bd16150c92e8", x"656a15df9fe3cdbe", x"9c2366b242b6f645");
            when 27169991 => data <= (x"7d8a0b1b21b24ae5", x"c52bfa634b6ddedb", x"3c74c37d205d956a", x"5a759e7ea836a280", x"e3003684505a0248", x"d346c89f66eafbdf", x"13e411a888998369", x"de842c4245c4ca01");
            when 2169584 => data <= (x"1e54fea8781263ae", x"f4facb11400b0fa6", x"429c488b2a6c7f8c", x"d6c0630ebaf63095", x"584308bec43469d7", x"5c2b52c681a88bab", x"29af0121b36b2234", x"4acae5be48055659");
            when 27209668 => data <= (x"cfba87ef5e1b15be", x"db8c5c4c5b71ef27", x"2dcbc7c5b53f0e6d", x"93a9b2e7d4642526", x"5ac675728636beba", x"d15a728c867774ad", x"183b65fdd38616d0", x"c91ad7e6558e0b2e");
            when 9780940 => data <= (x"48658bfb10156082", x"b6ed1906dcd8604d", x"cd12d2d934aa2265", x"c2a40bb59a5d8c07", x"2573709846d8154c", x"b9fcfdfb29cbfc24", x"a1f0849f349cc01f", x"3f11d8afce1b91df");
            when 31204505 => data <= (x"ee84d08e9f07d86a", x"7004ef0337420c71", x"41c2c493fc655fb9", x"c577a491b03e755c", x"1e4bb36275415a58", x"22a29397c351b990", x"f780243efbf135d1", x"bf58245e046e6727");
            when 32280774 => data <= (x"8a5bb9b6c22e31a1", x"07f5476e93f9a628", x"ecc52fbad029c012", x"cf75dcb115525fa7", x"2a054a0391062274", x"09965410e7d997cd", x"5d4094edb0a1c092", x"0b8871c151dd03c6");
            when 19451008 => data <= (x"e49485bb14b00e91", x"99dd4d737b6079de", x"d8ae921700a59537", x"faefb86aa9ed524e", x"acd10a985c4f339a", x"6d67988784e6280c", x"ab01a40b13997e67", x"441fd6e0ca32a78f");
            when 1221275 => data <= (x"597d9fc8561629ff", x"d3d3532998b80128", x"09aa03ddadf3cd5a", x"c09d41bc6049073a", x"b5e7990fcb8c6eeb", x"0d1c5f044c989a79", x"a93efab1f6fd8943", x"64cf85f08595fbc8");
            when 23169679 => data <= (x"9c081e56ba0b3b47", x"bcb791e75eb4bef1", x"c07523de62c0affa", x"932de571f4278cb7", x"a4b3832cd8af7306", x"cef1a3ff0b67f624", x"778ef377830429cf", x"d71340870a52a79f");
            when 22188419 => data <= (x"1ef3f02bdaeb447d", x"7777bbf12c7fce20", x"8cef366f9cf15156", x"50f2505eb8a712fe", x"edbf915c6ba6385d", x"5f541b508a316310", x"3ec46b776b982ef8", x"0024a1b21e38eaa0");
            when 18259572 => data <= (x"e93ae756c470e199", x"aa0f1b80a7efa772", x"b85bc76a889decb8", x"95d7665bfa957e42", x"2ab23751e84fd04d", x"cc29531ea4de39c3", x"2719acfc8b2f75c3", x"4e18d384a10f9e7f");
            when 15319327 => data <= (x"930d8a44370cbc96", x"e0e9f9fa33fef7fd", x"cd4eec995f601836", x"1494c78a5ade4f23", x"e1cef2eafbeebb7d", x"ac540501f2faa051", x"e23a64ba9dfb582e", x"debf862d98f7cbcd");
            when 33791088 => data <= (x"ed1ab020433fbd9a", x"8be523cf403b116f", x"5805ede895ca27d8", x"076a36bf03e74d9d", x"ae860ddf15bc5a72", x"30f0fa48a4277d9c", x"3d88adf2b412a299", x"37be276ab7db27d2");
            when 16695666 => data <= (x"c917543875fe8838", x"9ebd992724ad0e4b", x"05ce9f157090c343", x"56143236512255fb", x"ea9a289b84c29edb", x"c9e94d1c3aabab0e", x"529bcc289e62a339", x"28ca475b3157ec49");
            when 1866900 => data <= (x"a18b9888652b29a2", x"e2afe4b93eb4e006", x"7e2dcc2b245ac8f8", x"52ef0d5f6ad60f96", x"965399e875c89143", x"80006e070a39b2e4", x"942868b0cbbfd8e7", x"7285dfb6082bffd1");
            when 26743019 => data <= (x"e39d30882ab09a7c", x"6727f69d836f1821", x"5814dc3e114c0981", x"83416f9a943f9798", x"070bd03dfee37e09", x"641073aa21dd55ad", x"60e94e0f9947a7a8", x"9c2d3def3ad7c94f");
            when 9072092 => data <= (x"362d4bc75da492df", x"d761fdc8fc218a02", x"6ad367ce61b945c1", x"300d771a8df43f89", x"82d93a3be422a5de", x"006e0b7a87dca54f", x"14b104a72cefd56e", x"c3aabfb8f2eb6f3a");
            when 2610185 => data <= (x"855ce2b7e50f3070", x"ed8d1bb44bf9f9fc", x"79e747708879e545", x"19eb3551ac35948b", x"80684f6e97cfdc7f", x"3e5bfcaea0e9c13b", x"e7d2b8ea237a9c29", x"505508e442fd4fef");
            when 21302386 => data <= (x"bb5036d01b621d41", x"131fded6ec27500b", x"69b39fdf9b8da6ab", x"3a44ef447b144268", x"97961df55105ebf8", x"29a1f8500c08470e", x"5c0887a7244beaf3", x"097676bcfdc5fc7a");
            when 28481880 => data <= (x"13a8acbd59e4c2b4", x"d3a2245a55688d8c", x"4db29b04da819109", x"e7e81696984f01c7", x"07802bd047c8d5c6", x"940a1ee3f7351549", x"26e8fd25852339fd", x"8f40d9603e1f0f63");
            when 26029902 => data <= (x"fcde33e0b7aa04bd", x"75c7d2d341e361b0", x"b6100b91b9ed2de4", x"cdeff9321840e571", x"10f7b17f68a6ee5a", x"375be79ca7fcfef4", x"8537b0c19be06f65", x"a5b879491376da6e");
            when 5197570 => data <= (x"29938e4a42c159b8", x"cac8d5afbc1d15cf", x"a70ad70fd09d5ba6", x"79ec7f46b1757d3e", x"50a59da6d693e833", x"211e53a89f3afcf2", x"090a27dd4cfe891e", x"d7891c7c240cf663");
            when 15179419 => data <= (x"cea4823c71923336", x"a0cded038677490a", x"450051c4ab230cb2", x"47b6928017c47224", x"4fba1d7279f2e1d7", x"0661588ea4e3f5c5", x"2e8206c9e2a8cfea", x"3afe44d6c968199d");
            when 21284795 => data <= (x"429a43c5109b13e5", x"a75be2c35f1ac3e5", x"08614c9cbe74d40e", x"1d42d9fa8ff63f6c", x"41cf9c1f885eeb3a", x"5760c7e623b02690", x"fefbea7d1b691fa9", x"ac7fc04ac3c3f527");
            when 20302005 => data <= (x"f92185fa5a1dfbf4", x"175b318e8337571c", x"71d76fd7464995df", x"dda0854ccd58f192", x"d031dfda6cf230f8", x"feb28c5efb49295e", x"48cca213199b1cb7", x"d25a69e32451bd61");
            when 20996366 => data <= (x"65bc8783149aa963", x"a3814b438475517c", x"36f0802593ba4057", x"0c535aff6980c0d3", x"d384ac034f4d8e32", x"c28c9c5ce27fce9c", x"3762833b2f3565cd", x"f603c986e352b5bc");
            when 17503227 => data <= (x"52704a76bb9d5bd7", x"475c95820fde0888", x"f70b3d5633ffc477", x"eea55db8d67027dd", x"6a687f6a9012b177", x"8e11d953570482f8", x"c06ed8626091f852", x"9a4f0ebd49882330");
            when 13824028 => data <= (x"a36a5422b76764f9", x"9340f69ecccf70cb", x"cb944027d37594bf", x"710fd6ed79dd2be2", x"3d88a13b0cb39673", x"fe412988f82faed9", x"3b7b136fcd48888f", x"cceaa1153df0f6a7");
            when 18600838 => data <= (x"921e9ac22f9c1b07", x"8ee5d90eb3a3c477", x"6cf7ca223205bd4f", x"c78e3deb99818816", x"ab53b26982cb4300", x"c77dedb5111e821d", x"90c5c5d8f24a369a", x"259866d036d8508a");
            when 1857232 => data <= (x"4d95fb849f063648", x"6272c20164d041a0", x"14aeca153d691e82", x"c67bc9a189ccd1dd", x"8ea88cc665a6c900", x"3cdd56841d0752f7", x"fd9ee1cfe2a4ba31", x"2fd77c5b73cd14c7");
            when 2109752 => data <= (x"7f519f9651013e2c", x"5a7025e8ee2de207", x"4b457b80e6745ef0", x"f7b7838eb6f95dd2", x"7e4dc97992ea4fee", x"b7391f15b38b7d22", x"477fd296c685097d", x"51ca5dd286dc869b");
            when 33124014 => data <= (x"ad234645fb54c390", x"6cd34a0d1409e869", x"5665c82306b82028", x"5b18a8f9bbbed25f", x"11cbb0b1678cd030", x"0dfe5f88e7cb87bf", x"0171f89af9cf34ee", x"af56bbd852e20aa3");
            when 871600 => data <= (x"e00fa0b7f8ba0d26", x"afe0a03fae44cffa", x"911c30b0c31a261e", x"2195640f9a5a3c3f", x"6a765d868fc37785", x"f48a146a94e1ba3a", x"c465fa390f8e383a", x"fe7141cbe7eb4a88");
            when 14960037 => data <= (x"60af2b12195c49b0", x"9c9e7acf96dfb391", x"8cf179751b89e38e", x"7ca72dfa9e3b4a33", x"f3ce26ee9b42fc71", x"6dd5c427bdd3e11d", x"fa0b9f6632469bf3", x"3a5034bc0f8151f4");
            when 19093143 => data <= (x"c2db77c4a315e45d", x"069a3c0413d2c42e", x"b15a31ddf4f9caa3", x"035bce9699f28ee5", x"99b063927e098570", x"105204da5b0efea3", x"6bc6e17e73d6f63a", x"b07fb89235f06bae");
            when 25046997 => data <= (x"e559b88def6c8ea3", x"f8c17f3fb4959415", x"9a92a5fd9bd8db28", x"6084a57591f84d6c", x"d16cff72e5a86145", x"2ae157306da539d3", x"ecf01427d52a463f", x"ae323c4fe63004f8");
            when 1857274 => data <= (x"bb7620d8a1556e57", x"971537d769539375", x"5e8695ae46c71526", x"7524d7b1c26315e5", x"25e2b0b5eeb83318", x"ffae2fbf00139b5b", x"1efdcdece93e7eea", x"c8b2537ba07703d4");
            when 30422287 => data <= (x"02f594c74fac0bdb", x"56f8af314215f61e", x"017850ea52a6a475", x"acf434d2f7ec46fe", x"f1d2be575411d303", x"8f25c86f454c5ec3", x"abb5f823256df604", x"7505a576c903667e");
            when 22430684 => data <= (x"49cc4fb7084a5d42", x"ddf00119a6c2ffd2", x"13771a3206019788", x"63091bd18b791041", x"3f7f28bd21d7b6ce", x"b8194b0b97f5084e", x"f44c36062015b43c", x"f5e32a674fe24efa");
            when 18382296 => data <= (x"234282f72a260958", x"8dcc5c3f967a6c89", x"f9d8cff41b06db8b", x"e445efcd81af4439", x"a111be790717fb6b", x"d0d660eb932fd636", x"d142fec6b648bc89", x"4182d366b5cf54e0");
            when 1314927 => data <= (x"2d4ca001797f368a", x"242db7a1cc9e9cbb", x"90b57e9c639a28f2", x"7a9cab56297521d6", x"93c8514593dc779b", x"a20d20e56b08a775", x"f25e3997a3b63e37", x"793c5c25a3286328");
            when 11962520 => data <= (x"c267189e3328b68d", x"232e3211bb6f2b72", x"7e91ec492cd58afa", x"d27a3749ca08acbb", x"92ed8240a3977c3a", x"32c92e8beea46a94", x"3a089a6e02908175", x"cefea6c6de75df70");
            when 31705942 => data <= (x"2531e9cba1e0d09d", x"db72c10e555df08a", x"0c944aebab1667e6", x"6e471d72b89ca73e", x"09f533cb1d1c160c", x"e4ef317e58d75fcc", x"e5c8801529da9a83", x"802439865a5ffd8e");
            when 19120636 => data <= (x"f1a6a783c5b67b5f", x"79e14df029a97c7b", x"6d40997a9dee4b29", x"fe82ec60457d8088", x"f2eca07666578bd2", x"aa63395939c2e2ad", x"ac565eb92e53729c", x"e4d74201c82d7de1");
            when 11872570 => data <= (x"d972533ce5a2b6ba", x"ba106e7d58a56b50", x"26962fe61745d5b8", x"5d4122d8a1317c7b", x"d344d268bbe45deb", x"b8b3fb2731183dd6", x"053bed75f7dcd35a", x"0f3d0ee8e5561c5b");
            when 30695046 => data <= (x"6a841b0e27bc39f2", x"5a8fee2fcd6edbdd", x"6680d8ad3fd25c9b", x"b835a018a15b9bd0", x"1ed7f03964e5b4af", x"f0c2dc18ed214849", x"ade08ebefc09b21c", x"5845a365487d1ad4");
            when 31642453 => data <= (x"fe557afd08128673", x"c3a1eae4ceadc4be", x"14260f47530b381a", x"fe0f45031a117ff3", x"0099e8f34d86c1de", x"b354f2b59464c6a8", x"056715dd60d5d438", x"03fb64d7f960d7cc");
            when 19302275 => data <= (x"bc21ffe224e85682", x"e3415535da7d5477", x"117b988bbbd8489a", x"7bf7e91066f9bbf7", x"4871d514513e0a06", x"cf385aa03ea8ffb6", x"1e3047acbb66d106", x"954e44e74ccbc7f7");
            when 17959859 => data <= (x"9c20c93e4dc568a0", x"97cc64777b0e0a16", x"5841c167d597f2d3", x"ae0b2fdc07dd54bd", x"3d8249364e850563", x"2b471aa0c29581fd", x"7a132f999efac813", x"bfc521cbc2b34c82");
            when 2891594 => data <= (x"6220f727922ffe83", x"fad512e844a4cb7e", x"200d12374ce91271", x"46ad66bac763519a", x"d9587c0166c30340", x"b8d4a13732adf9b3", x"490b72f226b3f0e3", x"ab5d6f1b6cdfe25a");
            when 30170601 => data <= (x"c935832cd8a174cb", x"425b6380934996fc", x"938af2c9a4934b2d", x"bc0cc38f0aed9b8c", x"d2601c961dcc500c", x"52cab94370952b7b", x"b19f62e4a7fa3a92", x"a99749475ed7033a");
            when 33032338 => data <= (x"39bcd8de53861b33", x"ebf526b0bfe40081", x"bbf74fddeca47d98", x"86894b3b399e9a62", x"d53918fd3aec4dec", x"dfb2be053e80c38b", x"852785a14256ecfd", x"8e468554fcc4f85d");
            when 4985717 => data <= (x"0ea20c4379f3dce5", x"7e39805186ec4fb2", x"de11f1869faba4ac", x"e10084798b858989", x"c2866c345fd0f763", x"558c3303ba9c4206", x"09c640f2b0741281", x"b2594d299db25877");
            when 10211208 => data <= (x"5da4243a765fbfcf", x"3e5591bdb7c3ddb7", x"6be4dae061a80065", x"88834251990aa27f", x"8281ae228c448b86", x"d7cc36277aec61cd", x"79e3d75b8e4a6f50", x"a3fb92ac7cf48236");
            when 32711938 => data <= (x"f1b7b066c341aff0", x"3ae38ae790f26749", x"69af6122643a31fe", x"2e72febb0decfc8b", x"d9c9f8ace73e5ca9", x"44e487ba105ae7fb", x"56eb58e738849c2b", x"6281f4be41dd4651");
            when 19332115 => data <= (x"44e917d546ffaa8d", x"3f2b2864bade268d", x"84a9899b5313b3e6", x"13abd671545b391a", x"bc38792667253729", x"67352dd10cafc961", x"b5cdd37bc191b80f", x"fdb13202dc6e1099");
            when 428751 => data <= (x"0ad11cd09bde8c7c", x"020492cd916d42af", x"6ed5d9fdb5bd3a57", x"2d16e6886536f271", x"209f9f273019cdc2", x"f9e8b991eecdc16a", x"64e751a8d9c9b941", x"72252870bea5bfe6");
            when 11534937 => data <= (x"f93964b21d969d54", x"1be93fd59d526831", x"e77a8d23bfbd64b3", x"f66a3422a6ffd9e0", x"9704570c0a804f85", x"35b968ee6e5263f5", x"c89fcc87750c8571", x"2f14569447319677");
            when 14596304 => data <= (x"e387830ede367cfc", x"569f2f424034e64d", x"ca26371a9c92cbd9", x"29746654d8e2f80b", x"80b0931f67d34d7d", x"b923b9189ba3a778", x"9c9744c2bfa2f45f", x"00b60848e2d95d70");
            when 4391878 => data <= (x"0d96294727276411", x"9908936c69bd0108", x"c7f5c0efa743e9b4", x"a3ff7d1b5ef28ea6", x"f520219cb6d15ced", x"56ac0afe73b41597", x"e3fde764a2cd71d3", x"0e5ca7fa3fe79aa8");
            when 19726182 => data <= (x"5cc3049942478270", x"fe83a36c4b584197", x"9c6f6bfb1ff2b174", x"33237d01b7a13c10", x"3e908a884d58c7c7", x"a485a517769c7fc1", x"be69ef3ce027c590", x"0ae9bcaa7a79303d");
            when 15003724 => data <= (x"01e0425e5c2211d1", x"e9e636652f0b3fb8", x"54238c78a1cdfe79", x"7ed94fe398a03f98", x"04343fc41fadddf9", x"1512299906b11cf2", x"29a4fcce80e0523f", x"2b35981190accc2b");
            when 24569320 => data <= (x"980f0e007a8268e7", x"bf408484cd3e469d", x"07030a7483b573cf", x"033335234ab40d69", x"ac1ae9cd9ec74e75", x"57ac47740b195049", x"659a3434d94afa63", x"050891011497040e");
            when 25476575 => data <= (x"fa82e92f812333ec", x"16da338304692bc0", x"510f43549558dcba", x"38a7a6432b4cdbd0", x"0cc8194f248e5aed", x"33cb44c64b2c58cc", x"94848597ec49e8ad", x"6106ded194fbd941");
            when 8132336 => data <= (x"f419571c774b2a38", x"1967bf671bee2c78", x"af7387d1add93dd8", x"112281da9083b2a3", x"e1477ec200389708", x"d9efe1090aa866f9", x"fc76de59aa9d52f1", x"1533844887121b56");
            when 26160969 => data <= (x"810e7fba960e3d95", x"e495c7f04901a40f", x"5ffeebb6932c0c76", x"1fae882366397c5e", x"5132bbdd5fd23b6b", x"2af244564818fcac", x"79f1b87b00e698e9", x"81b37f9c36b5c218");
            when 8844388 => data <= (x"c9bff97740bd52d3", x"cfcdf6f95b2c8633", x"d5122321962e9453", x"9aff65624221ebf2", x"d123ff86db296ee1", x"b1c28331bce1fad9", x"e4f3f352196c44d0", x"3608d4b9a876a942");
            when 10730620 => data <= (x"afd59656ead582cc", x"210621d8afbb0c2a", x"fcc7c4ec95871553", x"00bfbe0617dc20d0", x"becf3511c0bd95cb", x"dfae7a3b43b92ea0", x"a032f69d657bb3ef", x"c0312b986ea2e6fb");
            when 23383323 => data <= (x"d3761cc1708c0d5c", x"218ab6126ed640f1", x"dcba44c277f6cd9b", x"9efffdeeb968d485", x"b403029f4c159f14", x"f302b54c2b17301c", x"5e215e2b4627cad9", x"4cb8fd062cb5594c");
            when 32865169 => data <= (x"3d46f540b66c339e", x"8c9e120166490c90", x"24727538836326fd", x"9027458d436b5eec", x"80a433926e0f8612", x"a9be8662391ecb0c", x"1c2e851f6217a0df", x"2838de729e58e8aa");
            when 12463869 => data <= (x"8780839abdea77dd", x"a127ffbd1993b8f7", x"8c8179c4d4141f82", x"5e43fb832f54e73e", x"47f2cfb2dd78f514", x"efb6f29020fe60bb", x"2408834d392fe4db", x"0aa800dce04463cd");
            when 4405712 => data <= (x"360014c45080d375", x"5656c00923282d9c", x"25ae7b7518f1e21a", x"e5003613a06d40de", x"24c2d0cebfccfdad", x"2c7f2a953b900cf5", x"3114bff3ccbac0e5", x"310fe8b178c5148a");
            when 28254247 => data <= (x"60b9d8eac419da89", x"c662148a7db99bce", x"b278b0805743303b", x"5a0d3d7d6d5225e5", x"d262f41bd34b177d", x"0961d915d7b7c351", x"3d959e791f8dc415", x"47b28bbbd1e1a32a");
            when 15118986 => data <= (x"dc65eb9079269ebd", x"907d7cae2e529536", x"097a10580d62d97f", x"52ca3b04c1055c1b", x"9cb0419dbd908c1d", x"b99e33de33fbb0f6", x"d8894abcfd22a88b", x"756b8635219dad53");
            when 4504637 => data <= (x"5dd76cf2807c7145", x"8a482ac418f37a85", x"8760afe2e44d2d24", x"a48bd793962a1395", x"591e6d01c81ff954", x"6a68ff228ebd3e25", x"c0b9d96d0cf0a095", x"29f11c5ee92aa139");
            when 23513788 => data <= (x"b724e5629472f30f", x"cf6abad7fd70c4fd", x"85dc697dada55dd0", x"e37fd4dfdfa423d2", x"db3180ca267e97fc", x"8ee78f41c9759ab6", x"2e34601268c63fc0", x"54ef973800e8bb13");
            when 22705851 => data <= (x"c42f2fa2688b5154", x"854b34887e925e8f", x"fa50ecb08d9785e8", x"508bc86e4565fc4a", x"b06dd22975ddd546", x"110c0eba55c53829", x"3594fa28d8b47b1c", x"1271e0e1c86aa29e");
            when 11338399 => data <= (x"d0d7fa4abc5113a7", x"8b75f5e2adc6eadd", x"7ce0e2019c582b09", x"a461f3e2dbbb64bf", x"bc5eba9de5a01b43", x"bc5f81561dee3986", x"b7b0335f2ebf85cf", x"0b8badd0bdfdaae7");
            when 7944303 => data <= (x"6be1a8a67658a8d9", x"71e469a004869d32", x"6b622c6d59fedd3a", x"fb69de074cbe64f7", x"321b67bea406a51c", x"788e7067324fed64", x"ed54f2a85d2e343b", x"825da8084d97d02e");
            when 5857315 => data <= (x"5021768898783767", x"ab03335a0b5a666f", x"28a0a8960ba22378", x"e83a1425c4d3155a", x"15c061a185d64480", x"33a915e395e82818", x"5d219072243c1eab", x"176b84567cfc0a5d");
            when 3179967 => data <= (x"a32d3766b9609713", x"b5af49a6286619ee", x"014dd8914123e12d", x"d361916ffd95f5da", x"6a25d5d884da0f5f", x"5272ec6285bb1e66", x"d621f06a56e4b99a", x"603a45578757294c");
            when 2195976 => data <= (x"adb13422ae265f21", x"5ff6e8d517f71997", x"2994f09ac27834dd", x"64be196c81400991", x"13abf74d9717633c", x"0b877fd0cb27a92a", x"3af93779f0eb59c5", x"178bc4c9e43962d0");
            when 12224004 => data <= (x"653703ff4f13dd5e", x"1702d0bfd036ec1f", x"a79d0f0af12dbbc4", x"736159f73f56fa3b", x"1ad3340f9673e50f", x"bf62db4df7ee7aa3", x"b16c9c68dc7aafd1", x"bef2723a1ebbe0e1");
            when 3453756 => data <= (x"d6a53d300c6d8ea5", x"406ca3e645b502d0", x"035838620cfe61e2", x"aab13e97cf258a56", x"37e60314fb092e8a", x"635f9741efc1fd83", x"e7347465e83e1547", x"f301336c7f26a6c6");
            when 8003106 => data <= (x"dcd8ce3a33dd66e2", x"c28bdfa79d551e37", x"0a445802538f2fb2", x"6804bb83e36ed077", x"dc303c9adade7a36", x"cbcef1cdb1303c34", x"39effb4b14a56f90", x"2722f726bb752cfe");
            when 31532599 => data <= (x"2e6ade678b54e799", x"88bb8d72b83e189d", x"6cd4b643bc34b4c2", x"4efcdf544bf51d69", x"933ff741f9e3785f", x"47be2a983ae27de0", x"2329e13661ff485d", x"58e9b998d8d59d8f");
            when 4125318 => data <= (x"ff0681e20ecdcb7c", x"1a8a562ad6ca7cb1", x"4e37b9d50fada791", x"accfe5f5b5c7d785", x"4bcbbdc397b35069", x"fc5ad504017f9470", x"ad8d4a6a5ecc9ca7", x"f52ad158f90562da");
            when 23691135 => data <= (x"fa2cca6c7db6b19c", x"f307d016cb5b3dc6", x"aef6f7c2e7ed25d8", x"ee14a0c3d2a1145f", x"e2fce8b5352ced6a", x"8edadd9fcae2946d", x"fc9170b5ba6fff98", x"81691d2b6ad28ba8");
            when 33712908 => data <= (x"1966e19bac09236e", x"285196301e44b586", x"7d9891fef50108ce", x"69dee20a7ac2bf22", x"43bb25db717c2d3a", x"249a8d4b836bfaf1", x"d888e4fda714f56e", x"a22382999f969779");
            when 7955355 => data <= (x"c68fb087b09471bd", x"510edf78d59a6645", x"cbf9d78f6eb55f91", x"28324c0cdfa4f1c4", x"e2ee091da66511c8", x"067d716051f338b0", x"ec55f5e573d8a1a4", x"0f80c019453bb8e1");
            when 9677398 => data <= (x"f851f359be77d1c4", x"2fcf5564978ae3aa", x"cbb2ec769dd94bab", x"f5cae40686ad8e53", x"763ddb3e5d49b61a", x"8d7b77035861a0f4", x"2bc82dd05a0bbb6c", x"7d12e03996a6610d");
            when 6194746 => data <= (x"2b8e5f667bf0a671", x"ccea568c771440f0", x"ce25ebc8724e54f3", x"e8d8c6c65ff2e579", x"1ac06db4171b8357", x"3c5379538bc7b00c", x"d3372978c87243c9", x"08a34cfea1142186");
            when 23817849 => data <= (x"018546d13c399fd6", x"ad6262aa2a26c12d", x"9609944b542219e5", x"1b4df8d462e68b41", x"ffa6103d33e91403", x"3c12f02437943ecc", x"923a5e4220047be8", x"4776b116a55fce82");
            when 26975941 => data <= (x"76e17612ce2c18cb", x"39eb4c4b2e82a1d5", x"68885ca099a52df8", x"04187be10e5350f8", x"1d1381105cd5753c", x"d7ea6306ac54b25d", x"4919f888c8b197e9", x"e402a1752fb077bc");
            when 30374335 => data <= (x"aa5a77568b78e56b", x"48520e3f3452389f", x"405f6eabfab8ec0d", x"e217c7cf0120527b", x"264aaf4036b617cf", x"cb981f8ba8fda07a", x"006d140cc8b298b6", x"666ec952d4d8fbea");
            when 11247586 => data <= (x"d0a6f8d19f1209d2", x"9d7ed7aee022d5f9", x"9d9b76316508f75c", x"b36f5ddeebf1a4f1", x"72ecab5ed5b6e207", x"38302a7565ef2bca", x"a38da0d3b32dfeb5", x"4c3620db1220b865");
            when 10374471 => data <= (x"fdcca0b094941e1d", x"24a403a23328fee9", x"74b7206ec0132f16", x"9d034e999d87584c", x"e16c5bb14f8e6404", x"473c8f9e490bc0d0", x"e344e87b7e281ee4", x"71222f5607e6a028");
            when 27091578 => data <= (x"3007447ea5813544", x"72bb7b14dab419ef", x"b85ab95de7034113", x"b3159548465c9884", x"f0c4dbbc5cfeb8ef", x"ad21ff216415562e", x"027ac566033e2bf9", x"0ed4660881073737");
            when 32204999 => data <= (x"d6091be819986028", x"72d50191d5144e7b", x"2ffb9f88d048f951", x"e23e607f66ec3c01", x"e03695628e8250a8", x"a933cc7e48f5e3db", x"264fd8b6aac5e2b2", x"a9abf9b1c1a2f825");
            when 21533016 => data <= (x"d0da246a645a9d57", x"d8d824bb9e0e772a", x"f580c7cb62a68080", x"cb8afc00fb8bda5a", x"df4855e415973941", x"55ac4594d52c5ff0", x"594f555b934fb22c", x"dad9ae23c1a240c2");
            when 3299145 => data <= (x"aa6e1648433702f6", x"f84aa115ca609345", x"aeb932d1f5464e18", x"44c6701d22b8b1ee", x"7f8db54030a5a2e4", x"d772ad7be37f53c6", x"f0d80af7f5043d83", x"297a83e273f949f4");
            when 22128049 => data <= (x"15ef2588258a9f9f", x"006d60475af3420b", x"c46130ae768f6ade", x"48c2d0ec98a17d72", x"d6b3366c3b2fb613", x"3627607d8c05241d", x"a6f7ad5195c398e1", x"ae7651ddaf1addb9");
            when 25743003 => data <= (x"674bfd611d9d51e5", x"b39f5fe35786e105", x"b3f0c364ef6b79e4", x"a66ce63b17ba49dd", x"7792b8f5c3334bd0", x"f93061ac2df192de", x"347a7bc5d560a0c4", x"984e402e5cc618d0");
            when 26214737 => data <= (x"0ca0e9a488d7a419", x"b8d4185794692328", x"ec4663c0c3c1ff87", x"5b99bdfac8e7a631", x"c297b7fd48537ab8", x"72ee979ed4062da5", x"8acf5585a2769dbe", x"a47be0bb70bafdde");
            when 31672632 => data <= (x"23b1feafced7ac39", x"80fd436cb944cad9", x"78e20d86bee522e6", x"05f3bec7df40b786", x"1288c1d70dcba445", x"fe1396a8ce73c219", x"2eb29a12416350f1", x"1585f784cb558598");
            when 9907879 => data <= (x"f689cdbebc4ffd81", x"66af69a4e77536e9", x"a217cb2bf159861b", x"c9e39d1b1c039298", x"c6c2a49301b1141a", x"20901087a6ce2d02", x"e6e254c5864ab6ec", x"a717ab6e3056f38c");
            when 27352607 => data <= (x"c28719ea27a3e9af", x"e8e5ea40cce8c021", x"d109b70e2f5c279a", x"fc95a713e49ce1f8", x"734f36e9ef1a2d93", x"e7046f17df7dce31", x"ad2b1c6ee0df8674", x"c1c448b33a4a51d4");
            when 20484676 => data <= (x"66f2790983f46fde", x"5d73c2d2b0812ce2", x"e452c8dd26ff748c", x"ab69b353fc9fb979", x"97facd0c1a241107", x"a2a78a16f52f676d", x"95e0d927ef35d564", x"141824a1cee15c59");
            when 17869079 => data <= (x"3f28b9c4ecb2d65e", x"0f64ad769b49c84b", x"bea38184b52c85c8", x"ebc1ddca5c66d2dd", x"5abf52295be2c744", x"ee9929ba219a5482", x"63095ef05d945a21", x"5422730ec80c98a7");
            when 1440495 => data <= (x"7c42a5b1ae4d35e8", x"36dff7c0210b98bc", x"d431000e8e9a19d8", x"ce2421b1b7c165b7", x"24c2c24ee60cb18c", x"91e35a7f15554f28", x"2a25037d0ee81180", x"ad590d98ee3a0b5a");
            when 12086755 => data <= (x"7a894c73ed0f5e31", x"44d8ecf07fbb3efd", x"f866d7887fa585c9", x"8387e28203cc036b", x"3d0965e0ad512ff9", x"060ba10e31058669", x"446e0ac217813a5b", x"20a7008cbc94778a");
            when 12572584 => data <= (x"d42c7fc9d795403f", x"43a1f9ac5e290a68", x"2086d094dd323c87", x"15113354c7ae3c12", x"3a1b45aef50f479d", x"3bc33a129f9fb883", x"83b18879f95c1040", x"b8cbbaf443bcfeb4");
            when 31141582 => data <= (x"8e6ef7b32e642e94", x"2f2d1d23a5bb555d", x"399e708336d7b160", x"57f987eac5f3eae4", x"2e3be986b31c95d6", x"06ed876bbf969717", x"283c50b1f8b8fac7", x"9441af1cc74ccdbf");
            when 28817505 => data <= (x"98fb79fd45fa2567", x"c3bcb451e8926ba3", x"45f80c0248442ecd", x"5e42b52f1ff01a5e", x"085b8b9baac5f479", x"651fb611e4e09d26", x"b58920acf8045851", x"00696cfc4d25f59f");
            when 24114448 => data <= (x"7f0d70e48e5b601c", x"c366bd15f2501194", x"cbb7110465ef6843", x"f3f6f96d426e1085", x"50e85bd2b444b62d", x"c47e8dfbc29d3425", x"32e7dadb0aa045ce", x"30fbeb1f4da262bf");
            when 20598772 => data <= (x"d1e0f809ca982310", x"1aac4fa87e1796cd", x"e64b248eb95456e9", x"46291f02f92b7ca4", x"2e7dbae12398f1f2", x"41e7d4ef3638ad9e", x"9e386ddefe378b61", x"5e82a5d9a97ad565");
            when 11618987 => data <= (x"854727fcc1836e8c", x"1ed11f2a307bf72f", x"76a164d7e08804d0", x"10ce0dacf7f4b6eb", x"406839c78860c1e4", x"54716fc883c58b02", x"0b63b94fd2e9d70a", x"b78fadd5a2ab138d");
            when 16744593 => data <= (x"13a1723cbcaaefbe", x"d13df884e5eaa5a9", x"c547121dca631acd", x"61aefc726d997640", x"3831d1b4b477ae92", x"676e72666e09faa2", x"18228727ff08be37", x"3f7c2ae58a49676e");
            when 15954736 => data <= (x"9531c30d968940f1", x"7a26936f6476807f", x"5d8eb1945d13607c", x"2ed3832abb664240", x"f67100123e6d1d0e", x"49bfa4b7a56cd3d4", x"a9aa0084dd2b5856", x"c56062a608c96ab3");
            when 7587429 => data <= (x"a85fa9ea33377dea", x"9f0df1f5fb7b21c7", x"e55ee1c8c993d76b", x"e64575ca72856cb8", x"ef118a44a90ed4b8", x"046e693dcd68ba96", x"ae559f8642781eca", x"00f32e926119828b");
            when 2807920 => data <= (x"658467965b25a78a", x"54fe889ca5cc328f", x"55d74b7cd7181fa6", x"7979e293a1c8c9d3", x"b55644f899b62556", x"6349e71a820ad268", x"bdee6a26e227afcf", x"dfea564e4860f46b");
            when 5745743 => data <= (x"51a727441e776beb", x"348368f69336ebc1", x"cabde3d0c75b4e60", x"ee62061bad68ed87", x"8443449af260dfae", x"5279b7a92ecc7340", x"331ad38b64c1a989", x"1243dcb5b957509b");
            when 27890874 => data <= (x"7d6d3c51544c89d7", x"25242495fe4c62e6", x"d8af46088682e958", x"f9f7e3590435e5bf", x"a9854b52747257df", x"1f720b557cd70e3d", x"0b97017693f5405a", x"62cd44f64574811b");
            when 17307805 => data <= (x"80d76ab6974b4cf1", x"d541ef531575fea1", x"9d519788276b0940", x"67aec5461710e05e", x"961e910cd78b6dfa", x"cc34f1597f043f6e", x"c66c26fa6f14d877", x"d82fe81a9547b95a");
            when 8397946 => data <= (x"df90c3664a937c8d", x"1e20cc397cd23050", x"f16875d6c7b17300", x"558130d8303463cd", x"454eb4dc909eb38c", x"d0c0b4d3f04f0d99", x"6430553e54f1dd9c", x"e066f42454ff9b1d");
            when 23363775 => data <= (x"26051c3dc79aea68", x"42657ec58c212e6b", x"0beed44cf47b8bae", x"81d2b5ee6e0f4ed9", x"1c344caa6ed861ea", x"66e0d88045a634c2", x"400a6f5b397b459a", x"144c11442090a0de");
            when 20868006 => data <= (x"3915beb8bc671d0a", x"69be14d90eec4162", x"80157ba428eed1dd", x"469b4e045e94ce98", x"e56be7bc13ea7b83", x"d74304feb0ab1492", x"e1e1b37fbc66efa4", x"8527c8648c981cf2");
            when 7054877 => data <= (x"983523026585f046", x"4e89da1269792041", x"0e96bfa219061942", x"ceee2e387c1e67a1", x"f55a2829f17cec12", x"58751482a4cc49cf", x"81bc838d886a744a", x"08c949d5be7deba4");
            when 16743547 => data <= (x"8cb00c8fe8782a43", x"d9d08b9f64332020", x"47a6c9b58db95724", x"598f9778b361faa2", x"c4fdce11962a7475", x"46eccea6330d992f", x"bfed5e619570088d", x"4b516c36769d3b63");
            when 3626931 => data <= (x"35335dbfbc9a7215", x"fa9cd48423a3b834", x"c1fde0d28656a3fb", x"2cb54e26e74adfb1", x"ca08b69dcbf0eb0b", x"e0e735d68f7ba4f2", x"ad47bd2c18276b64", x"bfff142959956aac");
            when 11997647 => data <= (x"e7241ed2aeb516be", x"7d2d852c6c68eee1", x"17b13cb87de6cdd0", x"d0415921e677d550", x"842d419a3c587542", x"589f73412f491743", x"3c36f6effdff5166", x"075d7e30239fdc81");
            when 1993515 => data <= (x"14b286ed3cc4821c", x"695dcb0869e67b2d", x"bf30b037f0390cce", x"40f2ee33869acaf9", x"49e58b6f33b08827", x"f94040abac029c12", x"fd890adc172e9ebd", x"b0646d5314edd7d6");
            when 27664811 => data <= (x"7395e24c57a8bc66", x"10fdf3bce15ea6bd", x"aea7ac73eab46b6e", x"2a1ef838d9f032a6", x"defb0c8002e5a3b0", x"03a98ae23d8704fc", x"ada60207f93f850a", x"87a0d11d0931885d");
            when 1473323 => data <= (x"84d5468a9c8edd39", x"0d02f68f6ab60e7a", x"de486ba38c11196a", x"1c7109553e56c050", x"e7d6ddccebbe2729", x"fd599cbd1edfa95e", x"8000358fce114ace", x"4b02008c37d9a51b");
            when 15441950 => data <= (x"b40fb4dd3699d730", x"e1fd1a9a7518bc12", x"86df4d18ef97df1a", x"b63446fce52a79fa", x"5d34779d499e0f26", x"80ad94eb154937c5", x"19a310c1f21c3325", x"7db28bc382c824d9");
            when 33741835 => data <= (x"fab7650aad819508", x"859c51d8d58ece63", x"4e15abb8dfe70a73", x"9c49976f51dc6ed2", x"99763ff33e73b068", x"b50ccd7fa1c11fa8", x"0e3a57e3f1d1db1d", x"2a0eb55c8b090f1f");
            when 21936879 => data <= (x"478383bc0d2babb5", x"b54d46d4a052eb61", x"df5953a0c7c1deff", x"46dabb78b06269d3", x"a728c34e7da9431d", x"c7c923df5d43fb1b", x"c2da083060aa8c69", x"33786c771c2ac6b8");
            when 29177065 => data <= (x"aaccbc4c8b4bbb9e", x"b44edfe4d4c67acb", x"1b2a49ad23ef989d", x"80a9ef8696f03a45", x"1c24c35842ea634c", x"e64c2bf9a1d2ae70", x"bde3cb46fdf8116a", x"7f30d2d27121fc1f");
            when 9888997 => data <= (x"09f0235967499861", x"0a4ce016031eaa91", x"db06a3767493dd1a", x"33bafdd91706fa6f", x"2399fc46502e9526", x"a441e50ea23b1f22", x"6d731b608a2cfbf3", x"68d0fc89ace66601");
            when 10181344 => data <= (x"df2bea3b98ffb4c1", x"cf9774297f19b133", x"fa6b6a88852278f6", x"b1cdc22a7e0cfa8c", x"b30886d5f0aac5d8", x"4f1cebbec3914038", x"9da6c7f5651dbd23", x"960634af3af6c071");
            when 3345085 => data <= (x"6982e8f3dfbd454a", x"16c355739409d22c", x"263ee8a49d073932", x"26e93b0a190172e4", x"b6cd3900bf7a6c5f", x"1fb88936deb8fd8b", x"188a287c818079a8", x"76b86ee468d68b5d");
            when 17316512 => data <= (x"890888891c7f2ec5", x"2765850fc4e39809", x"ae3110fdbfc9a46f", x"2f2e49a8adc633ce", x"8345cf61a8cb216c", x"73ab17bcfb8dacb9", x"e5b82cb1cbe5a919", x"34daff1e71596196");
            when 11354797 => data <= (x"b48c6702a72a24db", x"03542256df456706", x"94355117a0bd098a", x"ceedaaad6399a27d", x"657ad1d1684f77ae", x"b22755063e673fa3", x"3ee00d60797e7bf0", x"b81af109598fbc0b");
            when 6063738 => data <= (x"a3c0e87aaa0416e4", x"42dc30b9e213c7f2", x"1a4be94a8d6dff7c", x"28c6906774f93109", x"fe45dafa09f8aecb", x"c9992a7d40166f04", x"fc87c8ffff5d3402", x"6dea07c212898767");
            when 16604465 => data <= (x"a587bd80bdb2d736", x"2f881d668a7c5eb9", x"6eb9168155bd0642", x"1e926ed7bafa2f24", x"0b7c48bcd9c78b38", x"460baa0444a523e5", x"e9bd651e20619dfa", x"418881e5d4a04d9c");
            when 6831659 => data <= (x"3341a132359823cf", x"eccd7f97cddb6bfb", x"404edd1feabc9c06", x"dce30c5dae122e34", x"dd648cb9829dfd3c", x"df4a27d3a26ab910", x"873f8fba6c0ef613", x"d65a659596ba9904");
            when 16178096 => data <= (x"0ceea80d03b02f61", x"a116d8a9ffe67dbf", x"d005b872260db93b", x"4c801792b8672606", x"e4002314bba89d94", x"597b84c5a9e8543c", x"3ca9df824b7d4e9a", x"0d878526029b5095");
            when 21387587 => data <= (x"7c12d40af1dc933a", x"45e605bd19023835", x"7d89a5405c9c1806", x"2f0b39c76f5b4782", x"d0f889b4a3a45691", x"38fda105e61e592e", x"31db82ddc180a65b", x"0ba151389658d156");
            when 26384581 => data <= (x"4852ae1a19f40692", x"3f7ee2ac1fcf5f52", x"68fc3accffdfe8b4", x"692dc575f329fe3f", x"4ba7a33cf18f5f30", x"e47a4ba5969eb1e9", x"9a2d9956d333a0db", x"3b33fd218721a343");
            when 12705148 => data <= (x"aa607a13a63aef6d", x"9bef8872ad831d4c", x"34acb3b356105456", x"2aafe33e7be78b28", x"69bde57d6c4f1526", x"0421b45cd1072d4f", x"79ab2847412783b0", x"5718239f159c4587");
            when 21863307 => data <= (x"63049326fa58eeb3", x"7e5e97acb26618f7", x"9ff736384719a5a8", x"0813fda69959ff22", x"c2bdbb58ee49ce1e", x"47804607b699758a", x"81c78316b843a57d", x"007e4a6635ddd6a3");
            when 2946148 => data <= (x"600650bc5c7ffcf8", x"8aca015c4cd16c06", x"89b50394dea37982", x"4d0b76581d9d5a54", x"60b0efb5058271f5", x"011e03876f3fbda0", x"bea2d397b899da95", x"60bfb346e0685440");
            when 30380768 => data <= (x"9b5829d3de8bc2da", x"84d76e330f8d2109", x"9150bbf6891f7bef", x"c2637e7e4adcf2a9", x"b9c851d182b9d7d6", x"68d0ab4c7c5d7a19", x"608a579784e76ed3", x"73245698cd7a1e4d");
            when 26864814 => data <= (x"0863b8c322a0be01", x"5d8a1f541dcd5904", x"d7933ffcdfdf2db8", x"35e4827941c964cf", x"e78365ee9e36243a", x"ffa82dc7564ff7cf", x"1c1edc1ea65a2246", x"0a16cca95b5a3b45");
            when 29395918 => data <= (x"eef6797b9df62ec6", x"d891f56f0e3fa598", x"cca589ef89b93dcf", x"af11a61067f01948", x"c7b97d1cf5cf2685", x"752a7f3ed0842f91", x"82368ea96fb30770", x"3eb9bbaa833abdb9");
            when 21903424 => data <= (x"67db8c2491c02572", x"9afd47b8ec3ff01e", x"9e048e9247d66631", x"f3a195a547c74307", x"1919e05736f0e95f", x"5de4cbb3d3721bf9", x"1dd2416d854da33e", x"75314f3480002d65");
            when 10957121 => data <= (x"54a4b70da9d966b3", x"902a8fee7602eb1c", x"d2bafc6fac7b0b47", x"1ea5396e9b8698fd", x"980b6b407bb69881", x"15c4860f1c21acc0", x"50e4c549ad84cde9", x"2ef06097f7d09b3c");
            when 27513183 => data <= (x"0a3a8ae0932a9754", x"1879d38499372b3c", x"9063f907a213827a", x"51f3b8bf63c05549", x"a57eab4a3915c5e8", x"d502946141b5f4da", x"a7bad11027b96b32", x"714799342951c18a");
            when 9930554 => data <= (x"d0c7114f548658bd", x"2aeb9e9eea347f54", x"fc6802eca8ee8d3d", x"9083c7716c4406ba", x"1e802d51cccde469", x"049e2098473837c5", x"422a3a0538771e6b", x"5b40d53d87d17a21");
            when 27458357 => data <= (x"8cc9485bf7c5efdf", x"a438979fe30b0495", x"4552500a2a077753", x"d47528c84aaa7f10", x"6a830fa4d1df83a9", x"80bcc96670cca44b", x"7a4dbfaa134e588c", x"34abc74471c42266");
            when 18536891 => data <= (x"25a65542c24ba75d", x"2b26c2705827311f", x"194b3fbbef195703", x"fee92ef0df6cc206", x"56777621813810bd", x"f5814c20e903ed5e", x"cdebcada52a9a9c2", x"4eacab144276206e");
            when 31253171 => data <= (x"97dc6e817f544ac4", x"fd21882b3a3e90df", x"0daa275f23415092", x"d9fbb73df46fda33", x"27d2d327f027915c", x"1b4d5a5041751782", x"f9dce7009edbdde5", x"f20c21fc11d56c1a");
            when 10161710 => data <= (x"90c7efca04f91b81", x"5e0df04653738f2b", x"dc3197bc4c7589f4", x"f805650ef7579e43", x"f9059cfd5c91888e", x"2e85fc549d5a6b83", x"137705114cd99a39", x"87f0db5f9eca077a");
            when 24868766 => data <= (x"55758cbada1dedfe", x"ce43b6a2b9af5cf9", x"58f21766464df51c", x"22fc4515e900aa50", x"ac4e240e90e96b79", x"b1eed0b2dd9e1d51", x"81ce13a0256df174", x"6bb75c01e1c4f257");
            when 22137760 => data <= (x"ab099fcff1a63892", x"da435cdf2fefaadd", x"7d86ffe199b888f0", x"6b5e1739799c1c21", x"647742b9bc1c6f1f", x"8d3ce6c49496dcc6", x"dd57b393a49df273", x"e53e5122134a26f5");
            when 27530226 => data <= (x"c560f1bcec5772fd", x"e78ca610b48c65cc", x"f94f9034a628318c", x"a3b79caa8782ba8d", x"7f5e39b4b53a88e8", x"5349fc3dcc38976e", x"6c643698939f3139", x"240e6d1fa1ac9b7a");
            when 17395593 => data <= (x"be3df4b3f08ba487", x"0d28e49c284477b8", x"097a1dee984085cc", x"ef388f732593e1c8", x"965268315c05e5fb", x"7a35de45ae354576", x"973a6d8705d5f3ec", x"9d9466b280438359");
            when 22766805 => data <= (x"ec51e917c8568955", x"d742e330d9d6b06a", x"47a2c5b3c30f5608", x"91a21a8bc6347f5d", x"8606405daeb1482e", x"e88db838fdb15a52", x"30d5aae2936be4de", x"b98206244e95a107");
            when 32170849 => data <= (x"237fee7670dbf13a", x"7ab6fa8394e49f10", x"6fc59bfec612d4b9", x"1728e83c3268925a", x"02250601c8e2c832", x"cac87be0fe64af8c", x"88a9b65ec660e93d", x"510487faac6fce4e");
            when 7393635 => data <= (x"49abcc1f67ef804a", x"734686715db97f62", x"e47799ff7e9dea36", x"8544d90e3158dcb2", x"10e3e218daa5d6e1", x"c941bd59746394e3", x"fddc1096157e7d12", x"3f8ef975718dc52a");
            when 11510413 => data <= (x"472c90af6fa218ac", x"b5b8e1ff725a027f", x"fb2e0143332c94bd", x"dfbd8be45a1e7cb4", x"c27d74d87e632187", x"36cc65c791ce2916", x"60497312d7ab6c02", x"bf446653d45b0a28");
            when 22590355 => data <= (x"521caceb334dbb0a", x"fe4e7d62655d1243", x"77b57b608633949b", x"5b87be99caa54a4d", x"5c9e4bfd5966422e", x"4b9e1b4c8a644f67", x"0bf5438ecf43b7db", x"b05bd4ffebf913ce");
            when 9165464 => data <= (x"2ddedb4e52eeb70a", x"f1a6ed37b0020fa2", x"ff84f817e781dbdf", x"926d9bd0c9fa6408", x"7a97432c6ef12bcc", x"e26f974c9993beca", x"e5b9d377f9599451", x"48c0387c75502232");
            when 3047957 => data <= (x"055531be81a5efdc", x"e92a41682819f647", x"75a96a57a6de2940", x"afc8416552eccf82", x"8c61638aeba087b8", x"3d2918f00e195f85", x"736fd29b935c8438", x"f8b2ee713f48ff04");
            when 5412056 => data <= (x"8c2aec4cba188342", x"30a8ef42c5a90e4d", x"3840ca1950bbbaa5", x"8ab5842f8fce0e96", x"00236a261f79d03a", x"adc640e9650cab83", x"e9f9519ca6ba8c71", x"f36e761a2ad65cdc");
            when 20061593 => data <= (x"0243575dead3203c", x"8bd1185b01023d31", x"e98d7adeb8b3783c", x"5bd792ba00b1dd04", x"3efb1805ec359748", x"958697b3c56d0497", x"ef054427cf6f5710", x"877aedd2dbb38e71");
            when 28602097 => data <= (x"036e7afebf39d44e", x"12a68e6173c94dd3", x"73be6b314c2a967e", x"796cf0c299c39971", x"bb458ff8f19d6205", x"128e2eb0c964b262", x"bcf5d579ea724fcd", x"57a28132253a1a4c");
            when 6446460 => data <= (x"5fc1a491a39d19df", x"363d4f934a3ee203", x"9c41c7dd424f5bba", x"9c20cbd28a3cc091", x"966bae13e8adcf98", x"fff54dc5fd06bdfc", x"223ebcb9477cde8a", x"463509b6336e1c5e");
            when 11377824 => data <= (x"3098c8236fd5b8a8", x"838031a76c6c7ccb", x"8182b3b0d964dff0", x"756035d0c9db3573", x"3dfe94849670c2db", x"340b37a555ae943d", x"665cee20acca32ec", x"bed96aeb1e50b2e5");
            when 18416625 => data <= (x"baba4fa0b2880550", x"1d58c2213829f66d", x"07a00c7a8cdd30a2", x"a271bdc672e67838", x"b26732b12272e8ab", x"55ece30eb484490f", x"ee1de65d321961ba", x"ac901093004c03c3");
            when 11005654 => data <= (x"6e82f1f66088cd06", x"36ae6c91c22076b2", x"0e58b2ea9bb4087e", x"2182ecaa843dc667", x"31706616f596ea56", x"2773eab4f63c5232", x"691e274388ba84f6", x"5c22fc892cec7e12");
            when 28275175 => data <= (x"0ee63c0ac8c5156d", x"c134fb49ddb3767b", x"436f095faef7ef94", x"771732e60ff3e0c8", x"18e58656758190f9", x"6402e88eb7550df4", x"8ea1224809674083", x"23c9fb9922e52aff");
            when 3365203 => data <= (x"ad600d2275f0d1fa", x"5b6a920b7f017e59", x"d83dd53f2b4610dc", x"9b41b9220240e2bb", x"a93eb68a961030e9", x"35c7e3b969415a1b", x"f9f5bfe0c7ffa34b", x"7c6b7a3d7babbfd8");
            when 19591765 => data <= (x"b7bd106186527e71", x"e5096ae91ba6a644", x"b1c691983f860050", x"cdd403e36c1a6e5f", x"08aad40af697371b", x"8ec70eaf00bcc45b", x"18d24a20dcd9ae56", x"998cc55dc9d3ff73");
            when 30939560 => data <= (x"b999766fa64badc7", x"3ca8ade468108a8d", x"bc60408276b9974a", x"483ef6497b9d04ee", x"4e905b28118e4606", x"812ddb1954b9bee0", x"5934b83f221940df", x"f27a057c01b646d2");
            when 14471194 => data <= (x"0af5f6ad9ac04af5", x"8c4a784a6e8794e6", x"f30f793aa8624273", x"02ac7b69c90dacab", x"e32af60ec990c26a", x"b3ac94d1097ebd9f", x"76e8751f3c9ed1b1", x"a4d10ee1ca278898");
            when 31614448 => data <= (x"e12a80c4c0cbdab4", x"35fd61604b010d2e", x"0b3c04a89afa8d77", x"6b89d374b3946c19", x"80e89d18fb6968d7", x"92a3a3afd44cd8e8", x"a41473e15c5adb74", x"4f1527674ad6463a");
            when 13724333 => data <= (x"80777f1ba187fcc2", x"ec6a58848f3f54b5", x"a771e3cdd277377a", x"d3083c5879578064", x"92f32727c7cf36e2", x"c6f025582cdab540", x"62e937ab7d64e3ef", x"8d6a8bffe68eb09c");
            when 5111335 => data <= (x"d5a206ad049e6064", x"c0a272b0bbd2c75e", x"8ea150c2e0e56bd6", x"22e7567d22fc6028", x"78ad33c9d7219743", x"ab9b3397b768ed0e", x"cc2562e08796807e", x"34697b6d142ffe1e");
            when 1418193 => data <= (x"eeb6ddab1477eaae", x"99cc8665408a043c", x"5d15abd5f8141416", x"386cdfd498b5734c", x"94a1337c7b41ecce", x"371596a67fdf1f22", x"cfda16941a837721", x"27f908b1ff6edd2f");
            when 26404778 => data <= (x"aed42881c36cc255", x"f2f4a1e04ce76738", x"4546a4494cc80f02", x"d16e7a719a74f464", x"abf2d86d4c81b3fd", x"e63f6ff0b3012628", x"6cb4f26666bacef3", x"d09bc673a7b2803d");
            when 4701117 => data <= (x"6a975671ea985529", x"302fcf11873ba68a", x"84d3f8298738bda1", x"8c5667689da25b5c", x"bbb4a8693498c7c1", x"c18a3e1d5c2f2a57", x"72d50efcc3b3f381", x"daf05322384de1cb");
            when 11156316 => data <= (x"bb8e9710f5bb56d0", x"717534c666c0d361", x"a8d655ef1af3baff", x"469f416291151122", x"ac5d3b9d93246029", x"aae350476de81098", x"e3059eed2e608589", x"362e1b7a22823042");
            when 24629344 => data <= (x"cbfe9f6c920ac00d", x"7a566653359519c0", x"4edc5cc23eb45ca2", x"0c80bae97779dbec", x"b9e33ac9a9bd079e", x"b86230cd4c38f178", x"c6c58e4ef340b17e", x"2abaeeea6750efc5");
            when 25666709 => data <= (x"c130f38843fe2929", x"410990481750075f", x"645b846419e316ce", x"694f8a994f3987e9", x"2f3cf291296effde", x"0f8e2f765a5a648c", x"ff6215fbd13093c6", x"00bcc586d531aad7");
            when 22276747 => data <= (x"274c8525d3c6d381", x"4193af90264b7144", x"3795c7bce2a45f31", x"073762b10b289f9e", x"feab38c4b00c2232", x"9130ecd8b8c61ac0", x"d96a992d0e70f11f", x"1c98ee5e7e70482c");
            when 17071588 => data <= (x"da35750af2b24764", x"0f01bb1670058e9e", x"a05034cd532cc788", x"0fcd6b6e6f144e10", x"880a562f359d20d0", x"39c060f410e1f9d9", x"f60f75984c644fda", x"fc1e3579fb319fd6");
            when 30563278 => data <= (x"ecd92ef09c2d9693", x"4acd55cc81e61016", x"0048cd1ce1baddb1", x"038284932a345b5c", x"b48ed10506075dc7", x"7e8958f6975361a7", x"6b478ac5cf7326ba", x"ea448a0b9fdd1133");
            when 24330975 => data <= (x"12e9d2822aa77c55", x"c8858ee5db93b719", x"b1d1f041817b5a76", x"49f3f5cbf931e066", x"2633a5e46d92b95d", x"d1ed727852cb470e", x"8b3c75922fdcedb5", x"5d1fa66611b555ef");
            when 26687326 => data <= (x"aec3c2e85e1e2518", x"f8bd0a8a769b68f9", x"b1e468ea8db238ae", x"5d02ce03d5ad22d8", x"938281f731aea97f", x"e27155bb127bba5c", x"c6bb43a1421bbc88", x"0fdc7ecf32ae7f61");
            when 20392719 => data <= (x"12054941645e5198", x"5e9a71931944dc67", x"31c83abc361600dd", x"1c32032d4148d10d", x"39ef30787107b227", x"bf51cfcb6028acdc", x"b3f97a0373b9b1fa", x"35dc223b744dc42e");
            when 26093428 => data <= (x"1dcdc906d313f6bf", x"63cf0a6dbc14911b", x"4f9b4c7b6c6e8e94", x"624f57318f9caab8", x"636ba4592cf717aa", x"5edf36e7daf3cb07", x"9db423f6be584b95", x"93880f0d94afac2f");
            when 15645116 => data <= (x"6421ed3ca8774050", x"734e6c77e8103748", x"c7f308dab1147404", x"d762fd155e9979f7", x"fdba06c187506da7", x"75ff70fed0c0e859", x"97b4788d8de77ff2", x"6717bafcffcb19ce");
            when 19375628 => data <= (x"180efa1933ab77be", x"469fbae2b710787d", x"9cf10835b0fd6963", x"6ca35b8cce4ed879", x"8cbb0cf25ecf5e2c", x"cd900fe634fd1d76", x"18aa1500c7f84f41", x"4a7b9dbf6f7cbda8");
            when 31508437 => data <= (x"788783cb7447c9a1", x"2ad81d07f2e3c680", x"f9919e692d7fa5e9", x"c806ad7b910054bd", x"9235cae08f5f2958", x"5a1a3add29b8f07f", x"6c2bcc31da12e03e", x"abb184a2e96550ec");
            when 31408029 => data <= (x"5cdf7994276bc07f", x"91044fef25f107f8", x"48a94f938ad26e69", x"cbb2d2815d095f87", x"0988c64aaf2f1bc1", x"348f27d50abe3f34", x"4c1157363ed997ca", x"78e0e9bfbd9a9952");
            when 23771047 => data <= (x"dde2e3d74d9cc8bb", x"84772b4174ed0186", x"93eb03ceda6a9154", x"a278f5b59b239710", x"6cb38b6941b38fbf", x"a82eafa6de4cd329", x"2678ba23ac4347fd", x"8a047efa6e905026");
            when 28757522 => data <= (x"1efdefb0df469c27", x"aefd042a60e84e0c", x"e3e4922c129a3284", x"41c1824d7e236498", x"1df5cc90a40baf16", x"ddf2d94a690b1205", x"ac8db6b2ce23a4de", x"16a7d39b2d024e61");
            when 11833152 => data <= (x"7c56fa173d8743a5", x"5a85127392774b0e", x"7bd19ec372c1c1e8", x"6d25ecf51e4837f0", x"1e47e97d717fbc86", x"6c20b9882dd26c73", x"84ccd39cec27ec03", x"1e6a6f0b7d2081e5");
            when 427570 => data <= (x"ac850e1aab11ab98", x"b7fd54b0f4b8fb65", x"82db793183ecf9fc", x"ae0f073d2136a371", x"d5636bbcd8d10646", x"329f953bde01f305", x"97c479c266c6f65a", x"b2ecfb6601ac46f9");
            when 2915726 => data <= (x"2385be654f9af18f", x"6d258fa76674c7e6", x"f6af34fbdf4a0ee5", x"9ce7f58c0489731c", x"15b214d86cce8874", x"73940fae2e9b3147", x"48f72c7fe0daf976", x"153229d8a03815cc");
            when 15587662 => data <= (x"d6968c6b5754c20c", x"ce93d833c119da56", x"bfdcf1c8cbba7001", x"a91d32f7ce6b0371", x"374b1c1d0199c817", x"58ad450f88662131", x"3703d7bb04e1de59", x"450d7787b3a13d75");
            when 11041976 => data <= (x"2fe653902ad709a6", x"c24f3d2945c5886c", x"00c67dfc0ee2fe38", x"b6f570e3cf8b5cfe", x"cdd5d71224225927", x"b800766c03e552a1", x"be090ee8c2755084", x"b462e95395270b3d");
            when 16955774 => data <= (x"aa501ca5b7f50878", x"70652c01a5053558", x"a323c61221a8a02a", x"a2e73442b54fd611", x"da4d07480872ead1", x"0b04abf286f4ee0e", x"dd49795e24698ab6", x"e8e7f1dc5a4af8c9");
            when 5681836 => data <= (x"37896f925cd91b54", x"2d33dd0f2373a4cc", x"e59ab94b565a7ec7", x"1c0f7e8212505c0b", x"f54a89dbbd650a42", x"904fe4b98139bc42", x"340c8aae11da44db", x"1a60f28d725bd0f3");
            when 20709423 => data <= (x"b208932c671be085", x"68b0e7e1a0d4a339", x"ef1b322b7556c032", x"ae67a64a44ff3d0a", x"79245c9fd0d4bd78", x"de527615d78ba2cf", x"aa0abe6806111cd5", x"33a18a8ce83585ab");
            when 27916739 => data <= (x"3e6845d34f56397d", x"36812f0b8615be94", x"8ad319c9d99ff49d", x"ba6cb196a8de2809", x"97a5b6f7722ea32b", x"d515121fc2215402", x"598422d831df83c3", x"366b10b329579040");
            when 5370513 => data <= (x"605d4f699d85f752", x"02464d7201b176dd", x"7e8fcdc863153c97", x"df9ed85597099f4a", x"a433888eed01bb74", x"aa5dae73dac6e39b", x"d4dadcd9c12dbd5b", x"be91422e3e1e5fb2");
            when 24564100 => data <= (x"c3d6402535ded23b", x"044207d5427e3ee9", x"7591a734675e470e", x"5949eaa1784389c6", x"291cf39b3dd25f68", x"a5429bcea3cca9bc", x"1546ecd1b2d56297", x"1161a5b6c6403b77");
            when 22516355 => data <= (x"35ac560cd1b662dd", x"b509e798af7f18b9", x"c3c618fd430791fb", x"bce500a9479dc835", x"2cddb56599c45600", x"edf4c5ef06f9cbeb", x"a74e73bbe1a63624", x"229585c4d265426a");
            when 27917235 => data <= (x"c9f4f9907fb68486", x"d4ce8f5c2c8d1b15", x"9690f2ec8321b4db", x"d40d1d94045dd01f", x"f4218994cb67e439", x"e5fb064f4c4f84d4", x"f8b2937d02621ecb", x"7e656ecb7da87636");
            when 29664768 => data <= (x"0fff41024a72ba14", x"e0e041629d729399", x"2c533df748a53691", x"74dc6f7e90b71c44", x"fe21b13b2c7fe667", x"cefa6446e64a7c15", x"43345dd0468c52d6", x"af550a8320988bbb");
            when 20388759 => data <= (x"3cc0090383c2921e", x"138fbb25ec1a2d2e", x"9788dcb0ec20baae", x"cf4a3f7fe2d8c041", x"08bd8c9be79a3bab", x"c79717dc25e8e93d", x"16635a20e628b71c", x"b7ac67af88bb4d24");
            when 23835637 => data <= (x"872194753508c3f8", x"8a6c709238102bea", x"1bf1772b649edcf2", x"8919351376053200", x"55023b74b4bf2c87", x"1d2ebddf80d849c6", x"b24e43b18a3f21b9", x"93871af2a33ab01d");
            when 15431548 => data <= (x"1d545511f68fd291", x"399798511951d578", x"f923ba08164784b9", x"9c09924df2d43607", x"735f6b1ebadafa74", x"38a6c1414d5aaaf3", x"38fbcd9a31937085", x"66ef65efd3928625");
            when 7400390 => data <= (x"529b6a53b48edbfc", x"11f8763fa79d6a4c", x"8d68b5861f90e2e5", x"56928e69349e4c2c", x"c8c8a3cc59f73c23", x"513f58997872110d", x"25e58e86571fea57", x"0f62699fcf47fa87");
            when 7414855 => data <= (x"6141842daf81c3fc", x"d710d26b24fae199", x"37cfe25a49d46d82", x"d86d31fd5cb3767b", x"5c226cff09f9ca0c", x"5c58e6c6ffd16093", x"c3b09a8439b9556c", x"55eace355544a99b");
            when 11146285 => data <= (x"7bd80f3b3df5d58c", x"3eae1d1bc14df029", x"2ef8538ec33cb65f", x"a8e544c78b1eba06", x"76b39d173a0eb8e9", x"34f91d702f12d90e", x"d784440eb4f28624", x"620ab2bf1ff0aec4");
            when 33047682 => data <= (x"fc9d4819854a469c", x"c392b8c4749e25ce", x"ae6050e353a3cca8", x"e64ee12e7ac1d6e1", x"4c2eb44617e97b14", x"096f69cbf792b9b1", x"cbd65cd3d0bb0ab0", x"a35d9e03b4d86c12");
            when 3754329 => data <= (x"87d78304e4b828be", x"a6ff5eee7f40dc70", x"c67d6921fb07e443", x"f1e3f98c13659116", x"b976959f972e93a0", x"436e25ef2f2ea1e6", x"91f2c3de90c8419c", x"bc6373e7134a8741");
            when 6394972 => data <= (x"1095d5806880bff4", x"5923ebe7c072b32f", x"7ba90012bf1e9362", x"3391ef914afff382", x"a7f61c4d88fbd374", x"7b23b929f197d29c", x"f52f9f80b7d11baf", x"2e2fd210f7aedc47");
            when 27182173 => data <= (x"8d4ddac37eeed30a", x"2fce1fd9099d87aa", x"c1bb5443065de30f", x"8169ce3089fd38e7", x"8a6e91e35b4c7be3", x"da80e6455779d995", x"ee730997d3da3e8d", x"32a686528f36fe8b");
            when 18735087 => data <= (x"f1eeb917b8321840", x"3fae9a7668fd0cf7", x"31f177eb9c555230", x"dbe65724def6c16b", x"651ea8e6efa1e631", x"e3aff8ea8738cda5", x"625909ccfc0abf86", x"7aca11a8490ae9f1");
            when 22648434 => data <= (x"4c65fb99f4b3eb6c", x"118cb4956035fff5", x"fd4a5cef5c2f64a9", x"fd990469f9cd92d5", x"ccdbafea9fba37f6", x"91b7a4421c10ad76", x"d027dc1c5f627e24", x"0c7328ec8b8abcca");
            when 33311886 => data <= (x"37f4c6b116517ce1", x"fc4807d1832d4bb9", x"9bfffb14d1e08a3a", x"bdaef1726cd9ef9f", x"c94341b316219643", x"e15d15b7afe62bf5", x"a797d78f8ea301b2", x"e5d0a41f33920498");
            when 9812066 => data <= (x"73a5322541ed367e", x"678c1ce0c2bb1b63", x"e1135ee4bcc7185d", x"ebe8e1f063a2cda8", x"bf6b92d89f703c6f", x"866071b6e8b63768", x"d6d4e27bf2f443bd", x"848973c7e4aa8cdb");
            when 25014625 => data <= (x"a53b50c9985d2173", x"12fe8bf512f044cb", x"5e01583fc36b6d47", x"a644c73caba7beef", x"4927bff947f63340", x"f53cec0dc211c245", x"1ac8459c551ac1b3", x"89d3b80c8be28abf");
            when 12617438 => data <= (x"ffd97aca5a0eddcb", x"b7c9408108d2d5f1", x"b096ca192dbefe78", x"c38cd10c3f877cc8", x"530b83255913d07b", x"f176b5cd28ec63aa", x"d8420a292a104628", x"d532cb80e1b04dc0");
            when 20308066 => data <= (x"7a2859eec7f43027", x"7963f2ed85ea640a", x"8bd5df372559fd25", x"f1d97a3701806c70", x"99eedeb146f4e906", x"3c2188f07f19cd80", x"367e2f559eda813c", x"240ccbc5e94ee352");
            when 33629531 => data <= (x"10420a0130a4a353", x"d1f7f5269c3e1868", x"dd241d6455f06cf3", x"aaabc5928cdbfbf8", x"b37ba674591f0703", x"e7102c5ca0a2a175", x"d03357c6fd155dc2", x"f905a3ee67ccf884");
            when 5641211 => data <= (x"3efc2edc4e8d06d3", x"565cded81d0fbc06", x"c9b1bf0e695d4295", x"e6654113cc3b45d5", x"e2422b7ced6ec0b8", x"d009c91d2c289b9a", x"d2bb4260821d5c7a", x"0c9603b86011b3bc");
            when 16562884 => data <= (x"18662fc6232dc0fe", x"3b8f87a27d7cda89", x"8d573a36027e7299", x"c589d58619543241", x"3458b82858700051", x"147cabe02eae85af", x"6b5618b4d0909bd1", x"543462c74f18df92");
            when 4331596 => data <= (x"cd37a2fc322e4f3e", x"af1824a80dd6efb1", x"8d1b9db12f3a0340", x"9ed43f8b6aa241d2", x"dcb747ad30d87438", x"53267559eae901ee", x"cd79e873c6379401", x"3e25e32cd98cf88e");
            when 26550696 => data <= (x"632f94109dec5e5e", x"472075f3c0fb83c6", x"2b3136df8bed2d86", x"6345d8fde94c66da", x"a7beae136ad64512", x"84c57aac5e12f6e5", x"452749ab1c508f54", x"b5399d092648d560");
            when 14560188 => data <= (x"24fff7fe4fd705d5", x"6231fd5a8be1ecf6", x"a4dca4a072f2d66d", x"48db87a3a5e8c21f", x"cdbe31a95f5c28f0", x"fe86c1717f078e80", x"10d1941a8fd0e6be", x"9031d3e70c1e15f9");
            when 33439069 => data <= (x"85adc0e2ccd189be", x"ead47f5a5520d0fd", x"41eb57fffb5f9414", x"a1f1d362bda33a85", x"63201357176fbde2", x"6cc45b19acd1b720", x"6c7d0a77060d2c1c", x"8e7980b60f8db0e9");
            when 8199859 => data <= (x"03e31e3399438141", x"9e1d94c7db144a2b", x"fc63ac5a564a0805", x"d0cc51b1c1b9262a", x"6659f049d296f64a", x"ee2284884a9dd138", x"7da0a1f40a2d12b9", x"27e9ed888cfc81b2");
            when 7555111 => data <= (x"a4608868c4998870", x"232f8e7ac828a456", x"4a3855783d69f678", x"cbe0fa0dffc18b6f", x"51d0804998ca6591", x"c42dd9a0ae1e6571", x"2e881a2094e0e57f", x"c0dddab9708ab469");
            when 2158067 => data <= (x"bb23699df7e840aa", x"556f58e042cc8894", x"74678842e0110047", x"7a7cbcb825352afe", x"857df3e6d3d58478", x"517c7d3423a4a1ea", x"b25f1acc5bb15fcf", x"d33b433b0e69b694");
            when 23778134 => data <= (x"756213f5664ed8af", x"ea0e947c3c53d394", x"f272540747a3d1e1", x"c6500ce990765cb0", x"a21dd7dd35095d7f", x"f72d428455f15ed1", x"af091187c2a1d10d", x"e34e384fdc756ee6");
            when 27801192 => data <= (x"b300ec09e8552028", x"cce6bdb8fe7aacf4", x"21311293d6f0626b", x"1cade364c8aa6aaa", x"6e872e71f8db7242", x"b36ee74ba0111f14", x"461bb8e0ded061e2", x"eb3dc8bdb3d539d1");
            when 11595552 => data <= (x"c92ff8d04d1d4019", x"b18542750c5cafd6", x"22299cc3c9729b21", x"560329900eea5c37", x"2fb00a950f63764d", x"5dd771eadbf7aebf", x"d781ff3e037e37e2", x"e81d06efd3131e99");
            when 20355604 => data <= (x"33ed78fa51824938", x"d451f54907e37709", x"a2e2c2d5d982a815", x"fd35d41668493db7", x"09b3e613ea9f1aaa", x"980e64a8e8928be8", x"af08fea2c944fdee", x"fef7118c62f2be85");
            when 13750951 => data <= (x"d61499a7fb55f426", x"384ad63f93c0b8a8", x"3e79d7c6f03421f5", x"8b80723e04baada0", x"29faac921524ffe2", x"97d552aa4833d768", x"2711ac7d862589be", x"136e37ec99308258");
            when 1777631 => data <= (x"3860b89ad36ffa88", x"dac81a06e536aee2", x"6704937bb562614e", x"ec657c8df228652a", x"2a71013273605d5d", x"d78875e2447af508", x"ccce0f33ccfcac61", x"e1b1d9bd11bf0d25");
            when 22966634 => data <= (x"8d152bce654245c7", x"ac1c93d7b71ab6f4", x"d9343f669ab5a28b", x"a58c51ab6d1abe31", x"3c2d10b1a3bc9b0f", x"1308be37efbde986", x"e088d45cb8316d4c", x"c616ee93ec5bc981");
            when 14296937 => data <= (x"8c4c666495dc55d9", x"24738907ea1d0f65", x"fb3df95fc9d026e0", x"c8f243c78ac97f2f", x"83411f8c9dc7036a", x"df5b2dbb29c9cce3", x"9348e63d54aec6d7", x"de8ee56f31acc9b9");
            when 26809849 => data <= (x"85794f30c655b5b4", x"3b414bba40e48fa4", x"8ffc4d37f87e7841", x"576bf696a2dd850e", x"809a27ab698b9ebd", x"8f6911fc2e60e014", x"b87e09b21849b9b3", x"e695f32ab80b2f21");
            when 28306158 => data <= (x"32096b5f1996035d", x"c3aaf165659125d9", x"89b092bbb3ae0f3b", x"45b48b6fae458275", x"9be7d5c47895b447", x"287d91ec6ac4af89", x"8bb6b9a8af6b3120", x"bcd481367e4a23e0");
            when 33754567 => data <= (x"5682f17045f5a54d", x"a6711affee3cdf08", x"ea315507791d2bec", x"77e0b3ce5511f6b7", x"9e486a459e694f1b", x"b332ce0abae44c59", x"6ea96b5f2ccdfe91", x"da54c150551c3fa7");
            when 7645693 => data <= (x"63bd679b58ddc1cb", x"04676ca96fa4d314", x"4d933678f2ea1702", x"80d41aa0373dd0d4", x"1e56fb6e2cba3400", x"bfa891a949cde3b2", x"74ec89b30305a6be", x"e3ba478006e31f9a");
            when 12262531 => data <= (x"2ba4b771bb2e268a", x"164f4e2c19d6cd5e", x"7228434b8b2e2ad8", x"0229b754518311c0", x"941536c58718b368", x"63b7f53751da8715", x"7c938bd096b201c5", x"20c3f0f4ce8e15a9");
            when 13578886 => data <= (x"a6582120461add78", x"e039d6f032d4cacd", x"b68ed4f4a3f703b5", x"ae478215560ba468", x"bb9872d9c53bc671", x"8c5719124a6f5186", x"226d6b77ba5d70ec", x"293a1ec8f55c9429");
            when 16985331 => data <= (x"182f3b8c7d38cf63", x"7aa4316662901046", x"6130cd3c0eff5d46", x"d5d846edfcf596bc", x"ea2c4c70d0941b2b", x"b0a00bc73410d588", x"72bab5bec6d9f05b", x"66fa62cb181b9633");
            when 14109746 => data <= (x"0acb93c6b3faf98d", x"b484851034019ebe", x"04ecc511835c74b7", x"bc1c432a7e467dbb", x"38357ab11581eac5", x"89ee3cb97ec35876", x"bfc55b06b1bb0699", x"aba645951a563751");
            when 2314422 => data <= (x"23ad34094ec4ce7d", x"74922c82c9f3bc78", x"c708b2cb64513f8f", x"12c94dd6cc69bf95", x"9a48c768075263c3", x"16ce7fafa3fa51ab", x"490a909b3cb4e722", x"58f9c47c92f5fd75");
            when 11210702 => data <= (x"c35b16d57e71039d", x"240edafc0d878816", x"6ced36d23e488739", x"ff6e787705ccc2e9", x"d6381e8e44c231b3", x"50e007ea154b6149", x"d60af21dd34cfc9f", x"a5a3a6756dad0267");
            when 2659539 => data <= (x"fb061b34bccb1990", x"5ee3bc823decba3c", x"85a7dd1acf7f0555", x"bdb7e242bed5eeb3", x"749336502a3270df", x"c0e58c9837127915", x"455413eeac41e7a2", x"205a7931294e25f0");
            when 24407155 => data <= (x"78d53489bb538e88", x"9707744b71eb32a0", x"1690d46a050a39b9", x"f4be74de9bd04b20", x"bcffa6bdf2984150", x"846dc48e69476405", x"11659f22ffee48da", x"811076bab90867aa");
            when 25913453 => data <= (x"baf5475d266f4704", x"2682267490c9b978", x"f84d2b12dacae883", x"13c49565eeb35c3e", x"e5145878f2ae85c6", x"772e2d614eedd59d", x"192ed0c49e1acad0", x"6199c5c72a8c5b8b");
            when 13945036 => data <= (x"deecc8db2baefc49", x"7df611522ec9c487", x"a844e43e78def079", x"211d29c2aa03d434", x"a55469c9c6bb4f56", x"b24e201aadda74fd", x"398ca2d381eef2ec", x"4a6ca0e500e49835");
            when 10085977 => data <= (x"3229502fc8745324", x"7f9ee3a946daa3ea", x"7c529d4a115f5b1c", x"c53b56b04d73d5da", x"5f3d95c07672fa21", x"18ecef3ef9a0f333", x"7824596776d58231", x"4b7710883bdc561a");
            when 11511979 => data <= (x"04ab1529e1496b71", x"7dbed49fcef150c0", x"5d1320ac5c30ca61", x"859a39bd3337595f", x"c6dc94f85ade58c3", x"12bf6eb1ab3c743f", x"cac47106338e1ec5", x"d170f927f788a8ef");
            when 30709555 => data <= (x"e99bb09717164fc0", x"92c9ff3e1760bd25", x"451ca8681440ea7b", x"cbceef8607826b4c", x"f51238e890768928", x"774e01e7bebd6895", x"d44f5704b786fb63", x"4e2d1b43901fcbbd");
            when 16110861 => data <= (x"32452376b0e88040", x"9fc89d634d76b446", x"b390b1834d233aa0", x"23ff629db7011d0a", x"6c6c3680b1627e45", x"ce21fd4c092f95b2", x"4a309a8b42d65a23", x"a79e1549acb4c07e");
            when 10100532 => data <= (x"345830a0bbb5172a", x"2e975507bc8f8005", x"cfa9b0ac49f3d553", x"274e43223227cc59", x"4b338aecc0943bc9", x"f0cd52d13544bf7d", x"efdaf49c4b2b6403", x"5f987d2271fb1a95");
            when 29388546 => data <= (x"53c9efbca37b30f0", x"d78fd53197057ed2", x"e41b4b09cc2af38f", x"a354dccff3bef614", x"7f07385629b5b146", x"8205b3eff2a8d9a6", x"725e2112207edb6a", x"cb437028ca2f5da0");
            when 25063612 => data <= (x"cf8cc6b7a9f2d5e5", x"72b86092ef030c3d", x"9d7a2d9b6bc0cec3", x"923bab53210a147f", x"5c381bcd6966c7f1", x"f48bee789d37aaed", x"36d2d15acb46a94e", x"eaf5c1bcab19474a");
            when 18762865 => data <= (x"1643442e8fb4413f", x"ec9f68677c4875b3", x"aaf58477819936c8", x"2f85157b3608d479", x"67fdefea91da1ecb", x"94386a32ae21eda2", x"58e0512e374ac0e3", x"1084374f8d37bc63");
            when 4048435 => data <= (x"22741414443e3652", x"5c720bd4c6017c14", x"fccb4b2951f435cc", x"0564f37fca66a26a", x"34478addeec44d2b", x"e6a0accf210959ca", x"4d95b7bf20950fa9", x"47f8f6c51caa8f3b");
            when 24585583 => data <= (x"ed67cb38fda1265d", x"2bfd7da90bcc4838", x"96bfb2d89fc1d186", x"b5c925a184d3fe25", x"4e35c5019fed0004", x"bde05840dc81ba6e", x"66c3296f1b529331", x"584768459ff01073");
            when 16053275 => data <= (x"0319550c97077d37", x"b5247802102654ff", x"4eddc14529938a19", x"9bf111272f7b6990", x"dd0a4658df334385", x"900f9e7cde2cac77", x"1683562005e9be4d", x"c2b7efe10d8c4040");
            when 13349063 => data <= (x"b4f58cbb4b60ffad", x"275108a5f932ad00", x"82686d901ac28c5a", x"1bc7956893465fdc", x"0fe8f4f533de337d", x"c75fdf03fb7831c6", x"cb55b5eec69593b9", x"d2597e82b03e846e");
            when 6345569 => data <= (x"d304434a3f3e09fb", x"88aa1ae14f5c2179", x"34077880e416c879", x"6cb2d79700b60a2d", x"19f15c295547a2db", x"6ae441b518bfdcc8", x"4f2ad6ca16ddf945", x"a88ec92271e963b5");
            when 8593647 => data <= (x"8ebee1fea55593cd", x"1e8f3074974fc8d3", x"c2c629b5ebfe94bc", x"35567ec01d1de51e", x"a4a7d4d2b044fba1", x"196e533b1ad6a8fd", x"f7ce01e4ad95d33e", x"f9d909e3a319d404");
            when 12172901 => data <= (x"e4fcf1fb7f411b40", x"e34309526ae31174", x"4af24773c21f7020", x"8dd918097fbc2e92", x"593fbaef0f218d27", x"ddd428aa8ed48f89", x"fa96e91d80b1d8ea", x"01069e5ba457c620");
            when 2531790 => data <= (x"8456db5d217a7bc8", x"3b28daf940a3b579", x"0e99a11a86dc1276", x"dd3affc946364974", x"0669c7a2324204b6", x"0bfb10200a29630b", x"73e356051533f027", x"fa74654b5c77070e");
            when 20303352 => data <= (x"0019478d553bb3d5", x"7851d2a34b62f59a", x"6e8a81658f574d5d", x"dadf24a01a7e4951", x"e5282e8dbda46a08", x"57913231907143fc", x"960c6f9e2b8d504c", x"3daa2206834eb25c");
            when 7885354 => data <= (x"50b336ac60362c58", x"8a0251ebc949068d", x"aaf2c70282481356", x"ba41b57e5113f9ce", x"4e1efa7e18e3ae1a", x"8c8731a4089af30d", x"e47d45b735fca70d", x"10043da86fbdf145");
            when 2678344 => data <= (x"b0f0513cbbdcfe50", x"9b2d4981b2760751", x"49bdc1cdc96d4ae5", x"5838d3fae44c5383", x"98021c18fc6eaf45", x"825775c9996ca834", x"c9b1577413fcb53f", x"6d987cc366ded733");
            when 16223871 => data <= (x"a79aa62927c3ac4a", x"eb9f26f3563122a7", x"a3e0ad417ea0d385", x"cbd7ea86eb9c7fa4", x"f15edaab2105aab5", x"1d8aa2e864a50904", x"76f6ee68c5ff9d63", x"b5d60ec3a2cb194f");
            when 24429781 => data <= (x"fa7663715e496e75", x"d2075cc6e8e2f51a", x"9c11af272f818244", x"9292b45de3f239bb", x"68c7df6824a9d7f0", x"f9c1d2297ef7d0b6", x"413ba5bb3c04bebb", x"f477e514adb8ecee");
            when 17053177 => data <= (x"d7ce0b004889b70f", x"cf7306799e7689ab", x"cefd677adbecce2d", x"988ed12f4aa31f0f", x"695f75e35ab6ad23", x"07a4e110470fe7d0", x"e0eb95babf3d00be", x"0c0b489aed6dd2ce");
            when 28757943 => data <= (x"0624d9f5428e287b", x"dcfc979288d07c76", x"7e7aa3ba4c1d4339", x"664dad640e96d085", x"dcb43d3df63f5257", x"71e0e17c0c4bff46", x"93e1e1fdf0e4c0d6", x"cfa4e6cbdedc2b3c");
            when 3080894 => data <= (x"5cc5feeca286cbe2", x"c4324de676623450", x"06ae95d83a9c6b1c", x"2c9242b57bf4bfb2", x"8b78285ef2cd9441", x"2562e76924701cb2", x"45e1d8b92db9de4f", x"80cbeade66d88a35");
            when 19601663 => data <= (x"37de28d5bce17f23", x"acf0a10197d817aa", x"3e7fd990d53a3217", x"a99e70626748851c", x"ce20e632846c1ca6", x"c7db2b2b2fb6a72e", x"cba1994fdd3a840c", x"ab9cc9021626a259");
            when 825727 => data <= (x"1a3e8c7dcc17c7bb", x"5b966cdb7a06127d", x"62f7106247f30ac8", x"ad5776af2ef5d9b0", x"a0eb83ab02343310", x"3c94a16843f0a1b5", x"7e1139877fc70507", x"0138b23a40033a10");
            when 20697799 => data <= (x"2a57bee2d6036a1e", x"bace44b1cf481f9b", x"7f415467075deed4", x"8e020d32463d12b7", x"bfa9f21267bc9d67", x"43fb6ca4d887f463", x"bce0bd387799724f", x"a5c732ea19c1b292");
            when 2820122 => data <= (x"0677c955d73c008f", x"d0053c75580b501f", x"f8a5d6502bd37c01", x"cfc2974cd550b32c", x"59d687951205c931", x"505306311b680afe", x"3c7ececa91625820", x"ea7f32bcfeeefc87");
            when 19372915 => data <= (x"a163669de1d6a226", x"8c7a964993669d22", x"e99c3b365602a198", x"2e8dea2da0cb77a8", x"356a590eb817a97d", x"99d5e4e3e6f63453", x"b101b5f573d0530b", x"fb7eb89fd9cbb4a1");
            when 33819301 => data <= (x"2bd48d1ba1476f32", x"dbcd12bc5894cc1f", x"4c0b3333a0b26d32", x"da4483656802d6ae", x"5a65a03641f3534d", x"e620d2a37b0b8001", x"0cfcc428b9c3098e", x"23e905d4ecec12ef");
            when 26849320 => data <= (x"07e4c554a9a216c9", x"c3943cd0ca3fd744", x"a25d0e72b67570be", x"a481545150b92333", x"d84b919f57a78902", x"8349849143a43254", x"54787a5f2319df99", x"6e5277457a54d67c");
            when 10759182 => data <= (x"2445a454dd74145a", x"bcaa4ffc18cb62ce", x"3209c63f94de22fb", x"0497d08fd0f4859e", x"f5912509cf5c3e89", x"dfd1eb72a08a3b69", x"5208d90bc0a202f2", x"a1cfd00a1faa49cf");
            when 13126981 => data <= (x"562c21d5dec21f02", x"8e937c76544825a9", x"bbf55992b0f6e43e", x"b9e0d6b1aa703173", x"83550e4f5fce0578", x"d035b7b9452c7b77", x"6a251713c791276e", x"33c25cc452628689");
            when 29562575 => data <= (x"e823e998cd8a5aa3", x"afcbce47ca32be9c", x"34efb87254fbdb7e", x"77c8e9ba78ef8b92", x"8848a8723ac1cad7", x"86089bf784f9872b", x"9c3cd3196c4abab6", x"6e5325d7b366e884");
            when 9225194 => data <= (x"8079cbcdd1938440", x"1a83d15c52aa5ca4", x"282dd31180ace2c3", x"56217bf467134f23", x"b72c43c1c0e5f1af", x"79bb0195cc334fff", x"d42f4fd167ad57b9", x"06605b2e894ff19e");
            when 11241655 => data <= (x"244bb02f0058bce8", x"20758d1508097384", x"7ab2595d584491a4", x"9707b9c4856e13d9", x"69a1dbaddb756645", x"7298a80e63b1407c", x"c2f70dbd5a8b04b0", x"26ba5a9d93a7ea52");
            when 25870445 => data <= (x"6e012151af6ef357", x"2eeb8a60e3f1d55a", x"450d0ab63a4b79ee", x"c3db429613060ade", x"6cdbf31a5ce34732", x"dff71379fe8677f0", x"32b8eba6a3c5d5a1", x"441a7c0874618de1");
            when 28128149 => data <= (x"a11decdbadb3e9c1", x"3d6e421806db1078", x"199685c70121c022", x"1dc8ddfbc84e00f0", x"93f2398440bc8839", x"b72f4c069e860084", x"d11ebdffdbff5f11", x"be1175e750047f0f");
            when 4169815 => data <= (x"825dd8e1e8c447db", x"08ae4a159b888f54", x"a50b9be921e21186", x"b4dd0a7f27ca32fc", x"0e9b5cd9fd5de07e", x"b84ebe8e87249b94", x"baeac7f51a6ff526", x"8dd68ee1be81d1e8");
            when 7336396 => data <= (x"287bcd3ca731b2b8", x"b7fe7a27b41f8fb5", x"9c8c1e826e0b6b67", x"3b646da42a5dced9", x"d1f4df6937fbfe79", x"2f60d2a37b1075c2", x"ebcf5c3efad7e3d6", x"d6b11ceadc386556");
            when 16511583 => data <= (x"2f4793e70fc8b59d", x"a04539bcae78bcd1", x"ff3dce3cdff3e75f", x"dfd220cb4e78ccfe", x"542878d53c84deab", x"8970e584188fe40b", x"5dbb2f583484f200", x"a7d86fc4326ddab8");
            when 16954699 => data <= (x"5ec80c1adf9eb19c", x"f51b77e6dd7acf1d", x"a1c480d79a455b19", x"2c77ac87da8be033", x"093c7cc26a555be4", x"3135490aa0a991f4", x"c20641dc3ebd7038", x"214821066ba2d513");
            when 1987435 => data <= (x"485b633350d23370", x"47ebc6ccc2e5351b", x"20e03b43b75a723e", x"77fcd015c12bfb54", x"a72d3c76b0f05e1e", x"b742c86d751dbe93", x"5bc1a3da1442c671", x"1c440b3ff0553b59");
            when 9371189 => data <= (x"9bd3bfa1400fb953", x"e13ed6d172b6f851", x"d3f001294ba2ec84", x"e62e358ccbcb8dde", x"2776c280bc06e552", x"43857b83b5731504", x"420561abd886503e", x"f3ee4079e9e6c870");
            when 6531161 => data <= (x"2305c9635b304c01", x"612a6015749cf6af", x"21ad44641f5cc242", x"f87181596c8e10e2", x"9e1f4b0056dd1f5a", x"515212f2ede3ff4f", x"964402ca761b169f", x"c31d212b2a675ca0");
            when 30259414 => data <= (x"23c66e53df5fc6d3", x"b433bf064e409b80", x"dcd145aeadf0d124", x"57110abdec64d12b", x"1ca7b8d2e7b9131e", x"f47046df57a25f4c", x"b2fc03d9973ebcf4", x"573d761efc28fdf3");
            when 31613125 => data <= (x"70fd685b4725d088", x"af7fafcc78c3f434", x"382752c1cdbcfd43", x"228c384647b4937b", x"dc2ad93d142774a3", x"7a911f090fe9c69b", x"59905fceb5bb19cd", x"c33b16f2f40d101f");
            when 27546399 => data <= (x"6ebd6c9cd11a45d3", x"1ba6111b608ee5e7", x"5958afb32ce68e90", x"790feefbf4be6a0b", x"c5a76e8e299ad02b", x"fed7df5d79efd8da", x"7ebb354cff67f59a", x"ec1a055620f82b0c");
            when 13808519 => data <= (x"0e6b711b57861105", x"0108677ccc8eba16", x"29b420eb919acef8", x"8dba4955b5674123", x"f784846876bd0c32", x"768cf279e5a76e75", x"2de8fbf88313cbc2", x"e8b9bc7fa0b98ff4");
            when 33488115 => data <= (x"22bcfa32e1189b4a", x"830bdc24b83d4e8b", x"0dd55997528ffe95", x"9e074164b818d171", x"694dfdf335edfc2f", x"5f695703749b535c", x"4c8e621a0d360817", x"a6a162c5fc3278cc");
            when 7117313 => data <= (x"3708e52648a374dd", x"bf2828b114c4bc6d", x"e8cff19cb4d84c6c", x"91996e4c3dbd8bac", x"1610e7306ab92356", x"243ab357b4df6281", x"c0d815cdd28a20c5", x"b667a12c73ffa183");
            when 2030370 => data <= (x"41cca3a66eb34062", x"29a1ea26a1a1cf1e", x"bbf4a37485e85205", x"09ebf288987a31ba", x"4ce5b6b873370737", x"e91647ab1cf1a942", x"17acfbefa51dd08e", x"3d6a5bc8389dedc9");
            when 27465336 => data <= (x"98d2a79b4e21bfb1", x"b7247a7c8cc55b49", x"6cec116bf9484b74", x"4f643816de1dc5f3", x"79a45f18b6cbcf52", x"49d8b5c9d591e436", x"7adab9fa100bf291", x"3ce1a55b16bf43e7");
            when 8672832 => data <= (x"50695c8e4603d5f0", x"fb3bfbb1260de37a", x"5a4d389f6f0ac9a2", x"a3661d1c187c3488", x"fd1410c1750acd90", x"e493590481b55e32", x"aa37c9f8b721b1f9", x"48afe6673ceaa5c4");
            when 30519937 => data <= (x"ca1e46e08266e60b", x"f961e67bed12ebc0", x"630bbb9d095fab2a", x"8cd3537a45efdd88", x"9e4c2d8ddbe8f6b6", x"879b1690553e6550", x"3f36b6b5fa128811", x"d8ba995229eb8a4d");
            when 24635237 => data <= (x"b0b5738c1ba28767", x"f89daf2c999d5078", x"be7d57a4b358b9dd", x"0da6669e9e9b5b6b", x"b26ec154fdc2284d", x"16a29bc092b76f41", x"8095bf888b7a4693", x"8694a4deebd59553");
            when 13444128 => data <= (x"593c504811336793", x"8b45a0890ed1fb93", x"10bc96f80a0a4596", x"c6c6019105964e18", x"03d206bd53cf15e7", x"8b45413beb0c9665", x"0bb7d02e65df2732", x"bb77b0bf30500300");
            when 10103564 => data <= (x"cea45d4d51447cfb", x"d89f7953423e93c6", x"c1d8370d2b734aaa", x"1c4122156f85a97a", x"639254418910c231", x"732a4d1f6ccc996a", x"f43cc2bd517d7db1", x"2bd536025e1a6118");
            when 3918686 => data <= (x"b109028a7e58ce5f", x"a23f8a2a5203c95a", x"27287acbbc966c55", x"82b7d68725e31f6a", x"9d9526499ffa5c6c", x"1315113abb1f1160", x"5d6fa569b76ca888", x"6059a5de91969b78");
            when 15043395 => data <= (x"c34ed081b87e7940", x"18b6f43f99e15af4", x"cf39575d6bca1336", x"31e9fc245cbe3ae7", x"413576b2a6f141fa", x"d50556a40c649389", x"6606cf9455bf8a24", x"913cd73b8e656b44");
            when 31446579 => data <= (x"d9f315c03922924f", x"cb7e750ac06f07dc", x"0ecc949247c31eb4", x"d07424ce03a31721", x"106e1bd5936be1ec", x"f0cb27beeac74b21", x"b7695667cd064e77", x"711465b006a55fa3");
            when 32705443 => data <= (x"faa938339e39ea9a", x"366d6c0f7b79da9f", x"4a7694230976b9ae", x"07f26f3c6db53953", x"990ec58ca1a4c234", x"5fa4a5f781d7d09f", x"f7b81407898f223a", x"077b18860e6c1440");
            when 23466376 => data <= (x"b5daed01ab76ef83", x"c0a3cc179620132e", x"4cc5c97ddfff6bdd", x"9435051c7733ec41", x"a56b1b35895c7faa", x"751caf770d050091", x"b17c7ddb3f81e26e", x"1da895a4bda24730");
            when 10952259 => data <= (x"5c9b82f6977dd076", x"d1ecd269002129f4", x"7671175b64e13448", x"f318018e60cbbbd0", x"1d58e6747897c92c", x"c9a61fbfde8a21fb", x"46de5ea4644f6995", x"e39098ac5253f0c8");
            when 33771209 => data <= (x"a9a7b6a1f99cf10a", x"a600eb8748fd659b", x"5a78975c6f06a58c", x"a2c9831dbf2c5156", x"321bf7ef12f43389", x"131dd6ee0bf528c1", x"272e578a6543c15a", x"26fbbc2ed70a33ac");
            when 20521788 => data <= (x"8802e605477932af", x"cd87e36ab84e9008", x"d08d70d633bfd738", x"9c241a2b3e93723d", x"8334b9b2a9befbfd", x"ebe728f88c98501a", x"d037f863b366cb85", x"5d4907b5200d77e6");
            when 14847773 => data <= (x"46df9d1b4ee67e48", x"5c91c0bb1491fd9e", x"ba0d1c33c74ed7ce", x"db2dbbc6eab61f9e", x"a256a4d371e5d75b", x"761b3d091dfc7099", x"3934dd13526838bf", x"26ff5a2af883021f");
            when 13306884 => data <= (x"28cea22d110fd0c8", x"f99aaf293f7fd2b5", x"981476e45f459927", x"f90b90c05bdc6450", x"abd1ac01e73c8bf8", x"36e8b5ba834fdc09", x"7b9c1b7fae143c72", x"8ac54fb27acfbeca");
            when 17418023 => data <= (x"0787775dfb2e058d", x"ddceeccfc856de11", x"feec9af4094f907c", x"ec440553b7a23c3c", x"e6414a5e14260c70", x"2c0bd5fd33e40641", x"a2b34f4e114f76dc", x"82343d09e130c360");
            when 6574670 => data <= (x"af79190a7473a190", x"276ae3e131634f41", x"f4de7ac07039e2a6", x"c46e0542112866a7", x"cfa94d8bad955708", x"9864d2bade7b0d95", x"fef704eb291a03f6", x"a414b3b6ea5d77a5");
            when 33748130 => data <= (x"a29e022df9ef4560", x"7ca052dc0e901866", x"7ea719a6e91547be", x"420577b066aabd5e", x"f99ebd8a1815def3", x"c57c1a0fb5bb1f72", x"2981907177dab85d", x"ee129a4c2a3edbea");
            when 10191028 => data <= (x"75754cad4bda409a", x"f577241c069a6d28", x"573856e1113d8775", x"215d4ef763642e49", x"ebb6a643ba6bf97a", x"b53bbb74f0b320f1", x"62e73c42f4981387", x"c9b23f1b048876d3");
            when 25727860 => data <= (x"e16a0ae9512dd9ef", x"70e507abdb9ae6a0", x"5d907ab337481b20", x"6d8a7dd6d9941bab", x"384ee65b776d8d65", x"e5018d1f935e4481", x"88b98815166f06ed", x"0a1332450fa89d3b");
            when 26891759 => data <= (x"f00aac83356d0364", x"a170cf590f1a1360", x"baf22cee651c68c8", x"3c96df1598bed086", x"aa675d54c83aaeee", x"b41eeffd603f940d", x"cd624dc6e9b0961b", x"78bdfa7b4baf164b");
            when 19574675 => data <= (x"9235605b7359d777", x"2e7d1d144e819b43", x"deead5fc35733cc4", x"aec34df77ba5143b", x"c83a247cf1a26577", x"ced16fc02ef3da45", x"2b145384a81b65c3", x"0b6ea5ab38c1dffc");
            when 31414814 => data <= (x"edf563e7fe28859d", x"63e207626c357bf1", x"119a969533766414", x"f007921d7b0a684d", x"a78c59a126c4039c", x"520f59f858f71b36", x"313ed6bff6a0b138", x"1395146324064a46");
            when 10636976 => data <= (x"f369986fb15c24b2", x"393a513d50566d14", x"4151872bd0f30cbf", x"1f58cb66665ba7db", x"d8e28fd23d0f322b", x"2502c4474886a828", x"446f8d873cedfcb0", x"13f0e108e75faf64");
            when 11583277 => data <= (x"713214ef5a466602", x"f9ea0ea1520f9d38", x"26256260a4541818", x"e0e5beb0fad765ae", x"f3ee167e4f3c96e5", x"0628298cb30433e3", x"e8e63c6520bbdb57", x"bf5802b83bdf4d0e");
            when 22398792 => data <= (x"cc996aa88313a7ff", x"c4c777a5ffbbec1b", x"e986f440462fc5ec", x"d00564cbc5449632", x"c6e5bfdfd12b6ac6", x"835e6ce8c69ef6ec", x"b05ac909bb13437b", x"e6f13d34abc9f84f");
            when 21411656 => data <= (x"c6194f3ffbd37b33", x"f688233b37acadc8", x"23e7877155b72d15", x"5907fc6e08dce836", x"7555fb0b1dc98504", x"a0cbd286da04c8c6", x"66328f5f71d343c8", x"85be295f53ac0742");
            when 21836912 => data <= (x"0a34481dd7a5e450", x"04189e54a393836b", x"4777c933afc39361", x"dfa8415ffcd98cf7", x"2dc6e505ed53e4d9", x"c77da6e8cce1d176", x"846c811582c42535", x"5929752274e27431");
            when 13185469 => data <= (x"7b352ce374964500", x"3f55acf896d97f57", x"1e8957e7ebde5d00", x"d7ccdeeef348a875", x"117f3e061f60c19a", x"647b0b1165691dad", x"87733d045c9c5739", x"2325fb4ea993447a");
            when 11329495 => data <= (x"4d10debb7c37a1b5", x"e63659ae83d9527c", x"6ec915ec8c69632e", x"3d3a5b7160ed044b", x"1e5ef466ce7c732a", x"2c685296a3acab94", x"d31aa3d93df11b88", x"09e9f9023dcbf706");
            when 27833275 => data <= (x"b8245bdc230c3512", x"bd27ea9f00aa1c03", x"f059b9f8116e5d56", x"9fd5c240e47a57a1", x"708ebc101f26eb39", x"640a79ea2f02aa31", x"ee25762396435d29", x"0d402e85cd3d26a0");
            when 25025630 => data <= (x"f71a5bbe59d2a529", x"274f5f642c0d2433", x"a1cd7b725a0a9fa0", x"1c7846dfc432f7f1", x"aac65c5c620b2be8", x"4a1b02033965a040", x"f7e35427b699f5c0", x"77d79ab21b97f325");
            when 18242799 => data <= (x"744f9487dc655938", x"71351ad4fa5d8fc3", x"da5af64849e52534", x"511b0728aa4e553b", x"3710aa773a9f47f4", x"2f439d35f8c9739f", x"fad7fae5c46cb3e2", x"0001b06ae1cbb6af");
            when 10892647 => data <= (x"a2ede038c5fe045e", x"8d731cda75c8c370", x"9111a9e6ca3c89b8", x"e34731302c010798", x"eb7b4c62038dfbff", x"f75a90ba21f69cf0", x"2efd1166c8c4e2e5", x"85d52a2676225160");
            when 26562934 => data <= (x"ac8adc617db0fd73", x"0c5678c14dc57175", x"40427d3b0288cd2f", x"d1b4b0510543ff12", x"2aab05077e47e6d3", x"2d5cc9a991be0b1b", x"9dd25f66e40e44e2", x"ddd86599cd6e1601");
            when 33868767 => data <= (x"b8eea41afd117b37", x"fb9de21afa92c0dd", x"42ffe80a003804be", x"f15ac8cab9874658", x"d4dbbaee683da820", x"bf6d4b3eabfb5bed", x"663294c3ad8c87d2", x"226d3ce649ee62e4");
            when 20727619 => data <= (x"7525432038c01660", x"f1065116c0adb921", x"7ce2de46ccd176bd", x"0c6d69fb5cf31c16", x"c37f17e729d55c26", x"6506d7bb01dfc282", x"ac22756e3163ac11", x"e034aaabb66f7c5d");
            when 33041276 => data <= (x"a33c54adf4659e29", x"02e6d840d4c90dc4", x"78339eb69a61614f", x"04bbcc258b4e0b60", x"a0b461a528b9fe3a", x"0b35e6790a7eb4e4", x"2bbe42917e1e959c", x"b9df5c03e87a9735");
            when 605797 => data <= (x"5b85a87a57bea247", x"81c7ad5c4c6b1df9", x"6f173a9ff2d25e38", x"b009630b752c7024", x"eb7945576f9561b8", x"6de2e05cf1251535", x"82318df8d5e87ea4", x"b76fd9874a7432d0");
            when 20937559 => data <= (x"9d1c6d698b4fb2ca", x"edc72e5c9e7f9994", x"af84f7440f030fce", x"98929119a7d1fd13", x"89a0557cc22f560b", x"49dbcb9ac79d6bc9", x"9e88928fd3725ecd", x"99dd3c497f6ebf11");
            when 26921692 => data <= (x"068b0cef195f5088", x"c3461e75892c95d5", x"5e8b4892378abb02", x"650dcb3b9ad61b22", x"f89f352b156d2231", x"a57ca5f9bb406f4b", x"4b4deda5c6456d78", x"cc76fe9de4f4d42d");
            when 22933756 => data <= (x"b5afdab17efd0557", x"77a74ee9927853c4", x"1b9c1ecee084770c", x"9f354e27c8e517cd", x"06af85b74d7677e2", x"d1b6b74ab53b8edd", x"104fa8882d22e0d4", x"d17115819e437d17");
            when 33836170 => data <= (x"dec1670df6939864", x"5dc1b4ed6e1084a5", x"c88a52022da61c56", x"0ee684821404ed9a", x"99a72c0ac6a7cc61", x"708d7ea35d636d46", x"38fd20cfe87d6415", x"79855b800e5df068");
            when 900862 => data <= (x"88a9acfb5906d027", x"520375c965094169", x"3f94e7308cc229c3", x"a261424b378bccf6", x"16f1fe9c29b4a5dd", x"8aa6bb66f56982b8", x"518f9c49fb97bdaf", x"37b384df682a4714");
            when 1907122 => data <= (x"405ff31696803b9b", x"59cd40f4393bb83e", x"f4d9a87260202eff", x"b259ced780a84a93", x"962cf10646351ed0", x"9ab38c503c2441ea", x"ca7208f2d15c7ef3", x"c1c270b9e64bc85b");
            when 2144395 => data <= (x"45e27c81f331d327", x"3062a874b16b06af", x"55458b6626659c29", x"4b41d140a3b307e5", x"ffc80c2399a5cc52", x"f59d2125eea3d1d9", x"f062e1b3196b0f11", x"8e27dad0065afb4a");
            when 28135190 => data <= (x"37c3665153c84978", x"41981b0ef989a413", x"7164a7c914a61bcf", x"8268db3df5ec7f46", x"2e4517fd37ad5664", x"a22c2a126afdd15a", x"6779b252b85f7d87", x"352dec209029e4a8");
            when 25219529 => data <= (x"3f81a6b129ba58c3", x"4345f67987bd902d", x"ab496a827fc156d5", x"a899e449da35bc01", x"5de98155e9505dbb", x"c2783fb121c349ac", x"c57efd04b9ef7edc", x"115176cf6e626238");
            when 22108910 => data <= (x"ab7f724c61e2081a", x"e426341f9b1fc12e", x"3acbb7cc9001685f", x"fd13478dbf9ed568", x"88c5bcb7f833a79d", x"f9bda772ae75afc3", x"cae6c3d96cb6c096", x"a2e8feb594888022");
            when 26715761 => data <= (x"34c9c1981955451e", x"6775ff75178d37ae", x"06f3643d9571e677", x"2b81c5b2e64de148", x"c1b96b1c9a252f4e", x"13af3b472a7fad83", x"458c850201235da9", x"a392a12f32399576");
            when 7318548 => data <= (x"f63a65cbcc0f4fc4", x"a8bf3723f1d04499", x"1b3db60ecc3e3025", x"79b407e61042203f", x"0dff1b6ebadde701", x"7954d002977e920c", x"f944cb9623d43552", x"196e875d6a10cf28");
            when 6855632 => data <= (x"1788a1da208df686", x"ce042b0bf63bd1e9", x"05a9bb5594f00daa", x"36cc5f6013c2ee9d", x"2c6a2624c6af0636", x"dddcfbe9542e9bce", x"868c17e8900e8112", x"995e5dbe912e05af");
            when 17392148 => data <= (x"f70d1373d18795c1", x"9226c64390c19e23", x"d66d2f578c1de546", x"9fd5757a17868a49", x"4373494abab5afc4", x"13250d94b35113a2", x"fad9f0dd564efd01", x"5e0e74df00905553");
            when 5041099 => data <= (x"18eb17f30383b762", x"03605c608add403e", x"5bfce025b7dcc3db", x"015ab8b18f9a405b", x"bdfc0fe2ce20c15b", x"ab75b815c5b8e328", x"067d779eef56d2b8", x"a3b0f9d609f87594");
            when 14859012 => data <= (x"2fb3f62de1c6f873", x"67fd24b31eea5908", x"0a895437b5b26b2a", x"40b8518f8c57018b", x"9fee761a711a7b9e", x"c545ee665d1171de", x"33973ae2b861355d", x"b89e55d5d2c932eb");
            when 24310885 => data <= (x"a7869ef6cb4ebf0d", x"ff1e6891e51320ad", x"5d7a32c3724bf56c", x"affef96417d0533d", x"d7cc0bb43af7bf47", x"f2cef692335fd040", x"15d71344b9041cd7", x"cc034cf83c58da3b");
            when 13007277 => data <= (x"a37e8191949ee3a1", x"6ef18a64a47ba72a", x"6a6101427f442bb7", x"7139e83d4e30be42", x"9486e36726ade4ef", x"209f819a1e4e0559", x"c05ba4487c94c8da", x"e039636a0ee72a9a");
            when 17749297 => data <= (x"23ab93734bc127ac", x"8dde8c8638f2a38b", x"b85fb9855021e817", x"3fe4bb64e54d711e", x"d807bd30fd3c1f3e", x"5f4d3cde87bbcd19", x"fd6749a6fab32a82", x"d69ea33d3eb7ed40");
            when 29628080 => data <= (x"bc43a0b7220578c3", x"e13d33d567b677cc", x"4b4270cbb0eb3132", x"3d54981847890d76", x"0820b11aeffdcdc6", x"f9a51e5684eb9e09", x"f24041c972a6f4ae", x"d9a4f4cc9bcdede7");
            when 33341314 => data <= (x"6174b360edb3b2b6", x"56a5cdc6aceb367e", x"b7bb21f4921d77f3", x"9f13b3e96a511dcc", x"22559d8bf8296c56", x"8ac63dc89b1a228e", x"eb34ed1953aebb4f", x"e66338f2928ba3cf");
            when 24241189 => data <= (x"b9422757a3bad3e2", x"444c664157753954", x"31dc47ebaef49881", x"791bd4c677f0c559", x"52d124617fbf9f9c", x"477e39bb6c06799b", x"162fbeaeadf94c6c", x"d95e5aebc324af64");
            when 21470131 => data <= (x"d670a4a3c29eda35", x"3017605f0202d62d", x"3d41cb98cd25a4e9", x"8bef96c450fdfb30", x"a5f674306fd0d252", x"973d5093879fa61f", x"51b12e5f43b32770", x"b5eacc2a998e0bea");
            when 13347056 => data <= (x"ea972e38381345cf", x"8b4ce65bee297d1a", x"95a2d6615d2f674d", x"d3a005890d251ff2", x"0cf95edcdf119ae3", x"af47c99a1e278f6b", x"72b8385726662fc7", x"01bca4def180b1bb");
            when 30904991 => data <= (x"9d06e3861e6de77d", x"9f9cbd89cd3f3a0e", x"f7fbf822e1b54d63", x"5461b44082ea5184", x"4da8bf53376547e6", x"e3180b98759fa6d5", x"8221c44d99e13942", x"c4cbbf7b6281d315");
            when 3112496 => data <= (x"f223a03dd65f6074", x"947762ee9ff81275", x"09109163044b5c9d", x"1f443ac493e5d968", x"9480a459a66fd2a5", x"4ad3e1cbb261a120", x"e20fbe080f2eb209", x"205b3ab5f10c9ccb");
            when 24931681 => data <= (x"b4c12cf288470610", x"20afb8a50ac78d2e", x"56adbfb65634f930", x"5cd36681bf358022", x"e56bec0291e8ab61", x"0fca6afb4c1962c9", x"834731284362c0f8", x"03b1161a0b5984a8");
            when 16743531 => data <= (x"f191f65d7a3f5e6a", x"4cb91537437ede44", x"af9eb6b6de0a930d", x"20aa3c623b4f4faa", x"25150d1cfc72c948", x"270bf070f8560368", x"758c1c94049732a1", x"574893407b69651e");
            when 17482407 => data <= (x"22d0ae36a5c362c3", x"6d0fafa5d0de86fc", x"27de6c7724f79ab5", x"235535b243f75c87", x"f5c69d9fb52bc607", x"9504faf0f0f28726", x"2c74d07e5dd878a3", x"13c469c8ff8ab432");
            when 24248738 => data <= (x"5e98bfa73d408f64", x"c92d44338ffc2c5a", x"d897952b72b42937", x"5cf3a1a009382ae3", x"9137a7bcd3535947", x"59523ac4814f8d99", x"24c8ca0d36dc4b61", x"9c242e985cf12687");
            when 14149196 => data <= (x"06cb71aae50887f9", x"5819f4680b7c054c", x"721d57774955b915", x"b350afa352ade5fe", x"2a6809c0d342d85a", x"7acf85eb1b8e20d2", x"af5a27d660cf0386", x"437111d83115159d");
            when 13284462 => data <= (x"e0cb65889a411e91", x"38332fa06f6976d9", x"b02fdcf01596097b", x"e7b8d0081c9401c4", x"ce8776d3b44f2d98", x"50c9517693ba4afd", x"a95fc221446b1e0d", x"740263c0297d4c54");
            when 24058819 => data <= (x"e011636531508b71", x"46c7888fd1ac6f55", x"5b2ece493f03e81a", x"36b9e771d71ad123", x"528c35d3190eb287", x"2502fd1046e53f4e", x"f4cbc665052ae3cf", x"2ec008f23b14763a");
            when 16630800 => data <= (x"233b40214277f48a", x"9f631e87f66cf18d", x"e6884b3733374657", x"a6e9efe546e11038", x"bfd5ec61d3b901d8", x"33563ead32be4ffd", x"829756ab1300c620", x"71d1b7b80175e0b5");
            when 6244381 => data <= (x"de917279e88816f2", x"5ca28b93b862223e", x"75ca13d3c1436a90", x"b2e312fa5becc021", x"ec8951b15d71cc96", x"2c0c739fb0765645", x"fb5272eebcdd4f00", x"431e00fa0e3643a9");
            when 28513167 => data <= (x"6c8692a1cdb784ac", x"27d47d1fc7679218", x"1a71c06f74c8e399", x"f89360d2dfd94298", x"edc1879509ca58c7", x"395a6bf1ffbfeee8", x"b501b23eff13199c", x"6c1f933bdb5e82ef");
            when 27865022 => data <= (x"a4448a384f4dc621", x"9489da53627f13c4", x"da24f2a718437fa8", x"9b16dd2e6900e71a", x"7706ccbe47d02736", x"ffda14eb8ea2d7d0", x"7d2aaf9eccd3a1ca", x"792222854b4d1742");
            when 21684252 => data <= (x"7e643fef44486f46", x"f349d9d8adb32c5b", x"c621d15eb0d1ffd0", x"5be12b9ad073c975", x"d4c9505ff0a099b2", x"a018a7c5f228e73a", x"12a3538650a5b863", x"7f25f770e39c6734");
            when 17000318 => data <= (x"d2ad815fce29cf54", x"afefe04bb2a66183", x"8878423c479c88df", x"c7c640c5ea03b2db", x"98d33e3a06722d86", x"725971f124205f87", x"33b304508c1c05e6", x"de44afe071a8c374");
            when 32487055 => data <= (x"966d76e35e421c88", x"6b317b91359aed0e", x"346764fd21cc296a", x"f1454e451eac826f", x"b34c234c6fc0c8c9", x"73ee890c51bea5bc", x"18c18fee6202763f", x"16aa968e35f27c20");
            when 13280280 => data <= (x"e0a2c1ec44a6363a", x"d9a972083cea531b", x"61113ce1ba6b5674", x"398f4afd0f500385", x"4477dbbc7698d4d4", x"e2b6e0dcd5bbffe3", x"bf87e331cb6df3de", x"8e75242404d57267");
            when 4891754 => data <= (x"aa109228de8327c9", x"d80b3f93c020c922", x"e648be088bee4b42", x"79283e18e7045c11", x"81045a533112316f", x"73dbcf3f668f5840", x"803a56a4c0265f63", x"8fbcc761db7c098e");
            when 2814820 => data <= (x"a93ff3c778577aed", x"3a998bf5eb93d176", x"84cf2e55a9bcbc3a", x"cf334c64ba0da905", x"dc93f3cdb1b563f8", x"effa3ba1d811db39", x"c854c4f417301273", x"8b65a8f93f3d89f6");
            when 7277486 => data <= (x"1460695e00874a29", x"60775bdab981564a", x"077e53e0a716e074", x"a111bcb2541df062", x"b851c629ea87d496", x"6e5c5d5cc99c9f94", x"c868508dbba73aac", x"25263dbb34d9ac78");
            when 23710455 => data <= (x"6bb702db3cc05acb", x"5ebbbdd7ae61c13d", x"890b4512a481fd8c", x"b280f6c816e5550a", x"5092fc7c53057414", x"158afa748ef3ac93", x"fc36053aa32461e0", x"9e9267478185d802");
            when 9848120 => data <= (x"b09f381dad4a29a2", x"612cb15957e64524", x"3e7096079971b8d5", x"33c39237c5808228", x"5e0310abaf1af1a2", x"f12fcc217b7438a3", x"f63a12955ec0f23f", x"1eea7595494d0f47");
            when 21913122 => data <= (x"be0b7a6d302b8806", x"d414f89402a352f4", x"7c72d1b9ccefee46", x"5442c671675f50cc", x"5c88e2cfff3a3c75", x"a26776deae6bf13a", x"369432b84f3d7c2f", x"f342f6d7a7801486");
            when 3477943 => data <= (x"ea8a5af94c9f61b3", x"0b771318a3b63d8a", x"28b02cd830a46760", x"553551b48192fa6d", x"5aad44ade912cf89", x"188f31f13cb00b22", x"1883266983f679b2", x"080f4dee68a7a1fb");
            when 33086646 => data <= (x"8a5e9e38924c6110", x"fd4ac9e581965203", x"85a298cd79faf9d9", x"f5757a0bdc8556a8", x"33cffeeacef84010", x"1a6720a6f861738a", x"b28984e240bcce7c", x"7c32baee212f03d7");
            when 2986945 => data <= (x"25f4e37f5edb5547", x"b7f73c04ce647443", x"2621e76c645ed7a3", x"2bb097e692973211", x"b819be344a14e300", x"d66d6b6677d94caa", x"edb523b5eaf32fc7", x"ed8f6cd1a48de5dd");
            when 10824917 => data <= (x"d8f843f5a324d40b", x"7807d01a7376a69e", x"a4a5ecde069483aa", x"7389cf87293c586e", x"5b7c431ea446cf74", x"b00918ab763fbeff", x"69bb54b8695fe550", x"31e6c8a4c5b156aa");
            when 32461926 => data <= (x"041ac790b322b9ca", x"dc0bb4c2c2525410", x"dec6b477625e0d27", x"d915fc9580f1ce92", x"f87c7337ebb41725", x"827bfa4f5ed39106", x"9ddabece748e6209", x"38c05bf2058bcdf5");
            when 8031963 => data <= (x"812d3692bade9d58", x"52cbf819fcf652b7", x"e635a10499bca91d", x"b3df6fe56961fb36", x"929ba96a7efa8358", x"1be80c210f7d85d5", x"a6c509cf8d9a7b42", x"358d7b1b280166df");
            when 12418587 => data <= (x"165690e50dd1ac65", x"65c77547b27a80f9", x"059002f9067744e4", x"0eca6af74590ee21", x"dcd8ffab89e4619a", x"2847799233708621", x"2f9c6dffc9a14058", x"99b07c9bf42cc3c1");
            when 12127972 => data <= (x"b7dde901c0afb8ee", x"e7e0988a3608d66c", x"642bcc411a8ddd1b", x"003cb363eda2b8fa", x"f2027fcbe70a233e", x"77cf9329bb3c9c3d", x"1eb74cc070c57f8a", x"605664a4001e44d0");
            when 11050254 => data <= (x"1e691b5f928c3102", x"22a29d05bad87442", x"ce299031e2975494", x"e712b648403bb6bb", x"c75fe63ae63d0073", x"d690c89bd3504fdc", x"90bf25b6ec4e6951", x"2c0f4a5f201d2097");
            when 31670503 => data <= (x"3eda45f2d5dc82d2", x"4c4947883f80aff9", x"2e299f6894f40014", x"c30f36b7f1585906", x"1d6f25e8dab0bd0c", x"b32eecc83f63e54a", x"79e7826c87534afc", x"2a161f89e8ef311b");
            when 31495307 => data <= (x"1c90fded9e6efee4", x"280547a43a509264", x"169b039a5646977e", x"67993f1ef0f735f0", x"5c066b614de44ea6", x"3cabbc08e7933b0a", x"dbd93d5009c98162", x"24fc15646d23fe06");
            when 21994150 => data <= (x"550b3f6d7bec7e58", x"8f60d73e7174106d", x"d603afff47655814", x"f982a3d04c604e32", x"0a35d0d27bd668b5", x"0ad7867156758c74", x"9b791b35b6ec9fc3", x"86a6c0621d8280a8");
            when 17703334 => data <= (x"6988c2f1681cd983", x"d8ad5f7f3c593c18", x"94d44090b003c974", x"de9cc1de173af89d", x"0ea3e35690bfb6cf", x"e1ea51c71257f0bc", x"ba14cc617a059cbc", x"087a1bbb2ec4c71d");
            when 6027672 => data <= (x"d3adda5775ca88e7", x"546a3f35cd918bfc", x"987c6467514d5342", x"0b881fff87e77eb7", x"9abe95b271cbb8fa", x"ab875d63a1dba64a", x"c8ab1c5d0971f595", x"4472db82504f74f2");
            when 16109079 => data <= (x"c950b9193fcbc489", x"562f05689cfbf95f", x"27a086a4b46845ff", x"a36f5c52ea5dc8db", x"e79a203dbc11ef8d", x"3572262e29c5cf2a", x"7970890f86875ae3", x"85b3ecc419f59ae1");
            when 3524873 => data <= (x"d0ea03879b5728f4", x"98a6c73ff015123c", x"01c370c9ce89632b", x"db08c1fbdac651ba", x"bef229380c349c20", x"f4a6ced57c9d03bb", x"73b392c83d3e2bbd", x"a7a210c4f42aa059");
            when 33056629 => data <= (x"5819171024994c58", x"bd0c91f59d600df2", x"875acf3e0d8a795c", x"e9c4e810395b8122", x"09dfb4a1957934eb", x"d0ade0649bf94b94", x"44e5149cf4916932", x"2f33419fa711f8e3");
            when 2709180 => data <= (x"8d0a4f212b6b1d7c", x"47af1c0ced07829d", x"d830f1fe94675c6c", x"caa3479f80143879", x"f4ac446bfb7d618a", x"17e1f33546d40d96", x"0137a301e22d23dc", x"d29523cb7361eeab");
            when 23601228 => data <= (x"56988cd1ec264ff1", x"102a250995c97d0f", x"5b7148528a327446", x"59462720e53120db", x"98c26deb80cbc3b0", x"14623afa0ce25310", x"4626a32f67460dd6", x"2d995e2b865f197d");
            when 13052447 => data <= (x"4f2db4e5ba5fe5a6", x"08d5609fc8144fd0", x"f9afc1173e276661", x"6b28d192eac2e591", x"98c56affeec77073", x"3379be48122c62fe", x"857a780b8c19c115", x"35653a16550e450e");
            when 5355509 => data <= (x"a421571eeb6edefd", x"a52d434b292b9f6f", x"a2ebaa4f7d426815", x"1ad888ce3c46cabd", x"c01d4441d9ed5265", x"e4cf8c808fbbecde", x"02d361ce5a250bf7", x"918f0c9036cd90ff");
            when 11708413 => data <= (x"86edc479ea1d573d", x"ca51dfe4c1419edc", x"874db5391b600dbc", x"6c6e0c7c92d43e51", x"11be64c6c6c8fe3e", x"c2920daf34a209a4", x"0be844bdde1060e8", x"ebfa58969da79452");
            when 15780896 => data <= (x"337fc27ea1b4b233", x"7fc6a2843d4ed559", x"60a6660dd48c23e6", x"3886cd88d23a822a", x"329cd83eaf553e25", x"cf18650684e76273", x"14b4d7c01f824fe5", x"74fd2690e0381be7");
            when 14838039 => data <= (x"244d3176aec63ad3", x"7d7f30fc4e750bfd", x"fe8d632fd3e77ad6", x"87a8999fb573e986", x"b012103f61a963f6", x"53baf63de74c9ad0", x"8676c1eb7519def9", x"b7d97c8b6ebb5640");
            when 24809937 => data <= (x"b8f41c67fb4a6904", x"dd4b847ac6b0778f", x"2bf0e1d4e1248920", x"e2eeeed218142282", x"1087e2c8dce26f5f", x"d28766e448b700d3", x"4b263c1829f886f8", x"357e906e8715599a");
            when 15007846 => data <= (x"4c2ae6da9bb1298a", x"ee85467a4938c635", x"0f196ec316eb07eb", x"f3f88a895dbff181", x"bcb4d7cba6941559", x"d55f4095772c4af9", x"3d02fdd908f15c3b", x"12c0e2c4674cb1e3");
            when 2464606 => data <= (x"f7b6c9c97c4ccbba", x"286d167b6f38ba91", x"efcedb5f8eabf23f", x"21647dc6a08a2d2d", x"be2bcd1bfce32400", x"45f909148da15b7e", x"4bf520d22b57f9c2", x"8908f56673e697b2");
            when 25492547 => data <= (x"e00e11010311f6b6", x"8df6434ed5dddd7b", x"5802faafa0e47df6", x"08aa48e9d47eaa41", x"37ea55e701613723", x"2a3f0814f7e31c99", x"cbdd5851f6b4b131", x"5939077a2a2b4ac4");
            when 29680546 => data <= (x"dd2f1b3f6aad40c6", x"ca07b3b1b51447bd", x"d5eb939dbe4ebfc9", x"c8f9e3dc11fc9a4c", x"4cf7d9c78eefa59d", x"e697030d02ec3c13", x"40257f8274b8334f", x"e16000548eecc5a9");
            when 1509812 => data <= (x"69cbae7a8af6392c", x"3a8a49ab57de00b6", x"1d1fada8a2ea7e39", x"f3251c9bef11131f", x"c3f97b324d60776b", x"a3e42e4ba5a99d1a", x"25b592ea5cff8682", x"bfd4a35c427fac9a");
            when 10464299 => data <= (x"3fff771921a958ff", x"2ca49c3a6e1990b3", x"a320e3c454e55912", x"63d8a41d0ff45c06", x"2047d702795bf31c", x"d635c981b4489159", x"e4885614e2a99e97", x"d0627ebe1a77e738");
            when 13512981 => data <= (x"a5278ed8a6db184b", x"0784793fde8a7080", x"7aa613ab2dac6dc2", x"c442ee1ea9f658ec", x"f968527e59454bc8", x"0a6e089adb3839f2", x"b2d52f41cd47b1d3", x"18dc03cc3f039f3f");
            when 15342055 => data <= (x"44e44d41e80dbb03", x"fb3a691d99432532", x"315c36d16e5fdefe", x"3792344256bb0ebe", x"e923d52932e7f090", x"1d0982f1044df774", x"0a538c4d6d744e1b", x"012d2a8d5b156d58");
            when 32662886 => data <= (x"327c918b71dd946c", x"5354964e1e22b102", x"470b59ae50491c37", x"2e53303ffb6d5820", x"f4f04b57762d51e5", x"5038b4190c1d3f39", x"6868b09c3d27811c", x"440bb50a49a8e854");
            when 24066080 => data <= (x"16e380c5521045fd", x"7f857b70e8e4cb68", x"5b19161d8c547bbd", x"cd4c1e01c024672d", x"4cf8933c7ae3e647", x"44170455873fb3b3", x"3c87291ef01afa59", x"872e2cd0cde6d950");
            when 7818097 => data <= (x"a7158f543fa16587", x"a59c276d274679f5", x"af07d39209fc5dfd", x"e5d5ea3e52ff0d17", x"741b4b9ea5948d5f", x"d2631520c1f8e4b2", x"fe91bb2ea9e7c4a0", x"4ad77a99a747f3d3");
            when 26795335 => data <= (x"1aa0f700c54fffcd", x"a0f974f2b127ff18", x"f7c2c2b7537a0eee", x"f91ecdfb082ee130", x"0bf072653cac357b", x"8b67c722d1bb175c", x"842bde81ef1b7e22", x"8156d393129f3c3c");
            when 26458939 => data <= (x"b112c7c84e5fe3f7", x"b031de4ee29c22a7", x"fcabd7de320ee3d6", x"4325823d7648fbf3", x"db263a1b1ab2e8ec", x"7bb4e9757710a273", x"3446c334322d9451", x"9532904d2b284deb");
            when 11540540 => data <= (x"3fb237369e5c8b45", x"3950c3f9cc133cfd", x"a3fbd2d9afcbe76c", x"c0d1bd9ed4180853", x"649c1274622e3523", x"f9dfbc261d933fa4", x"f3c24aca51488d42", x"68f45e0cafd1db4c");
            when 30374266 => data <= (x"214eac6947e05139", x"40c2181e8d9400d8", x"dcbe4cf1557f81b0", x"608f43478c65ad19", x"719e220bf24ed408", x"b1ce5067995958db", x"ee40a325c79a8b04", x"e3264aa7b5ac92ad");
            when 8163668 => data <= (x"6fb69bcbb6ab1d7e", x"57e3d734b9c0de6b", x"f5b0dddd605fd41a", x"eb2f394539c503f8", x"f0f859dc0d782f20", x"594964803e4b59af", x"93f847b06eff504b", x"867b29c5ad870473");
            when 15093008 => data <= (x"2190d2400d0684a4", x"302bb7911ba13d64", x"dfe4d2d0de92a8da", x"31929c60e15df6f0", x"615ef30e5cbaed44", x"55b4a443a8e873b3", x"6963f827c5cdf495", x"ee2fdae7e52b8c48");
            when 9784440 => data <= (x"7e487a729e597fb9", x"0de194b3065fb423", x"7114ddbd2ecd3302", x"61c886acfb0beb08", x"b35ec5053792a760", x"adea41cc544905bf", x"76d2e9b3d7927ece", x"fe05992249460ee4");
            when 29492923 => data <= (x"3a402220f70cda8a", x"a2185c06e846d818", x"b16770b541c1b3e7", x"c9b3fb44b9fd4d09", x"73360ab4fb593cae", x"63f580706a8d3eb0", x"21209c71b0238310", x"35c3af8b95e983de");
            when 22513857 => data <= (x"6605386cce7ad637", x"d9961d652ddc56c4", x"5d03bbde474f14a9", x"c7ac0c835798caaf", x"5c17b671ad3ca08a", x"8b7e658fe09836ae", x"d305ac46d68443f2", x"36a4197c400bc8b7");
            when 1503137 => data <= (x"e3c20b540fa87726", x"9334f8637abdef7e", x"2091dc9c524f0f2c", x"82f16a1fe0b90113", x"2d3ecc4048bce498", x"66cfa358722fafb0", x"54dc3cfd6d10cd76", x"8aa584e28aa0bda7");
            when 7420474 => data <= (x"b62a3a4dfeb9fe7e", x"daa5cbd6fdfb5988", x"c52f2507d0a74c22", x"9ffea044ca38f838", x"eeb992b2e68841c7", x"d7558b357eff973a", x"48510b811bff583b", x"612ebb91a00be8d9");
            when 5420178 => data <= (x"b7338db203f3db11", x"3c9b13874ef46573", x"5095992ffa5ce28b", x"df549b5b34041dbe", x"6cad48cc207f3c63", x"b5d664304f413917", x"affff79ec77e2800", x"e7e31339044f6778");
            when 10830794 => data <= (x"9045b6607125d901", x"d680ef116f56303d", x"eebdbfbaab55e997", x"00daeaf94acf1909", x"0651e172dde1ab60", x"13437ecb7c34921b", x"6c00bdb03cf5930d", x"c30a651c9631a443");
            when 11260533 => data <= (x"89b140b6d8e106d9", x"d656702a3efb60b0", x"a87935d383e8ef45", x"bbc5fff380f73587", x"5f710f8905015d42", x"8f8bfcfa987e3ce6", x"d09a2ba3630ee300", x"6ad28dcdc03d2ed7");
            when 27389956 => data <= (x"f03a993c93aa2df9", x"89b9c44f8864efcb", x"ab8e37dfdb7ec2fe", x"68b7d36ecc3ca98f", x"6523aaa8a669b591", x"9ce894627ec40b11", x"dcf7007d6f9689fb", x"1b11e89b372dcc33");
            when 11754395 => data <= (x"0480de307267cee0", x"e3e63ec0031aa52b", x"c00aa1629e8db61d", x"c6a58da6a31f2a2a", x"b6a781c9382b965e", x"19dc5e68e483f1e5", x"8093dcef458e143c", x"98b7314e78cc50e2");
            when 18769930 => data <= (x"91983d09b5596c05", x"22a8f60e30ed9718", x"f6dac5e3305d3b83", x"c84d6f939dfac689", x"840e2467e8cffd37", x"6b69a3f4b28db5c8", x"c87b96cebae3473e", x"074e07853ddbb9d7");
            when 30719528 => data <= (x"a461e6930f634d8e", x"3404297d048082f6", x"fded4514a5238193", x"1715567b69e60ae0", x"4b13fe94b9567186", x"4070a2721f7ff7a8", x"36e9795e3fbfac5c", x"8b153ca16005eec1");
            when 32366549 => data <= (x"48d108b576f29489", x"d27f62dd3ee2203a", x"4300bef1da5d3aaf", x"d63a4ddc73dc137c", x"aa8d3e9bcafdeac7", x"60d3567da4692d61", x"8255e849b888cdd6", x"00f41f50ee30fe18");
            when 22317792 => data <= (x"a6409147c9c2b1e5", x"0f192e5ad62e5e10", x"4fee7dc6c683bbea", x"88efc041a60d16a7", x"96daa405492ba8c3", x"e729b0abe0831853", x"2502e511e56a365f", x"f3d3cc8aeed2420d");
            when 8876986 => data <= (x"bfee1c0246d0ebd1", x"5b8131666ec7b093", x"df323256955a01fe", x"8c9440dc81fb3f1c", x"a14ec272f2539099", x"d5cf1adf8817f3ee", x"428b554b84364634", x"b34bacdfae6ad3b1");
            when 12885464 => data <= (x"1c90c0feba87b77a", x"828417019e1e1686", x"7920f45bf3ba9ebc", x"1b95280098ee9a48", x"c789f4fe84ae74de", x"3319d006f063b939", x"717bc777c3d636b4", x"3b6ab267b849ef4d");
            when 28197106 => data <= (x"9c861f02d282866e", x"133bf824053b5919", x"cd153585f48e9063", x"4e644af114c24c95", x"84f2fa6e5ecd372a", x"d503d2f02ec905ad", x"c820aa92ba1ea0c2", x"cca8bc318c9c339c");
            when 30006393 => data <= (x"87a727865bc91ffa", x"f3e79dc06bc36f97", x"d6effbc12010ea56", x"9e7a310f71bacc8d", x"125dfaf31bdfe8ce", x"439f9914a732e469", x"037be8410450870f", x"a486d8331422ce71");
            when 22849864 => data <= (x"fff0f3c5490707bb", x"d03e4c3aa68b1e35", x"1d3ab91d4d45aa8f", x"717ac939dd3fc370", x"1a30e50c57be3546", x"5b58b95fdc73f9c9", x"cf59e9f0dceea781", x"42aad30fb3910072");
            when 380701 => data <= (x"f3ad9518f255a991", x"59b02c10ec3412b3", x"1120a6ad3e45e2fa", x"08c1b2be1c281ce8", x"d65284269dab664a", x"41d1a7c9d6d2c588", x"77c7c4703041c62f", x"5b48bdee89a01b05");
            when 12965084 => data <= (x"44998aaef86f7e89", x"5fab8cdc923da79a", x"0c14043e396f06ec", x"a9bba6236bfb442f", x"99e0a76967c3e84d", x"355989346414a3ee", x"cb212f0b77348ac4", x"577138af12ecebe0");
            when 17274132 => data <= (x"59dfb6ddbc65ee3c", x"65848f750a66d1b8", x"94a27adf0ca81db4", x"096c63c4dfcd3bb6", x"ecbf4af01af587f6", x"4b6d569cae92204b", x"6cf7b1af9b60d07c", x"1c2ee00d1fb3dd93");
            when 17457198 => data <= (x"34606fca4781c76c", x"18a1fba70e5a66b6", x"102eb9d520819eab", x"ab10a85b98c65193", x"50a4f158aff25341", x"47db45dd3bd4b4f5", x"3d72d25bd8bf47e8", x"25118cc9ac97af23");
            when 33133589 => data <= (x"e3db1c6925ef2dd0", x"1c630669c0000bbb", x"d36f0f3893175d67", x"2595bba766384cfe", x"645f20f9c4c90363", x"c50d919606c17f2f", x"e94e7db91a6783a5", x"c873220433fe9f85");
            when 15180464 => data <= (x"ec88d967715b75d6", x"1f769060b252051b", x"aee43b839de4c161", x"3ec0410e71b839c2", x"7fb78bb656e418ab", x"bca1bb50d4ee107f", x"eed78d5c509a9423", x"8ffc2aa0c137e2ea");
            when 21473515 => data <= (x"c4c58be12563247c", x"19ca518d2c2f5c2e", x"faa853059db82775", x"25665e06803dc680", x"eb69f2f8e1c227da", x"05e3db47c4d5e782", x"a493a6a002edf107", x"ca08c8431804e5df");
            when 10296947 => data <= (x"5df435e1e6d7d1e0", x"b75018baf0484fc9", x"2716681b466d15e1", x"70579f11ea16ff27", x"b36197a087506d5e", x"7de9ed2fff41e56e", x"8a8c6ec6ee693f4f", x"45f19b0b3be65303");
            when 8774468 => data <= (x"e561c0700a2d52f2", x"1a8e31019f397d89", x"929c0a74a01ebe4e", x"71e935f90b1818ad", x"71ed588465940fcf", x"1602aa0595479075", x"807fb9a4b63e0db7", x"7b19f5ebb33d8328");
            when 21884349 => data <= (x"fdba121a568c4bde", x"cae8fb55a0b7cb1c", x"5fb4a05fee8c2222", x"6c9d449e2dc6bbe2", x"67701e70410f931e", x"1ded508648f36b93", x"7e818f34f2fd23a0", x"60982d440e1ca054");
            when 21211562 => data <= (x"d65af4c387448628", x"6608fbd236479c8c", x"d87575aaf88fb4b7", x"5dbaffc34871211a", x"ed35a069c030811a", x"843361bcd923ebef", x"8f9846f4cec9b238", x"245e9c4f941a2162");
            when 14462735 => data <= (x"d4cac642531b5058", x"c2aa621e35346fb3", x"c8832458f879bf8d", x"ddf92c300d9da264", x"c4ea806b9443aef0", x"dc0e2882cb328289", x"a9982c297add7bef", x"b84a93a3057a70fb");
            when 18063007 => data <= (x"63788cf60ac94559", x"b7c4f109ba0be994", x"cb0adf8d7cc34e42", x"a333dbba79a129d6", x"cf4aa46a2fc1363b", x"0ae4929b9c9f86a2", x"88ad3bce9befef1d", x"51c44a4cdbe654da");
            when 29974905 => data <= (x"e6b024df81fd5cad", x"8fdf62a4a09ca07a", x"7c695d3d8930115f", x"28c8c8db70948f15", x"e8b1d72ac90d3372", x"89e04565ce788f73", x"5ee5e385dd89dcc2", x"ab8f9d4f128feae9");
            when 23043935 => data <= (x"80854e4144f29d69", x"5489cf68a56ad4a2", x"fad2c624bf891ca8", x"ee314f87ad4b00a9", x"bbf766ebb6faa7ab", x"a7ad818dffe82c21", x"2b9064839fa06991", x"89df169a453f21b3");
            when 20541613 => data <= (x"7e0af5facbd6e14e", x"bafae6909c2de17f", x"402611975eb6ceee", x"6a1cc1887345f5d5", x"b294600b9a80a6c9", x"6435d047a40c66f7", x"68d1f6962b20efc4", x"1c86684b1eb05dfb");
            when 24080803 => data <= (x"6b8a44c9a665bc83", x"49c018c83929b96c", x"886646b3f570c9f6", x"b670275d450fdee9", x"424dc2b0e37efb23", x"11425fd9e57d8b7c", x"3f690d9654d35a8d", x"349db41ed55399e5");
            when 27142529 => data <= (x"72991d7f7418ca9c", x"7ba4cb85d0cce368", x"fbbbc265762f677d", x"7db1cceae0129e2b", x"07dedb0634d46d1c", x"1a6a679b4068d8d4", x"39025a19e4e1aa40", x"802405f1ce410740");
            when 13084149 => data <= (x"c3ebeb4c188bf21c", x"5c19ba129c6bd62d", x"58c30ab812d751e0", x"5606844132021013", x"84eacd5e36cc6f66", x"a8bd1f4c550a7c3d", x"bb659524695cdea0", x"96f9cf85c52d757b");
            when 8050128 => data <= (x"6358a8f580fa8e46", x"c9438da843ce4e4e", x"38af0e2d999f9c4b", x"bfa25c1030f352f1", x"b14c4234f0d4b028", x"ed849f7a0af78fa2", x"f840d8d32bae81e8", x"80736b4c4aaf15c0");
            when 25544257 => data <= (x"1bcec2beeab986f4", x"9ebd1509da365d6e", x"c665815cccda3c52", x"fd5e4b3922d01f36", x"c3501a7afbdf8682", x"230c1fb5fe7775a9", x"376cd6edd7ba931e", x"982b2a3e00407ca4");
            when 1633609 => data <= (x"a51dc02bd2438d6d", x"89d6cb53b8edf4ae", x"1a7f498a57d1ef31", x"2643ff3f5f7eb403", x"6ca1945a17a0d880", x"7fd4d79338d12280", x"30e03342b67ff0dc", x"434c9615353b2191");
            when 12847022 => data <= (x"8b0f00af72b365fd", x"83c74efbae440385", x"fc775f94dca6c7df", x"bcd4939762fb1484", x"553df427a3ad886d", x"895f76ec0219b167", x"cb7e76d246af4a93", x"9b48388725cb34ad");
            when 10553727 => data <= (x"4a74678e3d5d7b7f", x"2e8d04ce7de6f57b", x"e2a9d8bb4573c1d5", x"a5a93f205f94ea66", x"2024257d95fe2a9b", x"03db97aeaf272b62", x"0e462b67ef08db6c", x"5b5e974920fe014a");
            when 16108303 => data <= (x"c5a2fa458726eca1", x"c02e182fdb15c78e", x"3908463b44675c12", x"069d71daf6786c75", x"4e66294efe31ebee", x"048d76a6bb5a75ea", x"be92cbc64d59ab02", x"1b84e73b1b11aa54");
            when 15692467 => data <= (x"2da76d1cbf01919b", x"0dc736f47d644dfe", x"ca25791eccdf1ca7", x"40aa7a0da1ba30bb", x"ddec4d1d7d051c2f", x"009e4cff6b5330a7", x"f9cd804ef91f02ee", x"ea357916d060dc11");
            when 25622955 => data <= (x"f18ad96dc3c2f76b", x"fee5212cd5a694b9", x"ebcfc1ac8220c4e5", x"e6da744da53e6f77", x"7ab6f6ca063142b1", x"d96b164b6c6d8e69", x"c4c2ed4d524109fa", x"1c7620ea3bc6304a");
            when 27142765 => data <= (x"f4e051a5484f66fd", x"c803e9b75457d311", x"2c9c66bb7840bd05", x"624b4de3f285f37c", x"9a6d149a61477623", x"61a9d222158d7872", x"ca147e87e7d8837e", x"ee0716ea2a50bc95");
            when 25792107 => data <= (x"0e2926ad51a99ff5", x"75ed06dbe05289ef", x"335b64a827485a5d", x"04f460bbea20ab9d", x"a435a771d98d94a3", x"680d129640ca6b59", x"101eac00fa9fd444", x"0c11b1aeabaafc40");
            when 13724689 => data <= (x"eea12e6935cdc18f", x"03684717bfa93c71", x"dbdd0c7cea80ec84", x"aa988d2e4a8c6759", x"8880886c297e2301", x"94aa178b96047caa", x"8c2c111aebefa0f0", x"dc706d369ce16e6b");
            when 13531867 => data <= (x"74b83ef5ef817fdc", x"2ff60337cb9245c6", x"02c2afa9e0f9e67f", x"68366bf35547e0ff", x"3df73e995c75c2a8", x"57a7ece0f2728d9c", x"ad63e5c667cd8d2c", x"33cbde75e2cbc9d1");
            when 27777638 => data <= (x"eb5ca54cacadea95", x"5ffdbc513f704ae2", x"d4f734b8c0a07f95", x"efef5d83e026f605", x"a8342a2dc5d3976e", x"4ec0419328cc7790", x"9002f75784d6a8dc", x"37ee8f7def7a9d77");
            when 7959072 => data <= (x"010af2f8b4288666", x"f06b647267f35ef8", x"61d5308357bc5621", x"7c5c6a638e414f32", x"ab69e826eff70337", x"8a7e0cc307277eb3", x"dd62c591c43688ef", x"f0d060dea7e81b64");
            when 21164701 => data <= (x"da0f706bf67e3cd8", x"4fe5210f5a16c0b5", x"f826f316a0121e87", x"5d2f50e118aa9253", x"4f94902230660826", x"985353519eb1ac94", x"94c1534935902478", x"49dba4e2c8bc5bd5");
            when 23561323 => data <= (x"4dd18ea950bcc9ba", x"d23af83f6317ac66", x"45adbc9ba637fd39", x"a3c053e4f29894d3", x"5ab7bda85adb6de9", x"d6d076b3254cb9c3", x"53b0a16629827981", x"cab6398156cad1b9");
            when 22672355 => data <= (x"78a205bca4214b83", x"ad4f97211ca24e92", x"49bf3114a82eda38", x"b1173c6da64564b8", x"8efa92571acb73a0", x"df41ece3f5ea3c6c", x"068df4f656318741", x"8f3d4695e0042e85");
            when 8582956 => data <= (x"1958aa844f72ce48", x"b70bd2de5b41d884", x"65f04b8a14ed66ad", x"a9cab447efda2bd1", x"b98ace24c5764b80", x"a0f6cdec942815f1", x"138bfb023a865e4c", x"a0b5e53c04b161a0");
            when 30809594 => data <= (x"7148f703bc6e26ac", x"b71c900ff794444c", x"ba7a790bdaf1b22a", x"32fe5e797833367b", x"d27834c82c356e29", x"ccf6f5462bcb6547", x"122c8c8dac4ee36c", x"4d39ebbefbd5a833");
            when 4279125 => data <= (x"4c2f754102ce42e4", x"6b781c9e5fcf7cde", x"38504bc8416b8390", x"7497870ac87de970", x"a81fd6a686723c30", x"e1c693f882b8fec8", x"6901e8aa1ed4fcd3", x"1e2ba07f4a3fc636");
            when 1580773 => data <= (x"ac4f1c1883596cb3", x"2b43eb437856a4f3", x"890089a3ec353abe", x"41b01296e9ce9a9c", x"91f8f833a4548ac6", x"96ec9e37347d1f87", x"a9d313f60aee1454", x"90e2c289a481acf0");
            when 23986677 => data <= (x"84865e036d88ef28", x"57885de0429be82d", x"46855ce30f611ac1", x"55e7cf2ac613b1fa", x"3da7eac65b0e126e", x"06f023b4460770f7", x"15fa9798c8950b3c", x"e7b855c247115022");
            when 3086501 => data <= (x"4ae01e61185f6217", x"def91530d8067f45", x"d3aa0cf7196c2530", x"12156415e60f91b5", x"1b7cc1fa7a0f0dac", x"d1bcc1b9791d9498", x"f2d3eb61c18ee3e2", x"50d7b0cf34928b63");
            when 22930354 => data <= (x"0ae375bd27dae8f3", x"9bd86aa51aedf4ed", x"d387e7acdd0bfd92", x"7096a1850bff600e", x"1ded536a76b23961", x"5a545e8cb38820ba", x"e1cde228ee6e393b", x"4d63c59a4946844a");
            when 31651714 => data <= (x"ecc03387d74cd060", x"9a130f451c479122", x"10d212afa0de3346", x"360f2dc702ba1876", x"25c19f5b3e9aac8d", x"96df4016d4c99380", x"cf402e52a6091e81", x"f6fda45bc501455e");
            when 23147784 => data <= (x"8698c273f4493935", x"bbe493f0d659c2da", x"d3b3d403f6a5925b", x"a7bc3455479a6340", x"377d64ffa9c02e74", x"a76a1fac3b646970", x"b29d7a3191baedfe", x"5eefd15edb5acfa5");
            when 14366403 => data <= (x"93775f69ab8d2d4d", x"d96f9fe4f4c3b9f1", x"ad446e29a8a082b4", x"a7477a3638ef6501", x"0e1323a09f769190", x"d473753c3ff7da41", x"ab7712aa99b4f6a8", x"d5aa5c70d0a7ba34");
            when 18897984 => data <= (x"10b52fc33ce87946", x"e109a1e1e0b326b1", x"a5f13bc7b264357c", x"91abeb80c44674c6", x"90248f85a2a070da", x"0629f717e2521587", x"fd0f4fcf5b100341", x"577320d639a46304");
            when 21778576 => data <= (x"accdb011c84f56b3", x"a801a33d2b915ffd", x"3782af2e65b4ab1c", x"28b8c750d77d1091", x"3e0a8513a29e2958", x"f1caa1b1bf04e1f9", x"02ddbc0e4586eb42", x"bde645a7989ba743");
            when 21519817 => data <= (x"25d9be36339c9848", x"5e444ffb9f243a6b", x"ad773d7d49ce3625", x"47bb40dac203c95a", x"a9d0d3a5302bdccf", x"d03791da1f97b27a", x"dc67afc716e6321b", x"019a4ed2924ede1a");
            when 8969488 => data <= (x"6c875e884e4fbc27", x"42a7ccd8f68efa83", x"ebb3e5a817b386ea", x"57f4dd304ea97b6a", x"7d436903e3b1f524", x"a0358fcb57905421", x"7ae9ee17d741e55e", x"307a3352dc737a04");
            when 6449636 => data <= (x"d9ad6c5b09394934", x"ef3613165459f71d", x"4ca8bc84813a0583", x"0d2a88a6d1cc8374", x"54011808bce7b6f3", x"cee616b03497e326", x"f8a3db0c6dee1356", x"e36c05cbc3332d0b");
            when 1623714 => data <= (x"2ace89d6705bdfe6", x"ec45b6ce6f15586c", x"ace500df80b25b22", x"62e58195389b2f17", x"57ba2d626ccd48d4", x"40222a764f0cf9ae", x"b154c1b254f7fb9e", x"b872cb779c405636");
            when 16844173 => data <= (x"60f3b8cbb1e4973e", x"ed3887af60abcf0f", x"4776b7ea5c3ec064", x"3218fae72a4af19a", x"ef5720a0c8f16b71", x"a54a082fb3530671", x"82e25a5e5c935ee3", x"c0f6a504468a56f0");
            when 8677984 => data <= (x"ca4d15a68e0d707f", x"4f82ca47e6835ce6", x"c500cb9c098ee381", x"f5fee24cae302bf5", x"d960bdf07c1dd490", x"cc04e7554906b661", x"7f757402aefdd9ab", x"421533b76d367007");
            when 23762014 => data <= (x"47f8399e9c7c2ab6", x"477f562a80cd428e", x"6bb894d12d02382f", x"34f03c15502925f3", x"bb0d65d57170147c", x"61f8a61e667f0101", x"e0f7a82165232bc4", x"e8f585b0f0579498");
            when 11663234 => data <= (x"3d290a17b56e0949", x"def5ea2d02523705", x"8a455558af1eb5ce", x"a58993194a749906", x"a73954789956789e", x"21186751a6418fb1", x"e9eb0b46e4cf4d9d", x"9a0756d4ba17d8d1");
            when 19810728 => data <= (x"218aa57f603b8d59", x"c5bd000a5b12eea4", x"29fa400d48febdcb", x"3b9b337e1756f00e", x"89d79da5afc13bc5", x"0008691dfb903924", x"d69b4f5ac7efced9", x"05d0bf0a6b9bc64c");
            when 31230607 => data <= (x"ac8166963adeb2ad", x"d73cdbc0744aded2", x"a3882b12ddd51e27", x"451dfed24a0a2b0b", x"6d8baa45d48d9fcf", x"5dd5c673b14b4d8d", x"1f1e1a357479a054", x"d36ebd6da161ac2e");
            when 2853512 => data <= (x"4a025872e1b419b8", x"373d6c303a5e992f", x"1cad9758fcffedc6", x"73e28a404b76022f", x"198f06171a4b81a9", x"212e8c72ae4eb112", x"9f932ae52c3da5c3", x"e2924ac93edc603e");
            when 23440139 => data <= (x"15039296b66f94e1", x"faf44dedefabdfb2", x"4aa09c5c1f2fbbae", x"e06b7732ed7b0d99", x"31ab1128821224ff", x"7081343afd781bff", x"f6e3f1c6eb5ddd14", x"24ed1becbe177541");
            when 6440086 => data <= (x"a6110403a5d1618c", x"97ce34cc1023d265", x"8ce596abbb7337b8", x"71a2874bf58fa1ac", x"546dd6fd14c5cf38", x"c36819b2b9af5fc3", x"679f9ebb51b1d840", x"9eee83d5565ba72e");
            when 18352474 => data <= (x"e2ca1be6057551f4", x"1ecf93758043f2d8", x"0340843cacde97f6", x"3a224ef8828d0f88", x"b8a54f8ae79af788", x"8a811fd3f6aef278", x"7730d79e6b97147e", x"a790274c1175457d");
            when 30697777 => data <= (x"aa09ec70feb75899", x"9cbc0c21fa7c5b15", x"e192dd2381031b7c", x"644491d7c7e0b6fb", x"d4fdcda57797ce6b", x"960e758aa988daa9", x"8d9ff6dfcd26eef4", x"57f0074a97a60536");
            when 32453716 => data <= (x"bc658e25ba40804c", x"49b58d72a07c626c", x"872b7d76f85a11c8", x"c79a6ef5466c4700", x"40ce0125656db416", x"13d08b6f4dd61287", x"a8ab3369abf17110", x"fcd6c93fdae23249");
            when 15794013 => data <= (x"86d01bc8edfeaa94", x"5dc9ecd0a16ec184", x"5458caa084cc1c93", x"d9aa12f86b9c4386", x"8ab3b19a97fd8569", x"9ca0305d182fe08a", x"34602fbf109c4e3b", x"6b53fb831f6f6167");
            when 8622545 => data <= (x"15682f17efcf38ec", x"498b12efc98c7f94", x"2b65b3c910143472", x"add7a8cc1258ce00", x"ceb90e9aa77cc5aa", x"11d7455cb38434ed", x"126aa92b590f7ff1", x"cce30f9298a3e2cd");
            when 20484696 => data <= (x"37e12bd33c16337e", x"d1a371613d798512", x"a27e786a35d8d65a", x"fd89422eaa9af030", x"6823631a7dea46c4", x"56db274bd78eb67d", x"3d0496327942d4e2", x"9f82cdc8ae53149d");
            when 15485814 => data <= (x"0399c31bae451eed", x"f6c602484deb355a", x"0080a67858bda0fa", x"74602e063c752c48", x"d46b6f9ab19a4519", x"b38bcc6b8876e014", x"00cc4033ac33ac58", x"0765e9aaba1d0a75");
            when 1642084 => data <= (x"ee8df5a2a03fda55", x"6c8bb829c0375ab3", x"419856b2e2b13868", x"36d67d456c754be2", x"ab85d7d074c1946f", x"be8b0d4fb43dede4", x"806aee82d2df04fc", x"5fc9cf79e0d7dee2");
            when 1258736 => data <= (x"36511e86e69f0f74", x"b6261b05d3a26d26", x"946eabd63a5693e3", x"29cd704eae122686", x"ac75b289eca90512", x"eefb5d8ae5947e32", x"9a7940bf004aa611", x"a524a91f67a4a194");
            when 27883253 => data <= (x"729e4ff5bc167861", x"431fb6f81e93ba9e", x"e70c0f6a67811fa4", x"6f88a8ed54f83135", x"4b22e02c94d0be9b", x"48a9a844d22211d6", x"93d3c3b6f5924fd9", x"e797b4fb081b9ef0");
            when 19429530 => data <= (x"2ae56cd0e7235dd5", x"63c89d55adc65474", x"b20046b4756e3a77", x"ad5e20670722b172", x"e49f7bbfddfd367c", x"366f795d3a4de570", x"bf03f521c2682536", x"439aa39004d7a930");
            when 15015676 => data <= (x"36f025df89868c6a", x"4ff8af1e406b8517", x"58a563a617549877", x"34e4ac60c28be60c", x"0f502eec912f060b", x"bf22bc28fd39f8c2", x"654449d271646c0d", x"bd9cae778ca3c206");
            when 9467132 => data <= (x"6954622a688f5401", x"e2956de126f21d61", x"a0fd93f6db926e4f", x"b52541a88ecd70e2", x"e06bdce29046af88", x"1c885b13e62a2c8d", x"cfb8c79a044d83ca", x"58d5a459e1b57a02");
            when 19445868 => data <= (x"cf31e01898b3dbc4", x"5dda72d69270ae8d", x"5df9787e1cc6d8b0", x"10015fd2581f54d3", x"e4697d9265938644", x"4e8b466a4e4fd1d8", x"4b533f8128ec92b5", x"3c5515c6cc980d22");
            when 17380280 => data <= (x"3f5fa98852479d80", x"4507ed32f44bfd35", x"0ea47dade2701913", x"6461fb5c5c2c23f9", x"b2bcfa68c8b92133", x"cbbbbd8e7a4097c2", x"ded02a38afee1363", x"8cb02575578a2193");
            when 7536590 => data <= (x"9f5a568c7d892686", x"11d97c4fb5a5aa23", x"3d5cbed8d6b7acc1", x"cf637f12b93f266c", x"ce1cf78767c04f6e", x"74a1ac7239c00872", x"756f8931625b3f60", x"b4da620154b79a06");
            when 19089100 => data <= (x"6919752ac11db382", x"1441f170ea65a87b", x"3ceaf5d8883bc4d7", x"5590996f7cc258b9", x"531ae415b96ed5df", x"89659f968221831d", x"ae2d2966a4c30fd6", x"1b3597cc033d643f");
            when 1532392 => data <= (x"df843dbffe96f792", x"8d53fa7c871d6e77", x"e82229c586e9c806", x"4a28bafd20acce0c", x"1131ee3dcbc42a28", x"3e264e45c60f4dbf", x"685824b81fc02542", x"98d816025c053113");
            when 29389235 => data <= (x"4825a959d1223656", x"a3adad3c5ef5d1a6", x"bb93924be6607386", x"81ee93e45b578080", x"ab5f4a4394179b0d", x"b5717df9e6c65f1e", x"734478b03fe3bd53", x"670c6d853f269923");
            when 11566879 => data <= (x"c31073c36bba4624", x"428373925b4d987d", x"97c359a06b384e2f", x"32ed3bdba2589bff", x"d0f359dd88d2251d", x"09721dba8ffa66ad", x"64b06714356e5ddf", x"4a016b59799e856c");
            when 1713958 => data <= (x"2372aa9591754cdb", x"c10251f58de47245", x"7316f73934baee5b", x"4435b5051ef7d212", x"6e61365cb46ee6db", x"998dd3f468e01efb", x"7b2851e70b596ee9", x"e2b9581cdcbab329");
            when 11152281 => data <= (x"da1ecdfad5938020", x"6908638b0c37d96c", x"c319738fae4de378", x"beaf45c505aed063", x"821a2b69adbc7839", x"1d07819741b98658", x"3886caafd8fa40d4", x"51f79ff0009c320d");
            when 26555335 => data <= (x"10614488476c2ade", x"627f2e7a62abf765", x"1927e9b12f56c442", x"bbc745c384108dc8", x"822d7324fec9dd3d", x"264d9e238dcf414a", x"d66ab125a4be718c", x"7328b234247fe2f0");
            when 1402285 => data <= (x"a2a096704b31377d", x"71a8cde618781246", x"40b2c7a485a1bfc3", x"a58279cc1726f9d5", x"8738968dd2c1090d", x"d581b6a23ede99ef", x"ef948fcca52d9604", x"f23e3e3c34a764b8");
            when 24731011 => data <= (x"5a21d86203ae918d", x"e1124ab1cd4555ed", x"5a73f53a94c7478d", x"cc140d69cc31cc78", x"c58637e83f2da335", x"3b14a22c550d9173", x"66d6263f6d50d25e", x"44dcfda81dd7f656");
            when 5482995 => data <= (x"8d2ac2dab437e5ac", x"a2b2a4d3b0e413bd", x"37d16b958c7940cd", x"db867831cac8c106", x"92df52d7891f81c2", x"51f4cde214238584", x"c90825023e1aa689", x"1bac37a4ca7f3aba");
            when 2231133 => data <= (x"734b51e02fc8f533", x"88005f451a8979f2", x"fb4a84564a35af4a", x"4389f3f6a3accf84", x"f5bd65b3eef3c232", x"167c10bf6e65d012", x"42d5f8b1ccc56648", x"5d37687eab34d466");
            when 17960046 => data <= (x"9207ab099b977cd0", x"c5c1421e6d1678e1", x"2343d9544253cdc7", x"a2133b9282f7e8a9", x"5d6a0a015974fc98", x"41d86fe627e72101", x"53a6a082a172cc65", x"186baac734ef8b50");
            when 33103735 => data <= (x"0349c2900d558791", x"9d042b110d322f0f", x"f2edbd60be63ffa0", x"74b4de88d2323162", x"6387afc40e2b290b", x"912c969a354aa867", x"4692320b471a3794", x"8c1fc921b088e429");
            when 18897401 => data <= (x"a2673b40427df364", x"8f091ba76fc7c1e1", x"987c0558273e0a9e", x"3ffff781c5ea527f", x"0eafef023dfa4d68", x"5e9ffe3313e6e96f", x"9dfc6810563a67b4", x"795c865c34488916");
            when 5581254 => data <= (x"23b8c30208bda237", x"0a6e5ff07ade3e5f", x"93bd415aaf1a8817", x"dac71094681a0428", x"435a29e1d57548e5", x"bbf4a1c15e61844c", x"a55b8396b5ba5045", x"3183e6e4a52ce95b");
            when 30376490 => data <= (x"48207b30b1bb008c", x"f199014e12ab1bd9", x"40701ad7d843bc49", x"c16d7a304a31005c", x"db5c686a080fb6d2", x"498a9c54adbf7e62", x"a74c59403237e05b", x"53e9b2ae2c9623e2");
            when 23888178 => data <= (x"1da0ad6bcd2e0e69", x"4b70fd3b703b454b", x"2f57bfc828c74d50", x"dfe270ab96348f09", x"53e00185672fcfb7", x"2778da804e0036d0", x"75e5237255cc8c20", x"eaee916f05f26b65");
            when 33795030 => data <= (x"255804cfa68f2110", x"1d412dfa68d8a6d6", x"4ec890c139acd933", x"4aadcc23ea296b9b", x"b20782120b82919e", x"bae081d856926da4", x"aa6eb6e66e38e22c", x"a3e3da1cde8b32ab");
            when 19141863 => data <= (x"7f9db5047d83e5a9", x"4b2f772820d21fc6", x"3377a69e89cc5988", x"646a92914a3f8af3", x"e728b54584407463", x"8a4b8f316cac0624", x"d6eb53bf84aadab6", x"d6b2b76cd445158a");
            when 593573 => data <= (x"55189464895785d7", x"bf211d35d698fed0", x"22d9af4d239735cf", x"5ff22390dc8ecf1d", x"392fb5228c719818", x"9352e4c0b42cdb82", x"ee1432df2191b050", x"decf5563b7ba4a6f");
            when 13480776 => data <= (x"108a1fe2176d0d96", x"a15c61781bb157d4", x"213724c4f2b670d7", x"8d00a655129ddb66", x"ee08a8ad824a4021", x"055f6a7eb04e3a5e", x"a3c5b2c2fe7a994a", x"7166e4bf8fe151f0");
            when 13975455 => data <= (x"595276726c1b2db6", x"eed7d83a6c1f8707", x"de7d7a6baf1a5005", x"887e163d56822ecd", x"690c730284fd39da", x"c9425bbd5148dffb", x"e92fc446ea139006", x"dfe5ae609d041ce0");
            when 1883941 => data <= (x"c479d80da82a2b41", x"b97ae106fa326e51", x"58586fd31beacecd", x"d9ef13591ccda1a1", x"a4d83bc7083ec355", x"ebfeef09459eb7cd", x"736a01933b565c22", x"3c4a5b46640ea601");
            when 25993780 => data <= (x"f068737adcdfa988", x"fb6faa966c32acb1", x"25dc4e5355d12a52", x"031407765797031e", x"031bd604c4d775b2", x"296aacee47246436", x"5d33a3d7e5e22faf", x"1500dd6299ad49ec");
            when 21562958 => data <= (x"13dded014c9c6683", x"ce621e60b67f5388", x"a519cf0072c877ce", x"291e9ed76720736d", x"029032d12eafa6a8", x"c728a5dd1cc70d65", x"e38b5bc65b3a2085", x"f0d1ad526ccae38b");
            when 7254108 => data <= (x"91a18cf6e715c04e", x"54e59aeace7e3483", x"9284c79ddc864b67", x"edd22cce5d4b4cb2", x"ad8b9ef0c5c445f7", x"c1f2208ff08651a9", x"f7569275423a267c", x"7ad7af32792b8e5c");
            when 28390719 => data <= (x"e1aa9fc5bef883e0", x"5d4b1d31ab4b157d", x"48357c9d08ae0276", x"e7a6a60f38242b01", x"034e57a36038c399", x"bd864210645a0fe2", x"6d03030d6486ece6", x"e3d80849c1cb0564");
            when 24877755 => data <= (x"91c5400dca2646ce", x"c26693a6786f5bae", x"68d619b6e7695fac", x"5139fa102a83dd94", x"ba6feb23b88f4a40", x"3fe8ec2f4f1a213a", x"c6a9392ed37af7b1", x"9bedf0b698b07a95");
            when 7032467 => data <= (x"97f29c2872ed01a6", x"d9ecb027b86d0718", x"d04c41003c0ed0b8", x"f1b0627ced1d6099", x"5075a1f2be95a606", x"93c9d46d9b1e6ef6", x"b1ea0fdf866c2d27", x"da7c75ebf990dcba");
            when 7396038 => data <= (x"20cdbee47f002c48", x"9abb1977c2b01e85", x"58b3a3134fa15922", x"85a708540c6ac5c4", x"1169ed467b009146", x"989e509a933252ca", x"62f8b5a6432ebdc0", x"15deb6e44adea4df");
            when 31000530 => data <= (x"d5e687225d82bf4a", x"188243491540651f", x"078f6df3cea4c4ad", x"5d0a4066822629f4", x"b1d4c367d4bed574", x"46db601a2f8d971b", x"1298fc13313ef1f7", x"79b8187d03aad0a1");
            when 15681809 => data <= (x"dbdf9ff56563066a", x"6ec24ea4f697c368", x"aa8a9447852bfc40", x"88b0a0c94aa369f4", x"f00cb4b3de7eb45d", x"81bfbe2898f345b1", x"b996185bc37091bb", x"d36dc37c0c2ce17e");
            when 965875 => data <= (x"34fbae909350e90a", x"7ad4dbff73381ff8", x"b4caf3062dc8943f", x"8175d62331c5b2fa", x"6ac8430950eb7ae1", x"888df4b64dfbe84c", x"843cc76c7082d51e", x"c8ef2c492b054716");
            when 22389474 => data <= (x"ddf8ab5617dec1e9", x"23053ee55cda8f03", x"56d9ad128e687545", x"ce3f6e500d02b45f", x"2fb82c2861fd6683", x"ab8f3f5a124d379e", x"0cc9abc7ba52c669", x"5b3269a6d0012817");
            when 32981210 => data <= (x"b33fd4f32458c5d6", x"1b608ded792d6340", x"ddd7c5f80388daee", x"b21d35d212f72a05", x"c3588d0417b796f3", x"7f8b63f9de6d8164", x"7092c2303544c058", x"3f9a55bb5d0b8340");
            when 31533996 => data <= (x"f0e7113a8972b3b6", x"9d74449678f9ff40", x"58b87bbaf2ce9fb7", x"061c744b7c03d9c3", x"a581f023490032c3", x"a30621214c61b9f7", x"49e9025060d2ac19", x"f06fdf72c54d6166");
            when 14797160 => data <= (x"ee095fc4eb4e1f9a", x"5a4b82480036a3be", x"a5a815ec7b414491", x"0f7a534ab34a514a", x"b40f5e4c0551b028", x"3f868decba632068", x"b8f83c0fd63b4780", x"f66b8d058deb4467");
            when 16948955 => data <= (x"51e7ab3d8e584954", x"da8da06db0fb90c6", x"a3fd4f5d75773f60", x"1fbc459072c4634a", x"d332adabe2d19e34", x"acc11ae04f8c6431", x"f66bc33d9e50631d", x"5f2aad84aea7985b");
            when 28571207 => data <= (x"59dbad4090bda38c", x"b03cb58a6dbbf08d", x"cf79e3cf1b16ea84", x"0f5bcc19d6a2b93d", x"9b3fb579a767afe6", x"b2c2044433d15884", x"22e5a6b6c5c33e7f", x"a2f2d7585fb68893");
            when 24658471 => data <= (x"98c2c2628ae4014c", x"5339e82ab02ad4e6", x"878850fc5a5d6932", x"669c979929acc6a3", x"6e8510badbc2e578", x"8af44d9ea44d19d5", x"2d5948292b211076", x"4301720cd8683eae");
            when 25619054 => data <= (x"5e3ae4a5cb283b26", x"acf8b92912744f52", x"723119115b2afbe2", x"9c3eb669f34f759c", x"4a0cb830bb0fd394", x"b91f97f6695adc66", x"408e536eb9150437", x"8b1749b5abf1dfde");
            when 12466215 => data <= (x"7d628e2c412922d3", x"e92d0b218591ebab", x"363263c6850df56c", x"f6c39cb9d7a41998", x"809a4d552348f4bc", x"a4ad34517f567b9c", x"f290a04b27d38ae5", x"6e0d383cce426e89");
            when 9720834 => data <= (x"2473bf9dfe7943aa", x"97ecd4dd76fa5afb", x"c6398be1ac6cd3c0", x"45a0493ec8d54420", x"296f6963f0dfcfa5", x"c095132ea6af3414", x"d32113a964e8d766", x"5517493bb559ff1e");
            when 10861763 => data <= (x"34221d0714bca394", x"0a5e80985ca6ea34", x"1cfe5f843ee5e207", x"02cd6bdb5542faea", x"fac642eea2b48310", x"8529ee702b133dfe", x"5cfc5e8a303827e1", x"9aceebf4556a0ff5");
            when 23762377 => data <= (x"392a420965f01052", x"61e99cded91e6413", x"9d741b96fd96db1c", x"f174fa0498990ee6", x"12524fc2fae013a3", x"97c6c023fa4adade", x"3863380ca0df3460", x"a3d3da31231d0086");
            when 32735766 => data <= (x"11829f8df4a0fee1", x"4026b52737d1110a", x"bcb68a09cf85e75a", x"8d8d9c556c883f7c", x"bc06ab334a16aa9d", x"7ac9fd6e03422782", x"f0fb4de0020544d3", x"e5fc6d9da19b9fa3");
            when 2990278 => data <= (x"7c4c63ce448c22af", x"936d47f6c184e5a4", x"820417f56ca117ec", x"7d436e39ca5d582f", x"4ace36c6165b2c7f", x"da9c8a83c8c7e56d", x"ecc2953ca6b30be3", x"4e4f584cd6bbdaf6");
            when 8979951 => data <= (x"84e012071c16a073", x"bba36305aa3766e6", x"3ab9fcb12d0d8a25", x"0add499fba2f981b", x"cfe01b1c047eaff9", x"407b4264ce4c80d1", x"796325948cebd6ca", x"ea82f353fe48cd79");
            when 13376800 => data <= (x"714fe4d244111233", x"443a35d153b8b2b4", x"ad86d58880599be0", x"af41fa969fdf621b", x"f017f19318318bf3", x"0c8db9ab47daeef2", x"8cf167f4d93bc2fc", x"74df0e6b7661ed93");
            when 13011446 => data <= (x"e360245fb846d941", x"31135ea9f50d6883", x"3822fc2e736e0c1c", x"5a249bc0cbee837e", x"97bee77ddb75c606", x"3ddbcac805d11674", x"a35bd9d69a6405ec", x"d1cd5d4ed44c521e");
            when 11278682 => data <= (x"6918e0f4d7d3e7a6", x"ff7245d77f9bf2ca", x"05466b444d93b458", x"4c2aabe53acd71ac", x"bbc3b744b264396a", x"9e01a6b8e3f844de", x"60d7d1c94fd74242", x"9d4a022cf65f8b46");
            when 32617718 => data <= (x"be2a5719ea50181a", x"a7a51ac7a9eb758e", x"0d60e2281f6f130d", x"a1c31f55ed614dee", x"7c0edcd7c5a3e095", x"326d1047c9bce01c", x"728b2b9f0e5b233d", x"e04af87f0d650fdc");
            when 2370047 => data <= (x"f719708652ba0ebe", x"ed88cc42cf6fe850", x"06bd44be8afd1258", x"4f844b9ff4af0a67", x"a0d8bb7104550955", x"399f04d3c5f410f8", x"a8ea6b4f709a4052", x"6a5c15a0bb56d16d");
            when 22105540 => data <= (x"a77476007a642727", x"665e4316b862b773", x"e12685b9d33524e4", x"58bf6919ad66f932", x"dd0ee6b310a48885", x"0d9672e279b8db56", x"eb39d6206b217d26", x"2433db21c720ec33");
            when 24902578 => data <= (x"28de6b46aa9ddf78", x"78b70c0649b28754", x"bca311f2f312560c", x"d62f00d35d198c9a", x"1d55fbfa59d7c278", x"0616491fec802f0a", x"60da44626b701674", x"502942819732c780");
            when 33749715 => data <= (x"fd09e4039fb1a9c7", x"3a1123428f2109d9", x"776f94c68698b018", x"1d356a490ace2053", x"8a474a021e3d04b7", x"a171aed342329da6", x"6c0a9cb5a0018da5", x"6a1d7a8db8908e09");
            when 6456743 => data <= (x"da504f52f3aa7df0", x"8f28db0944a49fcd", x"83392453a66069b8", x"b3c464c1c9e0ec23", x"9a8df72bb52b01dd", x"2264637744e19d55", x"fd0d05c462aa17c8", x"96d3319b540782b3");
            when 14461361 => data <= (x"b8f2ff166e072d54", x"331bb72798242392", x"372e747ce3e31e3a", x"95b4015b8d382aef", x"ef4922cbb7975b23", x"c5cc9b80bdf99919", x"9e9194ce91e2c144", x"f63c403251a5ac68");
            when 22412873 => data <= (x"52adf37949de639b", x"af657399d0384cda", x"9ffab9b800e46a87", x"c685385be97c840c", x"c32bd56ce6f75464", x"c1086c3dec11847a", x"790c2f3c072844ac", x"34e74e570b3b75d7");
            when 788608 => data <= (x"0df3df7f7eac3730", x"5b74c6b57bf230e2", x"60983eb982b107e3", x"0a04520fa7dd0da7", x"d2efa927f7e917f1", x"915a72a72233aa58", x"d20f9427a7a5b3f7", x"863d807c5f2ea6b3");
            when 8142855 => data <= (x"d7fb9c08ca7504fe", x"fcd33cf318922f34", x"6ff92a2701c54be8", x"850ebd3b24f264c0", x"7a8db2a02f241414", x"09e8220ce48fb056", x"cc3f76cc752db7f1", x"ba3f2b3ef37e0751");
            when 28049894 => data <= (x"eb3a058689b9acdd", x"0f8701f2125b4cef", x"61376ef67f891e1b", x"eb8d68d63f42f99e", x"704f33d187a02fb2", x"bf68f66adc517867", x"aec3343394ce9b2f", x"acc162cf4fe51709");
            when 5786842 => data <= (x"7e53e0d78f80f94f", x"3ac9a3368b50acf4", x"af78839c50db63eb", x"f1a1aa95b46cde53", x"c761edc0ccc7b297", x"291efb6b2d6dc4c4", x"adeec415ecb1f2df", x"a7b9196c8623fcec");
            when 25294767 => data <= (x"60defdef8def002a", x"d257c74a506c2562", x"68ab0bdc295c4ed0", x"e49ed41392446d7f", x"b5b81aa2b479412f", x"f089027b18148061", x"bc988ae2b9fd7710", x"35f460ec167db709");
            when 33412821 => data <= (x"50bd41b588902000", x"f7601dab29360b1f", x"8fe1e339ed1d818c", x"60315187e87db350", x"67444b3b5141b8f9", x"6da376b55f13f088", x"9dcb3815eca904ca", x"6cbefd059131e343");
            when 22920222 => data <= (x"887e0040bae3256f", x"78000019127ac704", x"82f6d201c601bbc7", x"5a16aeecaf4e0867", x"0fbb778ccd095c18", x"cd93c05b140a7f2f", x"56f957d7cf72f046", x"fdbd60deaf4c33f2");
            when 5513809 => data <= (x"d61ce085f57451a0", x"2e29b3a63bb976ba", x"483e4dc4a12e154b", x"7c23afd905e78f02", x"f95516ff91de6846", x"eb68a453a7b97830", x"ca61802f17f3fe5d", x"ab7e1b493ab85d4b");
            when 24020307 => data <= (x"2cc001452ea01856", x"aca2c170f5272e5f", x"6113551ad39adde7", x"d7817aa0ed5175a9", x"a38099cfab66abde", x"e70eb2b1dafdf87f", x"e6898836b467c539", x"73050121d7bad699");
            when 16983481 => data <= (x"0c348a82c82fb412", x"ae14f4245c1649b5", x"51764491ba5e4042", x"1c1cbfb27dc21b0f", x"0eff1b6e4db943d5", x"a18ffd00c5d42818", x"34e8872efbdec307", x"5c8f41e0aaedfa58");
            when 27453210 => data <= (x"39ba90351ca732a7", x"abe43dc42b3d3d07", x"1f17204d6b3a7cc8", x"f0468d50ee27a7b0", x"23c28527f3e20563", x"e21ce1b804acb9c9", x"380f8a2af94ee98e", x"15e3303f19241531");
            when 23047835 => data <= (x"b0cdcb414c2cdf29", x"595336baf7be716c", x"db8173ab72835830", x"07bd9ec96dfe3186", x"6fe06bb0747d9201", x"f0f0e075221be6d1", x"27dcaeab2233fc3c", x"9ef9068cbf06cc5e");
            when 28750264 => data <= (x"54546f4208525b9c", x"5912b682ee4ed144", x"64fb4ccde1ef23fb", x"c358c5996af7984a", x"26c94859e8215d3d", x"77e54cbe39ad670f", x"a04606ff7f103870", x"1e570931a83f6316");
            when 12222283 => data <= (x"9d67e382ba61a5fa", x"304c324ede7517d0", x"e05b2ef2e50e4631", x"5b3593182821f8c7", x"dbc7b8b71ff6332d", x"ab9afe2cba9f8cba", x"7255d4b1851600cf", x"dcacabf1622974d8");
            when 22812503 => data <= (x"c6c206aa38c72461", x"76010cbcb872631c", x"b9dae779473bdc03", x"d246eb2d0afd1e94", x"84ab32509e56452b", x"dea8b5e2cb125e0d", x"b4823688615719ff", x"aee19bfdaba3b7cf");
            when 19314430 => data <= (x"88b7d14cc7b0a529", x"b3d8e5be0c983e76", x"33c5468102610029", x"2b38f173f834367d", x"dee353ae7e2c970c", x"db56a92e5ea19365", x"c20bce882d383ec9", x"e17d1721e9ed0054");
            when 17278182 => data <= (x"8b378a463880dcad", x"da5f97b1276dad27", x"5d77f53b356eea36", x"78d5fd21ab2e9031", x"fcbcfb49f4de3a16", x"413b375e6584dec9", x"156d81d04f9a8cfd", x"ac342604f743c98a");
            when 28650002 => data <= (x"85fa2b7362a44d17", x"5232312362b14b5a", x"577c8b36e93e6eea", x"0a6dc8cfc0d28e34", x"8ac938c3e52d5fba", x"de5787039568c71d", x"05f4b512af35d3c9", x"5ddf94adb4d274cd");
            when 30941521 => data <= (x"9e709150467dfa56", x"b37eb97adbcd4027", x"7e740da5214bbfa7", x"587f880743554079", x"d6bb3ff478e8583c", x"cb54daa201af175a", x"11175ad52ad730de", x"50bfd114694d7765");
            when 4666733 => data <= (x"2766a63a11c1671c", x"b1f9facf80d4c621", x"4235d6fa52636e04", x"3b79ae89a048a8ef", x"130be7bc1ace54f1", x"eb86f048021988c5", x"b683886986423a40", x"27ff85e99a7425b1");
            when 24905681 => data <= (x"b77d7a4cb82c0a26", x"7d7c3fc272e0b8e0", x"477341c7daada3cf", x"0711baa87bd8c552", x"969109b8921355aa", x"8baea34e33653469", x"84b7143e661320ec", x"67fa559e7f530b8a");
            when 2338168 => data <= (x"52c270aeb11154c0", x"e559044666ccae23", x"03043d9901db5e04", x"56cde00b0304e71e", x"b478a16dea76d05d", x"38ef1787128a004d", x"0f7120f0d3e14f6d", x"fcb37a4aab3be0c7");
            when 24446586 => data <= (x"f85774a7c1e364f4", x"030a91ce3102b05c", x"9225a9f107f14927", x"ee36695be80a60e0", x"2888a6c95cb4ecd0", x"d04874663ac82d4e", x"767750b0a2f1c019", x"7dfa6b3f46e72d7f");
            when 29662885 => data <= (x"70d53d56c580ffb3", x"275865e19f6858bf", x"821906ada1e4b272", x"7a58d7acd9db4c0d", x"37d345054e921516", x"b2b73ee2ce0586cf", x"5ab1a7a74eb01923", x"0336291ddcdc7620");
            when 14263162 => data <= (x"a56500378ca76267", x"b3a792d8881f0708", x"ec5b0704648b4468", x"e5ac64de0b552060", x"a62ecef82c24de17", x"d1d3d1c97a50b788", x"1a43129e91dc4ca0", x"e64698d355d84723");
            when 33487203 => data <= (x"a4299414bda6c811", x"30fa5849a47dc9c2", x"3e5068c68a554b95", x"02fa91261dd13120", x"70202eb859c3a8fe", x"872e5081941a47a1", x"dd226f5ca42c0dee", x"a5ff380094075f23");
            when 14237608 => data <= (x"5f6b1e0fb824e107", x"e26bfe4bccf1efbc", x"6c5ec60028b90856", x"44c98b3421fbec04", x"50ec050bce1250a7", x"b1728781aaec9c93", x"f25a601b19ac3bcb", x"53da54cfef4df9dc");
            when 16791927 => data <= (x"d5f8d9647f3973c3", x"ca58b987b5e60a0c", x"b852c97aedb40725", x"5dc8337bdd69b6a1", x"a4fa5ba0701fc6a7", x"3ed2d00148161ae4", x"016e457b41918404", x"e0e320b0c5f34b19");
            when 11619768 => data <= (x"c1f018a9ddc8d04d", x"78bfc38690f533c9", x"b68b22b49c550fc3", x"aa18b4137ca5c14d", x"609038e9169638d8", x"b6b8d51a13d5b1b5", x"c1555072c5735063", x"95b409d7bae453cb");
            when 21520915 => data <= (x"4ee95fc79260a7cf", x"5f74f560588f3b45", x"8e9d19a00c5b5d40", x"d92f030b0a2bf4a5", x"ac1ca886903bae68", x"3ae4cebcf5973bfc", x"ac0c0579b1d182fe", x"2dc7b8d630ddf47f");
            when 4435314 => data <= (x"3a60422573a1edf0", x"eacea8e271046cf1", x"3c49464e0265f0b5", x"964ca3a287f248ab", x"926a60100a305788", x"90b54f34ebe6c57a", x"7c8240e4a66a35e0", x"83fd4a29c7c23da8");
            when 29053565 => data <= (x"6f03d8bc2724c5fe", x"22731d05bb4aee4b", x"0f5ea5e9c40cb2c4", x"2041149391bb5c9b", x"466f707115b7caaa", x"61130cab67de00cf", x"c1e0aade28ba74ff", x"789472b56eb280a6");
            when 4643962 => data <= (x"5146643c65a56919", x"6a7227ca31dc0765", x"9e527d64dc802479", x"d8805b1c5ca7482e", x"13c81093f08785bc", x"590fc09653c31ad8", x"f5ca313435846356", x"28d35ed16cd64b55");
            when 33078119 => data <= (x"31b97d95a3b89551", x"f205b50870b6c687", x"2c3858e2e7c3244e", x"62116fab9a77cb3f", x"49ffe0c66d70f289", x"7c55f7d6402142cd", x"49aa639220adc9a7", x"708fa5d0a2527a24");
            when 33695411 => data <= (x"c7137aec50ed50f8", x"4e1a02ef8392f71f", x"86d526b35dfa60b2", x"8d305d7c11a2084e", x"7293d0cb11176744", x"d40fa7ebb37fa30f", x"2196e1e460190437", x"0a4a869083df2fb0");
            when 25304908 => data <= (x"af333d07f2f0f232", x"c04aece1dabe686d", x"ae23c68d3f82807e", x"d7299646c1eeb027", x"1ad260c28db11edf", x"3f07be9cf992dd28", x"8cd2ec4cbb2b30f4", x"f5577fce0b349a5c");
            when 10501049 => data <= (x"bb8e0f3a74940a8c", x"713f00fa9c627495", x"cf1b41d090dea2a6", x"a2f37d787a53c5e1", x"0139dd28d720d5ee", x"ba8b75661cc286c8", x"918e64847342bb59", x"117b94ea6014079f");
            when 31072871 => data <= (x"269cde40b03a231d", x"e11c87bec00616f4", x"38fdc36b2df94fe1", x"7ee914ecfbd0a132", x"eae423f28533f8cc", x"cac7141f722a8365", x"74866ef22eb01dce", x"9f9732cf57f5432f");
            when 1648829 => data <= (x"de39ffcaaead749a", x"d95dc3033c794d4b", x"5021196923fa1452", x"87d0bb65eb836d80", x"e6ef0cacd2dad1aa", x"510dc1f0e2c51e00", x"8abda44876ecf146", x"2f918068712a9c88");
            when 31173269 => data <= (x"ab40018c470f1a32", x"d5cd0cd6459159bb", x"381c87f925ee306d", x"74b8c46d073b1d72", x"424ae68354534f68", x"784026701b5e30fd", x"5c9958721435a849", x"8e8d335f9f60a69e");
            when 23149879 => data <= (x"d6283eb7072f91f3", x"f9b1f4c4de2bdd1a", x"f68f60c316db9097", x"5e4476373e66d9cc", x"6862f2c7e6a04e87", x"4e863281f8a08d43", x"fa02a0dacc6abe4c", x"e4682f3ae710c04a");
            when 22118963 => data <= (x"4e212a77747d5586", x"4a6692d80db02201", x"f39e5079fb671221", x"a971ed3da19d7668", x"bde5a6448ff85959", x"c81c5574107a2d19", x"369b63878b2de5e2", x"38e6dafab9fa164e");
            when 27082086 => data <= (x"74e890866d0d9769", x"319867034f0544c7", x"4f70b4e88dd6b0dc", x"0ed0e957a13a9782", x"ba33cf41c9e2bbac", x"0e678e531c95a433", x"c01858327e05303a", x"c459880041ec9711");
            when 30627970 => data <= (x"7a592afe4e0d284f", x"1a08098b6374a610", x"980a3ac86a24ffae", x"70512035aa49ff9a", x"3960ae6e9ee28ed0", x"fdc2ef29e9d8c66a", x"e8c57985e3f1f7de", x"2be1fc6e6acafbe0");
            when 30302820 => data <= (x"ab7bf0d868be25b4", x"d2a755fdbc86d195", x"3be9eb00f9ece48c", x"8cfcfb4ef146b7fb", x"470b184aa9e88fd5", x"1a09c1d4acbec1ba", x"a802ac765eb6c437", x"bfe796c01eb4c606");
            when 28272314 => data <= (x"f316be4ddc10b045", x"b1fe001434bb54bb", x"ee42b3903f77008d", x"353562b0791c5ff0", x"d5eb1fdafcaeed4f", x"2ac8ae4049787c70", x"3f547b1607170035", x"0f9657438885c4c3");
            when 23386996 => data <= (x"382d6fd8d52330d3", x"c44763a9480c78c2", x"e1729dcdcdc03b6f", x"9ee8b738b2bf6550", x"e712388fd0d29015", x"e93cb74e527c732c", x"045e53c5c358b3b9", x"bc4e0ced3b6730c2");
            when 32671797 => data <= (x"ecb07ef6db8ea8e1", x"aa00eb10b3a88828", x"4a29543ccadee0c9", x"c9f161835009db29", x"6c819814712bf764", x"ef7358e424c3e3fd", x"06c1bbcd7ce4b069", x"5c8551bda0ef6b3f");
            when 4527376 => data <= (x"c11a010c326bd381", x"72bd002ed9967f46", x"2a667fa22643b866", x"a58ca7ac6c406e44", x"487baeecf9dfdef4", x"ca7a9c619d647d4d", x"69ee29f564bcee21", x"9bedec8847d34d2f");
            when 31273615 => data <= (x"030551a97d4236c6", x"e836fd210706e45b", x"bcaf241892e4012b", x"8478733ecbad5736", x"71b1d3ec631c44b2", x"2941e712a3f5fcec", x"f262c15cc178c36e", x"da8b70bc7d2fc434");
            when 26185671 => data <= (x"5e064179c1ca55ed", x"032cbfad0fe4dbd7", x"c845ad4500690cdb", x"9828176da157e930", x"6802adc8bdcd91bd", x"95ddaa44229f6d50", x"36bd9f54c090d9c2", x"8b4305492cdcd19c");
            when 31479471 => data <= (x"a5992e66d79e46c4", x"c9c15ddb92300120", x"0e790cd60f74b528", x"2dba81f5b22a0abf", x"443ed51ad5b5f9a1", x"b31835439e9fde80", x"45eb9cc80a8f4528", x"3ea7fd55438b29fa");
            when 19942200 => data <= (x"c26f414e11371f5f", x"3c770b89ecb2a8cd", x"8e8c29f5ab7dfdde", x"a8a411792ec24a2d", x"915e2b0d2671c2a4", x"3921012c7190a17e", x"974dd65b6c09ac36", x"05cb92181e45a4db");
            when 27637921 => data <= (x"bb00db70763a3f93", x"c9d249ff2f294e67", x"091f59246e3facd0", x"710cb741d0f36720", x"c712fb30b85c8f91", x"6c7f409a1bbfba4d", x"67c6f7fad6d12bad", x"54fe2efd5f3648ce");
            when 2784584 => data <= (x"35e8068b3b83c531", x"9d9a4e09b5e5136d", x"4fdd0e5075d6fe46", x"8e05cc0ca3278482", x"bc37b8ed7d396065", x"f3bd2a52c5d98a56", x"983e5f72c2e261c9", x"718fef1dd63f0a5a");
            when 8276951 => data <= (x"74d63d719b36046b", x"d1d91eea6209f45b", x"db79bf58952a18b9", x"c36629d744e3a57b", x"16443f5835afdb3e", x"df6d59df753c8c42", x"c13efd6b22cb2fc8", x"65a88611e130ca40");
            when 2255872 => data <= (x"bac87704f79f0890", x"1772cdaa36580c97", x"a4c18b382ecc9b0e", x"86b737623809176d", x"9630c7f43b995a13", x"4566171771d452dd", x"d58cde37bd8b4f31", x"ff7e70e5f5de0f48");
            when 17408880 => data <= (x"ce133968bbdb0b21", x"b4afc3c7b0f412f7", x"363417d39c12b660", x"0238a88ca825213a", x"6a339e6bf07577e5", x"633dc9eb6bdf8f77", x"9687dada0c8c1b70", x"38f5c739a25053ff");
            when 31484745 => data <= (x"294fc94f48c16f8a", x"c5bcdbd14ecb852f", x"ebd6d860522fee39", x"631dc616a663d6c5", x"3091226d25f5bb45", x"744f35c136742d23", x"4e3c1f2932d298a8", x"05c00f59d49f7298");
            when 8936680 => data <= (x"f10a61a3bedad151", x"7edd1894f63e586c", x"d7a61d10fb3fc9dd", x"c8ed7face46992b5", x"9fe050e593885fbc", x"297ead6f4a315cec", x"d28c05b01b3feae2", x"b8c109bac35520aa");
            when 12200391 => data <= (x"3d2224f775724c93", x"89d44429458f4daf", x"d91715716282dec6", x"d417dbc79b1ed494", x"50aa2167ffd20a54", x"48c1d379566915d7", x"c8fcccaff014187e", x"85f833bf3ddf1d4c");
            when 7281516 => data <= (x"4c7e86231bcf9914", x"5b7e3d317dada7df", x"106ff2f1d9007279", x"ece2b3a3eb15f465", x"5f63195da1e63c58", x"d1913cf6620752ba", x"bc1301a2ef8364cb", x"12ff797bfb7d55c4");
            when 7652649 => data <= (x"8ce52db4a93c8f88", x"8bba2a23b382b4f2", x"4d7a4d926c8883ad", x"b3c1fe3e95f8c577", x"7e972daac239255b", x"21c5478125290987", x"5bc80849a70a6f9b", x"0f6fc70e1916bdd6");
            when 12475514 => data <= (x"fb7d13612db4f786", x"aea8dcc1e4d32c9a", x"0810d5dc8d2b28cc", x"f91048468afdbe18", x"177ce2e52c6e2c5c", x"872d24721126ec80", x"26ce191b065b4eb2", x"ea8b6acd7ecc37d3");
            when 11539346 => data <= (x"ce6c9efbf0e0dec7", x"52068b13985cb2d7", x"a05d1ee6d0022daf", x"df9bfb76096c171b", x"24d9ab8cf20b9231", x"218cead6bc77c4ee", x"8adc78af5bb4c6db", x"44c17a813cd4ff83");
            when 30451146 => data <= (x"371aa5810ebc1062", x"e5d4164d4a5ad6fa", x"d3502419afc5df5a", x"cda4427185d6244d", x"ca549e5365379878", x"55f8977418a3ac9a", x"ff2bbdbe3da64c8d", x"6da81e013a04b6da");
            when 13694212 => data <= (x"80b310e9977ba464", x"56fcebfb94e2c2d8", x"ee06b237380b75a3", x"4a4ea0fd5e87a8a4", x"098ac3bbaec82cb8", x"c8da9987d7f90714", x"a75f91fd6b1cc51a", x"122b69148f229dd1");
            when 28074187 => data <= (x"ba2c78fa8fe57140", x"559286e49bf577c3", x"574e6af4dd29a33a", x"ba52caf70da473be", x"6395c711e0d2442b", x"ef13b962115573f2", x"d6f03d17cc09c99a", x"763279c69c305701");
            when 33038657 => data <= (x"f940a74ed4fa4d54", x"4facae73f29977a2", x"51acf9491d78b42c", x"ed2a89963e7df4ea", x"2a191725fea5876b", x"f8de9e36bb39f5e6", x"b97d652dc22c58a3", x"f8ca744c0bd5105c");
            when 6635425 => data <= (x"c4a8f1cbe120e362", x"5dbcd3b1d58275b7", x"bdab74fbc9770221", x"bf76d48d830c2339", x"cc549d8ebef7828e", x"8b812ec4a7234c56", x"996c141f62bf9f61", x"6dfe069ceed11d9f");
            when 28045090 => data <= (x"2d590aee516de32f", x"a6b4516ac8dab1f7", x"c16bae2dfc1f15ac", x"a9e5518af420f850", x"face72524c256aa6", x"a92afe565f6782e7", x"014bbc11a31a67c0", x"b136b75f844f8256");
            when 3040230 => data <= (x"46581cc7d7d53cd9", x"410205d90c450bb8", x"3699d5efa1846169", x"69ab4db827308829", x"0e2ccadb8508b150", x"24b4c3527ad92ac1", x"d94275a0be1e2ae0", x"f35d065d3656792d");
            when 33919242 => data <= (x"7edddf48027fca06", x"6faf61b9b1bd05a7", x"b8e802a6a316aa34", x"7bc4b0c9e3c46855", x"52175c258018b0f2", x"2565fccdc6de9a86", x"eb7e90a7fd9acdc8", x"ebc195bc07e4d135");
            when 21363009 => data <= (x"02d0e20643833684", x"2485fafba5c211f6", x"ce608d0acd8e6fbd", x"d1bc3cc38aea3122", x"40856b220466f9e9", x"de1b9518e8053c9b", x"c1dd37c0ec935e11", x"f105bf6914cae433");
            when 13305047 => data <= (x"b8fe8bfca4473544", x"0e058891bfe2ec47", x"95ee4095dc468c49", x"e1032684a1107745", x"90e1867a70d0d590", x"f0efc9fed52cd445", x"acbd9085a6a6ee81", x"e1198fecfbd186aa");
            when 23305727 => data <= (x"434f1d5265897fcd", x"5687110e13e31d68", x"db0121f477fc6403", x"ef12113ea1d2e142", x"2abfa5d7f6dc95a3", x"bbd9513f7f5aeae2", x"6eda8f4a3c2b2744", x"e64d4244845ea8a0");
            when 24401390 => data <= (x"38f7b3b385c7994f", x"15e6b8f9c6545314", x"8aeb39cd6c840913", x"28e88ac6b43e4f31", x"2f2506c5f43ed3d7", x"feeb670fb741e502", x"054509143ea911ea", x"a4a2add55768dd8d");
            when 5547341 => data <= (x"ba586116d9a8254f", x"148468960e0de538", x"33ebc7c9b426349c", x"f0081614ca8ffba8", x"b2f61af042ac7d3b", x"74421cb4d75ca0d4", x"7299d2f0f2de27a5", x"5058d9c16649be4e");
            when 22901875 => data <= (x"c4cd22058dc2a51c", x"dc4bd9a04c0f5827", x"2482a65528024cd5", x"f9ddcb826dafb4e7", x"82e710556f80613c", x"134b20376c06fa74", x"0144ed57e714d656", x"bba85e66d4213b76");
            when 1411972 => data <= (x"9bbb9fd879541fa4", x"a3dd7f424e9dd637", x"3298d71bdb6aaf4f", x"a7b2252935fbf69e", x"099fbf8019bffa53", x"99c7631bf15f881d", x"b5d1942ef3035f93", x"4fde2e24aa30f5c2");
            when 3784684 => data <= (x"635ac2c9545f188d", x"08761a93c2191269", x"d44338bd7c986b16", x"bc731328ce906611", x"25684359638fa40b", x"4d04f0c655ed8c92", x"0c3665c37c8c370b", x"36dfcdc24a80a3b0");
            when 4055217 => data <= (x"966a86d7b7a909c8", x"b716f4b3358f424e", x"06b0ca485b48903b", x"892ffda574d4683e", x"8538396dddf801c9", x"448ce40d9567487a", x"b42584aed4fd6c8a", x"180c163dd9ed82da");
            when 24757306 => data <= (x"5f80283928add22c", x"736e55fa65280bb7", x"2d26558df72f3884", x"e1dc8d92c0aa324f", x"1c0727560deb22d4", x"688d112f88c810be", x"24c8426a5d9717c4", x"6cd05a9ea40c5905");
            when 31727731 => data <= (x"b2744563b6712f1b", x"e52ff00fab26a02d", x"2b368e4ddd75795f", x"3cbb6f2547909569", x"abd411637bc1293b", x"ff8c83fef056afed", x"486003add1f3db9c", x"2465d370c1d96951");
            when 29368350 => data <= (x"34a6a302c271c85b", x"ac4d9dd001462b33", x"b0bfdc2372d68622", x"6d6c42368a1a08e0", x"14fe9e143850023f", x"a7036e3a4a59a199", x"8766838d734111c3", x"d850911cec1f4ff5");
            when 2136542 => data <= (x"efd0c2ef3851d1eb", x"3531bf964d15742a", x"50a61ae54554fe8b", x"2cd253eca7546bda", x"931442ff3169fdf1", x"24ab158c1ebabb41", x"a434d12f08156ee0", x"f47aa5fca917feb8");
            when 19087838 => data <= (x"100e6a55f3e75de1", x"ee3c93247072338d", x"6e881f8ee8a76eef", x"b1a5c56efe0e96b3", x"aa3938e9df8034ef", x"8d0d6a942870da8d", x"653eea45cf1c16af", x"cb28bfae97c692cd");
            when 27224490 => data <= (x"fd71823f396d56c0", x"c035eeea318f9c20", x"24ebce01515c8204", x"9f7eb4db9015198c", x"7d809d6ff5310665", x"f47b7d679e45ee64", x"136cb1f53477e428", x"fafa12fa781338b8");
            when 16699077 => data <= (x"b5a016f67fc2e2e8", x"290644aadd559906", x"47039e0d4aa35afe", x"4f86e3a485301768", x"5e26cebca936df30", x"1ad38cfd4ebe106b", x"26ddf2791eb64d7b", x"536ed599eaa19d5b");
            when 17924116 => data <= (x"e56b2ba8f54db37f", x"86ae727389435944", x"0b6fd8e91aae2d11", x"e38f9d24fbd05484", x"b312954cca108c06", x"6304c53480bd9c10", x"c54febaa3df43644", x"18c1c9f15eb48f98");
            when 27247470 => data <= (x"3ec75f7e8ab50502", x"99d793acaf3da3ac", x"fc63053edd20ac35", x"178ba823fd6464d4", x"68e12d7030b43fca", x"481bf8a19c514954", x"d78d986867da41b5", x"a2418d4d7a2cfc69");
            when 32649567 => data <= (x"97f90cf08b416e88", x"597c9dc51fa678c3", x"591c80b03fb651a0", x"cac4a008451d0222", x"44c3c521e7d5edb5", x"2deacd4f819a78d7", x"df8e1f8c2de98a9f", x"1980f70243fb0094");
            when 17237547 => data <= (x"80a2e2ab9d78d057", x"300ecd3a7f895d91", x"eafc1d3d1990be74", x"3272a5e90cae9a96", x"d181e733e938a9a5", x"fa4cb15c61be0fce", x"66b89ef12e721139", x"bd165c0d744cd363");
            when 30311448 => data <= (x"383458fa13d02298", x"fe9629431055c2d8", x"5c1b0fc05f5785b2", x"17ca469ce086e158", x"d3c04d55b43264d9", x"e46fefb9cb9bf8ec", x"556785b17e0fe7e2", x"fe4205dd4fd06712");
            when 5294696 => data <= (x"f18e0206f9a5b899", x"1f22c54920aa741c", x"6db62488a70c5959", x"182dae45fdff54ab", x"cf4f0ea91507de34", x"d1a910a888fabc84", x"0346992607d089a5", x"299b33bd0238f3a3");
            when 22579215 => data <= (x"8990046c55c3ed19", x"3db3da1e61dc9226", x"165593c4dda6c206", x"956836f4ad4efba9", x"eceb6dc51292e884", x"8d5afffaf3c6e199", x"06f977ef50b36a54", x"2e22c7fd929fd65d");
            when 11317517 => data <= (x"000e6f570bfa4ecf", x"bfa776ae95eab174", x"69ca771e4ededaf1", x"be0a6b897c52743b", x"44a5ad165c900b41", x"e8a46ea129f504ef", x"f7f47fe8da162a81", x"3389f93ce859cbd8");
            when 15397336 => data <= (x"6078066243a8850c", x"ae03b82b69a67c79", x"b1232c48aed50db0", x"7e672a8d09f51b4d", x"e1d5a3519b259279", x"1be893a2fcfa043b", x"24a882a26d2f8637", x"f38dae7d405d4a9e");
            when 32177501 => data <= (x"518bd39a47786f97", x"a4968448a3988bef", x"d94b6cb7edcc4670", x"a6e0c893d9160c79", x"f422e1b92ddd378a", x"b0694b98cf07537b", x"2dd4cb23efef667f", x"0dfeee4e83287501");
            when 30770453 => data <= (x"8822c767e30cc9ef", x"d28adc40a44dd702", x"98f0de6cf347d32e", x"5b22d5cf8be4870e", x"342ec937d1015e16", x"7b84fb7915cc8b8e", x"456a9d76d91456d9", x"4c9b864017dfd474");
            when 4523579 => data <= (x"6c4b597460b0a263", x"ac9dd65c85bb275d", x"9e6dc90a6906a319", x"cf5ce5704cd8bc73", x"90b0cc23274e2ec3", x"ffee4f0fdbafced2", x"16e566fa3fff9464", x"a08f835cd024b556");
            when 19863879 => data <= (x"796e9783351661d3", x"ddf5248a5051e1fc", x"c4fe43e3774c283a", x"b22975ebdd1f1496", x"e7ee2b0810beffa5", x"2c4c632ff6e03b52", x"13b208d70bf869fa", x"f9bf8c19fcb7fcec");
            when 8801014 => data <= (x"ee7b64258c0d3c4b", x"070e59ee71a15143", x"5214184956cd2a92", x"ecb9e06ec547fec0", x"77e13ea95e795c66", x"0c41d6e842ae787e", x"427c3b738014c594", x"87975c2a2d65d05f");
            when 9786011 => data <= (x"77e6571076b073f3", x"9ded35f56b159a90", x"574290bc10afc6b6", x"ff54b70ec0407390", x"db1886cc4b3403ba", x"11f245be432e9b77", x"369c2b802ae45c3b", x"771c66834150f960");
            when 33014119 => data <= (x"00eb9f428ff850b7", x"b60234a46304083f", x"03ed75ca234c353e", x"cd6e6e341636f626", x"c370529ed53f9a7a", x"afa2d1a98b979d89", x"48c9f5492c69f0f7", x"7f57f19b9b0c9e34");
            when 8594016 => data <= (x"d43621fd9318a0f6", x"fab5a4498a1f947a", x"b5ae22b43394c595", x"2d36af1a19a1d36b", x"4d90751308deeda4", x"e3e5df7db7de5657", x"eb8594c42453cc2c", x"fdb6cf0660ed08df");
            when 15654688 => data <= (x"d8058115c01bd982", x"9f68951ae6b98353", x"f4cf7a52f9b038d5", x"0fb32a76fb7e371d", x"7e410cac527ca86a", x"f2bdf852d504d735", x"13e84faa824a02f3", x"6c2b342f09e0c881");
            when 25476177 => data <= (x"e86bd0f58dfd5bac", x"08e7a73cc0358298", x"923eb9b40ea6c307", x"d4690cd4cba71a28", x"138ac9ba2fd28936", x"26334e57ed1372bf", x"ba7f67bb7e5ba81d", x"85b6c3d04614c18a");
            when 31894419 => data <= (x"fabc2bb0a0eb8310", x"2bd09dca7e26211c", x"7309ccbda4bccdba", x"575d4b9697901007", x"2a2624cf42aac2a5", x"08c6b147835e4de6", x"22d96432689e6c12", x"14c20913a8384ae0");
            when 26208420 => data <= (x"82edc721815e2336", x"a1e8760c440c63f6", x"c4abac150abcd1fd", x"1c0b0d7c6165397d", x"67af9f1e5852a72e", x"1bfb00f3377f4a93", x"0229a12a3b6ecb72", x"144d7cb8edb3fde2");
            when 32428779 => data <= (x"21a6f934fbe0ac62", x"e9fb466d3dc0cd4e", x"baf0e2a6f1a591cc", x"d0d054b5396738f6", x"06567c8cfa49880f", x"49671d89704683c4", x"ec6afd1be5a1e94b", x"50476a54c8cff166");
            when 31548608 => data <= (x"3b7656bbd9195359", x"20d742786d48c845", x"b2e1cdc8b3d57133", x"43296b4a68493460", x"67404de7cea88622", x"a2a0641b5c814fc3", x"fc626018438e53ac", x"c003c0f103b1a678");
            when 19860951 => data <= (x"456d1c29455def73", x"d3c148cd9be45fb1", x"27da6857c7b7463c", x"cabccae69c8a3ed8", x"6873ccdb305e27a2", x"99d0c4fa66941638", x"c4edfc71945958ad", x"6f5123a674b90fad");
            when 20844171 => data <= (x"d443a22a87924733", x"74e3caad56686c6a", x"43647c2722e58f9a", x"6a0872b25dab7a2c", x"966c5a9d6abef52d", x"078a5a5db859f9e5", x"9e82839075f812b7", x"59c96ee9aabc5b88");
            when 1810451 => data <= (x"61d67ca5674b6fe1", x"900a7f37bc0b1d1a", x"46b79c27656cbc17", x"a85ceadd30f29af3", x"6d8a29ac63f29d0a", x"8fd7087c1e015ecf", x"fff53ef0327dd67d", x"3bce4797d89aa47b");
            when 21771173 => data <= (x"e264e9c6a4e56ff5", x"88aabe2afe190f91", x"d376582fe3d9f4f5", x"e1d406aa99ff42d9", x"86aad9f6e37c4a69", x"6601a1fe7cfc0da4", x"37baa181431f0b3d", x"0905bed6ef69ead7");
            when 15088377 => data <= (x"21012309eb68aa32", x"976db1a0ef62f39c", x"31ee61b5fc749601", x"79f316928c175014", x"c3cb3daef362c72d", x"0102670b08b5e8be", x"d184e6e91abca1a0", x"bda25d00877eed9a");
            when 27374085 => data <= (x"c9ab0c1a5feb4c62", x"437f6693ba68d2d3", x"b548293395047772", x"0ecc4864a2b5b983", x"1ef452befd454bdd", x"bec502836ae92580", x"b4adb53e6889a4e3", x"ae6bacf46caab021");
            when 810796 => data <= (x"a0cdbbc31b430d8b", x"348d3c4945585f2f", x"29e7dc8b41e85d89", x"8dd12e1ebf5bfe6c", x"93af4504f3b613a4", x"38ff90cd63070064", x"96bdc99d0db18678", x"3f42ee28477d2c7c");
            when 32166975 => data <= (x"ee6c995adda51c98", x"e99c4ead2a7f9e9b", x"512f996fe86fac03", x"8e8bbbdf03565248", x"0c8b831f0433dbf5", x"9907a04df555d32d", x"fed1fc3333d9c377", x"efd2b9bb64e5b7f6");
            when 32625402 => data <= (x"2aef0747b3c51491", x"847db461680c762b", x"b334b69c8bc64b05", x"15efa2a563e343f8", x"6826d7c04223772d", x"a6bf0922693e7441", x"45cdc22cc14349c2", x"c1fa297f392e46be");
            when 25722828 => data <= (x"c710be8c2fa3e780", x"9f301f0b023d8d29", x"5c2ebf854ca141c0", x"03057041a48c78da", x"6f3478e804aab1dc", x"92ed55081d86d971", x"851d19e1d51d45f0", x"eab867276d7c4003");
            when 5404724 => data <= (x"044e7f789c58560c", x"4d9b74e1e56de10b", x"05eb2d85cb5e6506", x"0fc6b779f56a76df", x"9e968cac7e8863a9", x"53d5b265750cade4", x"77d0d5f4f9e2e85f", x"cd6c53ee823877b7");
            when 30618224 => data <= (x"b46ef5fff6f79e55", x"0c76cb9ba62f3af4", x"14e5fa3e0a9fb285", x"693dba83d29305cc", x"4684adb9cafb71b8", x"3cc438ecd97b84ce", x"7255281e993a9ab5", x"557806674cba6ff1");
            when 26373436 => data <= (x"26843bd26e2f821d", x"60a0d2f990d343b5", x"0bd295597f4e4c25", x"215fa0bfd2aa0e8c", x"cc1de20adc75f0ea", x"d30a26cd14b89d97", x"647adee9469cef58", x"4e7d3c1c83767f33");
            when 26776729 => data <= (x"1ba0812a1d25eaa6", x"e089d2195d56fe1e", x"89c9f5da85787d42", x"f98e3e329b6e369e", x"305fec3e6281c698", x"726b5d89c4d765f6", x"2726842b9b50d22d", x"2423f87769dbb37c");
            when 1490184 => data <= (x"397db918fd3d7e3d", x"23f926cb1cc76316", x"f0e7738a74dbdc5b", x"e60b65e9a96bd2ed", x"5b8f48c5aa7cc109", x"d323f319da979837", x"48b735214557abc1", x"d2be898b960088da");
            when 8851637 => data <= (x"e24e6aa0e8292c30", x"aae7103b17b8d7b0", x"a9a50fc67620a155", x"ad6ffacf6022a03e", x"b7c5df6972f1c517", x"de17ecbe9d8066c0", x"ebcc5b273c899f80", x"89e140d423bfadfc");
            when 1282942 => data <= (x"b90045d41bd0dede", x"d8d96f05f42d55e1", x"c7cf65770d30251f", x"44609905bb148c6d", x"4daf319f7ec82336", x"56b5d51889d842ca", x"989bb662eb474db2", x"5a9c5ec14f17c39d");
            when 7170852 => data <= (x"d2bb6c9117c65e74", x"b1831ef9fc456ef8", x"9cdfa439a739e53f", x"b3b16519677a4406", x"f00d17822a1ef596", x"d67503c0c0d884ab", x"1265dbc809a3fdb7", x"91cad462a6ea2785");
            when 14419081 => data <= (x"d07a3791d7a5cb09", x"2cc0814615a1bd84", x"25986c9d83e38f6b", x"834885ae74492ec5", x"f228d90ec8eef7fe", x"a43e647dea39f61f", x"2036d75ed8ca115c", x"ffcea0edfdc82720");
            when 8181793 => data <= (x"e43a86bfdb61e83f", x"e878161070889188", x"23a4a7960120ee6b", x"e279795256351d1b", x"e1eb7c2d057ff403", x"8a3f1e528c8d5517", x"cb0f76914d268fca", x"54722589595ab8b2");
            when 17347914 => data <= (x"9e2b842667732dbb", x"fd44443dbbeef389", x"ac02c901a8693607", x"42c71dece261ab5f", x"93a79cb51aba3da0", x"0c27267a0703fbdf", x"e517bed20eff7fa0", x"eec24b54e6954e71");
            when 13578055 => data <= (x"142bfb15cb5b4477", x"aff238ef3e2269db", x"3772b4cd22ba8a70", x"840ecf27860ada57", x"6b68d045467c660f", x"44c2b1545e584a19", x"47b7c29234328512", x"06b9b3b56be11539");
            when 18710901 => data <= (x"1b2685ceb0b2555b", x"9ba5f6274b77a411", x"67d220799714705f", x"d94760b5bed1b48e", x"22b7cf4a229922cb", x"65d1d096c84615bb", x"9fd314fb12246a6f", x"808c2f7757c15b2b");
            when 9271404 => data <= (x"0e85e373758f6fc6", x"5699a5b35b88b72c", x"5abe9913e609bf9b", x"dbab18875ec3615d", x"7eec609ce619b971", x"29af5fe0c1bfdbdb", x"6368548963f365ee", x"c711b44dcd61bc31");
            when 17282616 => data <= (x"c9104da6f4974788", x"1c95bdac272c11e7", x"1a91f56aef4882b9", x"1caa331682fb66ef", x"91d27ed403fc5389", x"6bbfdccdfb64dad0", x"b2e9d2d82bf931c2", x"98fba22e192b4a4e");
            when 12494468 => data <= (x"b1e7ecff9a11e7a8", x"cde171f0be3e1277", x"ff1e8b667a749ccf", x"3ea29e55b0f33f03", x"f867e7ef6d92957a", x"8e54050cd072d104", x"4582d1298d3dcb6b", x"2942fbaebdfb34d4");
            when 20033213 => data <= (x"e524c2b77b1f125e", x"cc4dfeb94482d873", x"988063aaace9c4ec", x"5f21e782264c08ef", x"7fe9e301c5129bc3", x"24854525f29a7ad8", x"3c9a488fb208b1a3", x"3913f969e8251432");
            when 9114220 => data <= (x"b742059500431822", x"14823e22d120379d", x"1579852ac80f394b", x"a61a30b2049bfb22", x"61b79fa3014f8234", x"7b89a3cd725fb99b", x"a11d71b7253caf1f", x"07e204efe833352b");
            when 16738881 => data <= (x"baf076dab7fe0fd5", x"605fb0e0fe29ebcc", x"ecc84f0e504aee10", x"4d3a98ae640c1083", x"f6cca5d3fe7182a7", x"58c5d92b1e47eff6", x"2e902c81d397a75f", x"3a896b8d43311162");
            when 1353868 => data <= (x"2fcaf7bcac28c9e7", x"c2c29f1a41c4b599", x"4d1745c41630f883", x"ca56fab73489ebdc", x"9db996d1725bc5ad", x"0383109ce16b66d4", x"c155941cbf3ab74e", x"b39f75f67d178326");
            when 13758597 => data <= (x"afb67999bee4c218", x"e02bf55eb8fd42ad", x"2f0d0ae5bda12328", x"1791db1af7e2ff47", x"bcab45dd9318e4c0", x"62270d9cbe6262fc", x"b95b1fd6b04c5d28", x"f75be249039f8e2b");
            when 32946578 => data <= (x"d0f9cd3f6e040949", x"8508a398c2064858", x"dbfba7ad6ad288a7", x"d598a6ff3a25a03f", x"5c2f790fde10881e", x"352433d01658480b", x"12341f6a46f8d568", x"add7555d8d0ededb");
            when 4869880 => data <= (x"fe18d3ac844d3202", x"c4d23b7950bcc183", x"474dc938d1f47283", x"06b41efeb5a4007e", x"83f230221e5709f7", x"f74f714526f3cf1a", x"b94c6a65d907b85c", x"7c954f6a11b7055d");
            when 2657076 => data <= (x"50262d6d43bcf4ed", x"74fa44edb1b76dfd", x"4f3a1a252d8e146d", x"77f534ea2beaad02", x"4de260a48014a3db", x"b78f543482db8e1a", x"5b7a090491df1d6b", x"bd5375c35e9dc793");
            when 31774067 => data <= (x"677744ece8035058", x"3c20db314d2cb38a", x"6da72ce9e5381d73", x"e9984a54565dc765", x"4442cba1a7a6d88f", x"1ab2b6da3b4945f9", x"c115823a318e26cc", x"13b7bf9f8fe1408c");
            when 26388387 => data <= (x"118007f093b3584a", x"bc2e7555802671d2", x"2dfe6e9c6557af75", x"aaae46ebd62f5beb", x"6d3af0dffd6e3ad2", x"ced9dd0488a172e3", x"ebbff9817c382c73", x"1298bcddffff287c");
            when 19813737 => data <= (x"86d06d77b71cf980", x"97ac3647b48e6a22", x"b91b143ee3014daa", x"5610e0077e8b0503", x"f68bb3f321fa5d5d", x"f52d9f7320a14080", x"8832b29e4c262853", x"8073aa91c6bea49f");
            when 21318862 => data <= (x"7900d2b0d2700e49", x"c98050c5b6cb2f2d", x"2ba9a29996670e63", x"367611aac2d9d72f", x"667fced50b7e461f", x"ab3bff7eed89127c", x"8d0bc1531aa8c3a6", x"d21c853fe0e51ff3");
            when 3407291 => data <= (x"24f10fa4dc5691c1", x"25672f2fa072501c", x"63a0443bda464696", x"66abc8d43fe37f79", x"a1a77a986691cf87", x"fab59a4cb8c5e676", x"9f67c3fece77fe2b", x"18f7f15a6a9a2d5b");
            when 20729364 => data <= (x"57e61eaab39cf188", x"8690d49b1b2706e7", x"b502e251341c7948", x"fdba0a0116c0589c", x"9a7d7f87db72ba68", x"7aa67b08fde3f139", x"2a154cd3fff0418f", x"974a01c15c8a436d");
            when 29761089 => data <= (x"38cde5d2114be82b", x"75a22b696e72fd2f", x"03925d3335b32af5", x"a2e3b4879af38888", x"604ad3c59f9c91ef", x"0c64bf3d2e8954ec", x"8497299ec6b31e93", x"7e3c329b0047157e");
            when 24628276 => data <= (x"06624ca486a508a2", x"1a64b78b2b571be4", x"0cf216fbac66aace", x"0b560f917b2e9d07", x"97f5f95887525c16", x"0f3921b6166c1a51", x"df632d8f2e132617", x"1876cad40cf5c4e1");
            when 25819137 => data <= (x"953c9a9869f11289", x"edd5d409ff2ce44a", x"4cd4f2e431ac53bc", x"0f5da4a597d6d36b", x"e69c5bdff353ccc1", x"2acbbadddca67226", x"b0e2466a66bcef6e", x"246a1b4bc06a8b8a");
            when 33740791 => data <= (x"9213a55e4444a197", x"87bb4c3eaba985f3", x"f626c6394fc6aba2", x"f7083b5d4cd8333d", x"c8b86342929cda60", x"c676ed7ccb1ee664", x"c6c3cf93b16ba79c", x"5ec5e17936fc171d");
            when 2487401 => data <= (x"0a8b50ad2a9b2a54", x"6951d29631064397", x"3840c5f9177d7324", x"913cd95d8d01ddfe", x"0d15deccf324e019", x"8df2a35175244dfb", x"9a374a68ca153381", x"310e2ab600454d3b");
            when 9019955 => data <= (x"40c42ac46cbad9f9", x"1dc8624b2652bcd5", x"180987eaf06bdee1", x"d9be22bca1cd6c57", x"3286b7e0d8789e0f", x"d5e0976e940a06c9", x"2aa89771321ce219", x"94ca3309b5dc173b");
            when 853960 => data <= (x"6eaedf314b0e22a7", x"6276dc7fbceef7d6", x"6728cc410ba3dd8f", x"cb0bf2fcc8a46504", x"86fb98def281cfb6", x"e40ee8e2888b3335", x"1af090303fda20c3", x"622c8d7bf6cf6083");
            when 29918787 => data <= (x"09396a63063f6d63", x"2b8e83342c34b294", x"7172d05fcd07d648", x"cb2dfcc66f16614c", x"d294fd0bf6ef2590", x"15c2382b274d68b1", x"bf9d318438876ea3", x"6ad27195b7cdd4f1");
            when 3577266 => data <= (x"072e8763dfd0829a", x"6ecca36e52f0ba75", x"037455a18208903e", x"9bfad67fbc4da0aa", x"2fc73f1a400123df", x"2759442e9d6f7ef4", x"e6ed5ec649451035", x"912e2a369ae0db2c");
            when 7985927 => data <= (x"18285c651ba61c53", x"5bef40afe07b5b93", x"6cf4cbf80682c412", x"ab87428cede0fd56", x"81661bc737f401d3", x"85643a20c190aecb", x"f0ae600c41521822", x"c39a4365e424c472");
            when 9955133 => data <= (x"ff9a023da8fd3723", x"411a0a267b847ef7", x"0ca2fa95b795aeb2", x"2c5c2ed20d07a6ed", x"e701edb4c7ea54a8", x"0cf26e64972b05d9", x"6cd105a09b86f2dc", x"44697f90937a6fc1");
            when 18666198 => data <= (x"ea263c0ba3ba16dc", x"a3f8f457e6e98898", x"2de4d1876026ce01", x"7cd81e23b2a91abe", x"4c6e621daeeb336e", x"77fb8ca5950a01fe", x"9a1bc59145215566", x"7109e0721d701c3e");
            when 9894479 => data <= (x"18bb22a158eeb1e2", x"9df8b591cfa14b81", x"f98387ae40333205", x"ac722293955dc445", x"414ed6b2e87d0053", x"3224e9fe52641571", x"7ad007e364b29c64", x"93d3c24ef08d6f3f");
            when 28046891 => data <= (x"48afcb89610db8e5", x"967e0e3cbe942915", x"d5a0a115af1fc324", x"17f7848c7a616083", x"e8469c4e21e42c18", x"548b51b65f92c8eb", x"546047c1737dc9e8", x"27637dc280f0b0e4");
            when 5024427 => data <= (x"7b5149337df23472", x"92bb4612b0115c6a", x"a1adaf8c496981b7", x"ea428d8fd3c44441", x"4960f900d10c7424", x"2ff1e7f39e96089d", x"b802e0a0ac519486", x"12487f6a3bcaa80e");
            when 23758844 => data <= (x"21bbef3415d6292b", x"13bb8f58312144b3", x"296733454d07d2cc", x"31f60e9bb0325458", x"d39bc4e10a70acb7", x"b6c64f672c945a6a", x"174049d99cc487b1", x"b9978ed8fe5f08c2");
            when 14673414 => data <= (x"b23df5dd3dc855f0", x"2011f8c48823ab6a", x"9785294b3f84bf6c", x"dc667a4312e2e75f", x"fa79bb3dc2e4c457", x"b641546774ede469", x"34204c2afca2e3fd", x"bc42773bd825d017");
            when 17700426 => data <= (x"8aada88634ea388d", x"1608cfcd7e88748b", x"6c73382f666de7e6", x"68db261408f06580", x"a84331850302c1c5", x"f8b5241f01763b4e", x"fecf4a3bcf6d3234", x"a9a2f59d7fdd6d28");
            when 22420071 => data <= (x"8f031707161c3bdc", x"4c3a010429bcf728", x"209aad4f8547d3d6", x"9bcbddd6892c8d50", x"e500c29571445154", x"71d78d5f0affde31", x"b34d6692b906685c", x"5c7be3cff07f5062");
            when 31378495 => data <= (x"49dd03ff8b650e2a", x"2c6ee0032d0cb328", x"3fd84866846c0dae", x"a824bfc63ba8a529", x"a43de3498c2ee147", x"ad42e10427cf014b", x"d57dd54db874b699", x"5ee68b0731817f16");
            when 7602316 => data <= (x"6b59fb4d9d0ce6f8", x"e282d61ccad51de6", x"f299b70a39936e7d", x"b3b61370e5831016", x"94f573b3429cce69", x"f22866c6e60b3d71", x"11a473ee40f8ee32", x"a8fb16412c85f4fb");
            when 13271091 => data <= (x"793a4aec929c99ef", x"e909ee3ac286d485", x"488783f5aedd6398", x"12cf2153a808d3d5", x"55af7cadb2f5c89d", x"d3bbc5dc759e77d6", x"57330b92f33f51aa", x"09e242257dd6ad27");
            when 12155856 => data <= (x"63aff78c8bf49937", x"088d1d431386583e", x"9dec6be043a357e0", x"9d1534a96c26a45f", x"559f83825e3b6ce0", x"767df63ba58ded3d", x"8e8230a42f0e6841", x"3cdd3f3fd6a7a3fc");
            when 18925192 => data <= (x"26c7afa55a03cc27", x"c15d2a2a51bcb97b", x"546df3f075a8a086", x"448d0fb67c369332", x"28a2a943b081b20a", x"c8614cc25f36bbec", x"2d58acdda39ea3a3", x"832948fc6b465988");
            when 28132482 => data <= (x"2da377e86404bf3f", x"56c12fd1d429bf8e", x"2e1cc3b62671713d", x"6791f398e42780b9", x"40c94c2899b59902", x"06aea3a25f176a62", x"42ca78dc252baa34", x"4f9b84ac98492bf8");
            when 30996879 => data <= (x"ea1dbe4c154c4389", x"02ab9186a57b905d", x"1312cbde48d8c9af", x"e97e05ce1b279090", x"3ddf80dedb4a1dd5", x"1d239ca703721a1a", x"b2af5e7f39ef7766", x"29145a05aa32c8d8");
            when 452037 => data <= (x"e05039a0b28cff3f", x"a13d0bf398bc90eb", x"b6ea224d7ee966e6", x"42c7229f98b39d24", x"8ecbf83f78e49b7a", x"ed2ccaca0a494d86", x"0366ee6f11455902", x"707cafacd1f182b1");
            when 4929945 => data <= (x"394548ac03c137c6", x"0c9708c6bf9bd2b8", x"8a3b141fdc22f104", x"c2e135ee18415135", x"66a624903aeb7fa6", x"069550e34bbc317f", x"6f934b2d8615629b", x"74bc3b0644516f88");
            when 18628560 => data <= (x"e1a500584574a1f7", x"875036b2ad92c82f", x"477383b2fa8fabe3", x"cee90a41a68c4140", x"fe364cc826ad9bc9", x"e7756e289949436d", x"ffb635b890b4aed2", x"ae4b6b84a3d293d5");
            when 24375656 => data <= (x"c24e567ae360bdd7", x"d1b67b057eab822d", x"1338b4d50ae56d87", x"ff89d9d0cf37592d", x"509b76eb4ae97da0", x"bfb82fd7623ecfbb", x"d19f1f1d10a680bf", x"d8296d4ca09277c1");
            when 29343930 => data <= (x"ed56b68de2914c0a", x"d84350f58aaac66a", x"a57d7475282255df", x"e97598742b1faa04", x"51446eec2809793f", x"85a13ae3e14d5e45", x"f0232b56476d07fa", x"5e014239ac4e0912");
            when 11449529 => data <= (x"414cc15f022f2d2e", x"bac99ec58043a621", x"13b3c8b8fa915a4b", x"584f8f2a1d4d02ef", x"7ddcd6ab1c8c5612", x"fd00c83aa7b00717", x"467de9333bbaad62", x"3f3f4e64431d3500");
            when 19813392 => data <= (x"ad9f0741ac5925fe", x"b86760d6cd59e2e1", x"613c1bd8ae8963d2", x"1c1f696d44334f81", x"b67a7aa2a30ac985", x"c8531b1ce13fc228", x"a5d1612d536e8c2f", x"97a3334714be01c9");
            when 30539650 => data <= (x"5c3ac13d4206df62", x"8492b0a61bee69b0", x"6b7d5eed8ac57d90", x"3d6ea5a45f2a6bd4", x"a130f209c6de16bd", x"4293d8876ae07c42", x"bc1e33fda28375ec", x"def4562acbd6c466");
            when 10793674 => data <= (x"a0f21321f2e7b00f", x"92ce6416453d7d10", x"b04a67582156b1c6", x"d8e8f461bfa4d8dd", x"af7e1cdda2a09c01", x"97eedc69ba4a145d", x"1c92c37982470db3", x"58c241d167df6bb5");
            when 12840170 => data <= (x"4aec88dc33322549", x"ae6b9567475a0415", x"d02c40d1bb48d342", x"e077819b28da2120", x"0d9dfb5f259952d0", x"c5fb7eb1287927ae", x"614e336360dcccbb", x"94b1e4d94d3e5d88");
            when 24668445 => data <= (x"1e8c4825a8ac5f8c", x"b53ff7a7cb92b533", x"e8845c5ddf530928", x"0a9265468f600f82", x"17d491efef18f77e", x"9b3e70e0bfae20e4", x"9c56def920cae521", x"42c0c5a069a2443d");
            when 28510129 => data <= (x"a6c9807532bb83a4", x"da371820236644fe", x"116cf4189e186375", x"6b664f0702f01fbc", x"2bd87be317610cac", x"b7d29bc112b2385e", x"03ffa94f30b0adef", x"cd4c8d6b08df522e");
            when 27651072 => data <= (x"5b9a92e7edbd866d", x"5dfc27801eff25f0", x"cc624dc50eba25fa", x"b52a9f0f2c2ef5ef", x"667cd96c14d9c5b0", x"41f3fb9f192d9782", x"521de0ec56919fe5", x"a80220f18d6a6cf6");
            when 21662621 => data <= (x"3b6272bf8f3fad42", x"c62c212af2b1c3f6", x"9e0f9c6c3967850e", x"16a32cc0dc61c80b", x"fa99582fb6b55e31", x"23634a9bb02e9664", x"f78bc313d555577f", x"4b721a69f1164001");
            when 5194176 => data <= (x"684c58e6aeed627c", x"a0357459d3e75e2b", x"adcf09b4ddd8064e", x"98d2a14bc87b1a8b", x"58e9456d92b86a9a", x"f44ca2cf3f6c6c29", x"6a40a888bb696f76", x"d8f0914ed70d741e");
            when 33261880 => data <= (x"ef61e6ccb817386d", x"52133af8e0aff85d", x"3bbadfd514c14f3f", x"d6ddb839427a942c", x"b2fb6b882a9aa8cb", x"b12d2127196768fe", x"7f6d70c32d374e4a", x"d7b708c377542076");
            when 14336220 => data <= (x"ade182a522560301", x"1af1dd50a36bafe0", x"ac7d588d45d4b5f9", x"39af3cf520981589", x"7dfcc7f32785cefc", x"6ffbc6ee5f300f01", x"96ab857b10cf9260", x"b75987a23f6551d3");
            when 20318235 => data <= (x"05036bb6ad860899", x"5ec156c35a3e241d", x"4ffab658bfbd30d3", x"e15ec336ea5a0b9e", x"91be666f8af0d14f", x"786b96523416f9ff", x"33b0b44b92098b5d", x"934f358068785556");
            when 27461544 => data <= (x"4d1ba7f5f7a72dd2", x"b4f830c7b219cf43", x"a788cb6f03e7e93e", x"6a36b796ffb3d10a", x"b3bd410636e5b787", x"6d70d62fb01004a1", x"4d11610efe96db0d", x"98cbc323d3737bbb");
            when 25847752 => data <= (x"09c6c854f6efe422", x"d49f8154c9b5425f", x"6c8d45d8f7b81fbe", x"98280cc60d502478", x"92b932dd1f8640d6", x"2d22b58230a39fb1", x"0ed7ceedb1769326", x"920e714c9a03dd93");
            when 13908867 => data <= (x"25e72b84a9b847c8", x"275bc76ce80e8ce0", x"0af30768c50d4965", x"78e4cd31d6221061", x"c24ae99a08efe0e1", x"5bfc33d7312e8399", x"d0d2575e28e6cee8", x"97b726bc85099d81");
            when 18824470 => data <= (x"23a62bc482f24840", x"aa9d5bb79c61dfa3", x"16cc22e62ef540ef", x"886ffe843353da4e", x"52f455d879c5122c", x"d0dea10f5a38dc2f", x"f06b8dcf01125e8a", x"5e313d6c73810f1a");
            when 20540611 => data <= (x"ee3602e0f551c874", x"4e70d409460f2467", x"5d56bd07106bc83e", x"9d1f6982260278a2", x"cfda9bc61ee9b127", x"f5984b63e2492d1d", x"48e9acec59053263", x"f7520e10feb38a05");
            when 33585556 => data <= (x"1f365533d51fa8e0", x"f3fda38a0aa40cc9", x"990567b2a038c550", x"50199586768b5571", x"00e1632528a34ba0", x"7738c2fbecb190f4", x"917e39ba72870c88", x"14260dd77fffa8fe");
            when 25351371 => data <= (x"5e3b606323d911ad", x"237842d9890e3b24", x"7ee42f8ab8672001", x"3fbc244ab0172a3d", x"e561cd235c62af0b", x"62d8741efd02cb60", x"0ebf3ce72db63c8b", x"a1f3c31b5e761e2b");
            when 25228829 => data <= (x"7410fed02112a57d", x"e1e0bf2d290568b8", x"935a884a97add5aa", x"4737ee5807a28c80", x"a06ebdabc067abcf", x"48aa38f3c990f06d", x"21a807e8a92c5f84", x"1ef738099ef14171");
            when 28489719 => data <= (x"48de71bed273317a", x"7bb5789cf71ce978", x"318c8103de7c8e20", x"49dd7048da3023cf", x"280223dd6745aaac", x"330e7f9e5c800257", x"31ecd4090bf55510", x"1d19919ab51c7c61");
            when 25036289 => data <= (x"5d80c27cedd682c8", x"c99b76eb42be381a", x"a8cb662a8cbe4e93", x"7287843988b390e2", x"1a70f8858e760230", x"6cc18bf01f0069fa", x"def8910a138c1463", x"8860aa7cc78137c5");
            when 27261716 => data <= (x"f696600664285c88", x"0a09826cb5553a99", x"429b57959cca15a6", x"d6ec42efd6fe6f28", x"e17b705bb2335ae5", x"ca972c0c5cd4c0e9", x"d65c7d4a8454be8b", x"affc02a964d6648f");
            when 32402539 => data <= (x"8d07e9d91642e734", x"f07e3b677cd02249", x"79674e054f337c69", x"0999dff31a5c9406", x"36fd072764f9cfcf", x"1dd3fc8dd337edc4", x"c92cd5ec385c717c", x"dc0aff3fc561f58a");
            when 18889803 => data <= (x"691f7328cfce0da8", x"01fbe254b8fef7b5", x"f7a20811c03e5564", x"8817b18033610d5c", x"8dacacfabe210ec0", x"1f004578356d6476", x"ae861f9d2366140c", x"86560f62fffa2465");
            when 25373075 => data <= (x"a6039b6d2cd21375", x"6689603b6c3b1acd", x"753361b858ecf3bf", x"a0ed07ff93aa6cda", x"550162fbd0e6da8e", x"a3d7846029866961", x"b5b977da3bd2b679", x"cec7cf240be99368");
            when 32027570 => data <= (x"e5724425948ab660", x"b8d3fde08346ed78", x"9778e1c014c0d708", x"0269da3d10ae4246", x"ce9e3c4b2d250898", x"be94e02fb5d101e1", x"981c19db9d7864f8", x"c7162ef23414d344");
            when 8466926 => data <= (x"472f31cdd0fb998b", x"60ce2b644ed36131", x"513789dbc354b530", x"5ee819c45a2b7ec4", x"0bc2d6c9c1f6cf9f", x"d0be65d9d3ad2132", x"052c0884cfc52a38", x"d38531d35c891875");
            when 13500178 => data <= (x"8358dda508a21153", x"dcce76b182ddf762", x"8d32cfa895af737a", x"3a2dc7b1f2d63d43", x"9d71f8c832e8b2d8", x"b83b96c90e57b16f", x"cf646105f8242bd4", x"1aed7e481a46732b");
            when 33132306 => data <= (x"fdca5db4d05e0d5f", x"63b626a08cb8626e", x"342fdc49435c7776", x"0d0e2b785fab772e", x"113ee3451cdcc372", x"e3faece1639ad144", x"02f78f60df04341e", x"d1d03d57b28390a9");
            when 19914251 => data <= (x"9992d2e3bb1e6dda", x"bd8e7117957c5245", x"ee7589eb1e14bda2", x"f5bcfef485574c3c", x"c5624411265da875", x"e7e694c0c4ccd23b", x"7a72216c83818c27", x"dedf2d198bf32179");
            when 15766369 => data <= (x"f1d88e0f98d4239c", x"a13471518c13e016", x"ab954adbf5cc1a2a", x"824b3b52f84b2028", x"31556a8fee6bdde2", x"3461035e52d11914", x"4b2948953ea84beb", x"13cae01111f1e301");
            when 18195858 => data <= (x"ce68c69c3cab0ad8", x"321d11e004fa4072", x"16b990bc874a8c8f", x"c80c9e3157c35189", x"d59434d713b0ecb3", x"69e2ac53ffc91dd4", x"a14eef9f533bce13", x"03bfb029786b881b");
            when 951713 => data <= (x"f72e4fdfd4461169", x"d7b53c196164968c", x"8fbceeace3db851c", x"b08db84b26bb73cb", x"28c8f06a90136df2", x"790c9ea4664ce261", x"4810f05864104974", x"1f8e0efb3d70efae");
            when 31966378 => data <= (x"899497f09803c71a", x"f75a091d7384e79b", x"0b91b18dd139c247", x"a0d1962284eb7445", x"563f788739bb3d72", x"1317a3fa960e80e2", x"21fd1784c0f15556", x"7dd29bda6d37c49d");
            when 26527851 => data <= (x"71058a64e854883e", x"980fea03cfe7596d", x"1320b08e3d487a5b", x"cd532b649c4a916e", x"486827140bfdcc89", x"915592821b32971e", x"552f25a2b7af087f", x"6a5ed93e7c0de329");
            when 5511299 => data <= (x"9a6988951a224209", x"578bb8882a9861b1", x"c0823a679bba146d", x"19023146e356ce0d", x"723b1fe3b639f376", x"cea35e6852a3f50a", x"d43004f2515af0ce", x"c4055dfa67dd879a");
            when 4066034 => data <= (x"a13089be8cafd78f", x"d7c717d49ccdf60c", x"ce23f889f424853f", x"5f53d82416e089d5", x"ba4a77e212068c1d", x"491ac2b5f9d47afc", x"10536a6e83ef31e0", x"ae2a45f2b43da08b");
            when 31185482 => data <= (x"b47f5fd458cbb613", x"bb3a7b3428cd7a65", x"71dbe4511977dd37", x"a8f739da4d50626c", x"f7cf8739bd96ae20", x"6754af8b8edaa943", x"401b03dd316fdfde", x"28283f7f7392fb04");
            when 1468541 => data <= (x"7aa9039cddc57220", x"0be625928b5e9027", x"59928482ce4d5fc5", x"2534237b1a7c4153", x"a76624ada7e89d5d", x"f1bb7cca11080c39", x"e56e29ece60e595f", x"92431d55ebc5e6d7");
            when 22679341 => data <= (x"b626763144876ab7", x"e0d2f2be1a242b01", x"5b2fa9801a489d19", x"0830381695b7a925", x"bd42c31a2146b953", x"4854324e60f66cfa", x"c5e2098a68987d10", x"a989403fa87d41e8");
            when 27780045 => data <= (x"c7cd2a9a3f797bb5", x"a0e8a961509497e8", x"0337a65bedd85411", x"3fd2e9aff4bc689a", x"6a65beeb8e55be6f", x"3d97193f2edc9c2d", x"96450bf0c27826b5", x"1375be5b219eaf21");
            when 3928671 => data <= (x"a73c97c22dacf7f3", x"1645eaee21434ddf", x"73162b84266baf23", x"868922bb489c8c39", x"b6778500602f28a7", x"cd42cd3c4beb00b5", x"c04fe725b85b67c4", x"d71d0944894feb46");
            when 18204660 => data <= (x"2cffb0ad5af35454", x"1826ab3543d94705", x"92bec775e45b5292", x"b4916f1f2f085a00", x"927159b8e23af622", x"d3c80d2e98c7762f", x"8e79c651e8ddc16e", x"b4a4469da5eff51b");
            when 25252673 => data <= (x"46d91554c7276e2d", x"0b7b3a41d030a1f4", x"463614984755ced7", x"94136f4f3ca0a668", x"430c85169c326abe", x"305fa51936aa408e", x"91b5e8ae61e06cdb", x"8290c544599a1cb1");
            when 17844244 => data <= (x"12421319bf4e3acf", x"d0cf511e22f8f482", x"889c1d038ddbd319", x"7cfd504c4e73a444", x"c9009e3e449e179c", x"a1b804bb6fa02834", x"b0f68b93505dd219", x"eedeb82c0b6c27e8");
            when 10966150 => data <= (x"4027d6f164faa472", x"40a56b7af9c0c804", x"305cceb31e05e34e", x"8ef503cc44b883a0", x"3615b6d05f90e646", x"678aa5b4212c866f", x"c5d7fb0815b37d14", x"e2667ae0ec24c265");
            when 6256103 => data <= (x"32aba5f5270f26e5", x"e0a1a1e7303ed29f", x"ef06d1ec2f1eb4a6", x"331fbac97f296097", x"2295ef0306363048", x"8a652f79a786abd3", x"15f56aad2d4f9541", x"fd94392942c4c611");
            when 30880642 => data <= (x"26a8eacf9bd60f37", x"5588ac6822a19e57", x"1b548fb2af8ce2a5", x"1b37bd76abb2686a", x"e89254677a36d2f2", x"45a06a8fdf701b79", x"9dc29b19ba644f8b", x"2663c67b879f1680");
            when 22305969 => data <= (x"1ba4b61f5a32cac5", x"05e49e2a3a955e3d", x"acd8cf36b67ecc1b", x"98e1c6b46cf6b4a5", x"e8252d813c6e938e", x"6966f27de091292c", x"52c4a796a795a3ec", x"49b90b66c1da6095");
            when 4532645 => data <= (x"f11b2400b50e27c0", x"0b9b36b7c15e8a1c", x"3ea16cb7f2845c9f", x"7f135accc8ba2dc2", x"fdc8707dda8bad93", x"9c555fcc05994753", x"012bbcd2d471b0e1", x"f161a66bcb41fba1");
            when 21678279 => data <= (x"5910223b0c70838f", x"3090422226c8910a", x"57e81513755e26a4", x"f05c804162e4142f", x"9ccc49e0cfe687c0", x"ee4cb4eaf0257938", x"e15b5e134a6086ec", x"434473693a6bfde3");
            when 17964764 => data <= (x"aa946e3dd448010a", x"390b8206ac807e6d", x"94f4bdbff2832da8", x"232beb936b433134", x"154faa469c74c418", x"f4478d21823bb069", x"de0c6881d9bdaabb", x"3f7b9b1b0f4765d0");
            when 24391780 => data <= (x"591b571e6778596a", x"6cf6dee1a28a0f43", x"3cd65b53dfe10600", x"6ca7d25cd88152f8", x"7cf9a36ad1c34895", x"16d44b04eccedd04", x"1e0ab7712f54942e", x"8552497759bb934e");
            when 15897664 => data <= (x"84d6317ec705d930", x"8eec52788f077407", x"cf09d5b01be70cf9", x"dd9a259c3864649d", x"3e5e8fb06f0813e2", x"51b8d499c90e1bf2", x"a288ca2c48f58dd0", x"b2a1dd0c2c2370df");
            when 2900508 => data <= (x"e9941f2ed60157fd", x"eda3ffba410d66f0", x"274e539a9dfaf058", x"8b5d6604921adaa8", x"a38ca06fee1d4adc", x"23919a6a92f98bab", x"b4c12329f19a464d", x"a2409f4795cb2819");
            when 33080761 => data <= (x"a6cbc7d1784e85cb", x"8a819455867e19e0", x"cf83079fc7350dad", x"78fa660f9024d23b", x"3f6b5077687d59b8", x"f6f1cb4704f65e54", x"41a9b39ed52efa84", x"e06abf901101b233");
            when 912509 => data <= (x"ef4dc00de1863f0d", x"92d98547a7389669", x"e20252c2933de495", x"a372315462fa54c2", x"d6abf46130c7f26b", x"cee50eb5b254fb0b", x"97d467fe0405ff67", x"a744681f259c0a74");
            when 13870088 => data <= (x"c5822360478889ec", x"e5806adfd6df2913", x"ced09037e4855413", x"5c0a68f74461fd79", x"f7b35c6febead29d", x"6f4370097aafbcbf", x"091eea6192bd0bf6", x"59b1c27e5ca75cbc");
            when 25479696 => data <= (x"1e8e6ada2ef6a614", x"ffbf512aba715f59", x"b70ed70c3d7e393c", x"5802c00dc3996fb9", x"48033f632be0fd4e", x"41da9748a2fa1b82", x"20a3b7ab3ebde4e0", x"1ee6126f93162f97");
            when 12943281 => data <= (x"d49eef5034c1ce9a", x"f7eb9ead161d3b1b", x"46d58abf3ef714a4", x"464fd129c2a8e949", x"fec67d1c2c0bdba2", x"7b9e1b06a17df35b", x"cc03a38718053e3b", x"2ff7ed54e71c51f9");
            when 25447029 => data <= (x"6d8bb68184739dae", x"bc1f099b28e72ea5", x"e319ac8434d9fe9c", x"b88b5ae8ee682785", x"fa4a3932bfe7a11a", x"35d23487addcd6f8", x"4cfb008ba8659a5b", x"912246f9bbc80b8e");
            when 9183869 => data <= (x"5d8df64252188c3f", x"a376fe8a024a63ce", x"33151890893409a2", x"071dd673074bad5d", x"b32d65a0603b27b8", x"61c8f143b504d87a", x"f6a907d22003aba9", x"4c17be7ccee52073");
            when 16497083 => data <= (x"9a210e4ad3f57bd3", x"09483bed6019215b", x"811471bb2e0e73c2", x"1c20626434c5e2db", x"ff20d9bca1c66bf0", x"ffab4ba5dd91dbf8", x"f124b15ef153d2e8", x"d377f9b1aac45301");
            when 32603069 => data <= (x"87662b9cb10e87d1", x"78618b123fddcb6d", x"c587fcaa9d5bd8ff", x"1f81ca93a102b6a4", x"e77c3662d006cf4e", x"9db6f43717d93f6f", x"cbe43fbedac3910e", x"cb55a2228be43b3d");
            when 27748643 => data <= (x"ef2b68af388100af", x"1a57ed7496c2b5d3", x"9af1ca29a46d5b70", x"11a758d862e58dc2", x"f41d840780d03d25", x"644f93e3db032962", x"d84e84b971ba994f", x"84ae3e3fc80d3287");
            when 25089355 => data <= (x"6a230cee03100e8a", x"434813217d3b54f9", x"5ebaadb51e60f06a", x"ada44fe8035738d0", x"09b461fc2b934ca7", x"d021a4e9753f6f9b", x"1ef83f1942b470df", x"d60b5e9bc339a045");
            when 20731187 => data <= (x"3ced2ea06b53fa41", x"b5b862b725becffe", x"20a717937ddac8aa", x"70f96b8c9db776f8", x"c2e12ec02ee88589", x"cbd7675280aa327a", x"57e5526c9b55203a", x"e670e6ad61b803bb");
            when 11545351 => data <= (x"32833371754d7af7", x"8b3d5b9a47506826", x"5d974375852b89ea", x"61ae70a7cacd257d", x"7ae40855158af8f0", x"1c4f8f61a83d7dea", x"a9fb386c8b1919e3", x"b9dc9ef2101084c6");
            when 11941929 => data <= (x"966f9d744cc4e6e0", x"2cfbdeffcdb832cc", x"03319abd37dc1492", x"27fa896548904e19", x"1209ad5d2436b44e", x"a26f4153a7bd9283", x"609e235ab5775c19", x"63443c20ad32545d");
            when 7887895 => data <= (x"e761d9f5657b625c", x"e9167283bfa0a724", x"d87719d186a1c45f", x"cd17a4d7524f389c", x"de4b6b537e89f9ce", x"75802e8e25d43d2f", x"35e024005b0c75f4", x"8572aade9463b23b");
            when 17406487 => data <= (x"c4260abb47ad4af2", x"76da8dbf6c40674c", x"1e17e42bfa1f69be", x"430410c17c2cdbdb", x"5eed80324e70d392", x"d111a5a4adfb93b8", x"7644cc05bd4be276", x"5556ab0a7cfc1966");
            when 1042889 => data <= (x"3f527ffde67d056c", x"5cfdb0dffda4ff52", x"0936e44b4c301bb6", x"b9d13687593910fb", x"3e072f603d6c5dcd", x"b72f938b02a2c128", x"1829b64a2643605a", x"7b3371e3f4232f6c");
            when 3044348 => data <= (x"2b24fbffdb79e981", x"d7a34da9c66ee54d", x"04d25a08334d578f", x"0dba14ea2e3c2bad", x"47ab70c2c750c9af", x"68f6ed6f68a7bcb7", x"edcf484f3ef4e956", x"5158871ab9171323");
            when 9889422 => data <= (x"50e4f37f83b19b4a", x"a88d8acf8f58a29c", x"96010f82be7a083a", x"2908b335b7fcec83", x"fa9d472a18ce11ed", x"88859d1604e74e26", x"71456efa4ff60c0b", x"d250d9d105dcdae0");
            when 22685700 => data <= (x"431844ecbf102cd2", x"af31ef91dbc95147", x"73dc08a98c6610a9", x"c0489453ed2d2a38", x"99719e8fcd0ac501", x"54385ed92997e88c", x"857bad399a8fe442", x"6484d0593db5c638");
            when 11926949 => data <= (x"9da7e37606920381", x"be8769c35e7bcf7e", x"bf62588e23c1cd7f", x"6da09560476b053b", x"18735c3407170dca", x"e36acb1954d7b72e", x"7f1e964c3b57abcb", x"55a315ec57950238");
            when 26286225 => data <= (x"75d08589b76190e0", x"6ed8208ccd82ce20", x"d5fc96846c976b45", x"5d6a3106a338d4e6", x"c002e7af0d95cccb", x"f40a75a1f0735be2", x"66e2c70f2285b997", x"b7f283378d98d8c4");
            when 5459273 => data <= (x"094031d6c4ae4d03", x"290ff0723975fd15", x"6bebf2e94f4601fe", x"fe04e822663b4507", x"cda7bfc958a5cc56", x"be0112d5dfd45f3b", x"7094b18b9108c693", x"d2ba7be47c6de042");
            when 25577418 => data <= (x"43d7a0c9a2c706db", x"cb1cb7bca998eb5e", x"a38fb4ad5e088dca", x"9edba8198cac7b35", x"00aa0c88a215b83f", x"6d5f9605c6ca4dba", x"f5db5f5b9c936a1f", x"e15c31bb840359ef");
            when 14679700 => data <= (x"7e891e6a134324da", x"a6c476a69bff4167", x"cebd7a783f963ce7", x"311fa0a348fd9892", x"b6a4169b5ad03dc3", x"e458506665c42656", x"99a64f9649a33c30", x"a05d6a55e9e918c9");
            when 13198834 => data <= (x"91881bc0d3c3e0e2", x"9dd9abbeb421906f", x"a5bdbdf5109ffb5c", x"2a6ccf1035db6b37", x"8f5128cbe046eb5f", x"a14e014be9775f03", x"35f75af5d5029a28", x"1ae7ec74f246dac5");
            when 10450861 => data <= (x"b81cc9bffbfc31dd", x"e7d5c427b28214e0", x"b69b2e89616d46c7", x"8ddb167997bdd935", x"337b5738f680b650", x"7a40dd8a6647fd9e", x"f313768caf81a196", x"0c72d91c64de9470");
            when 30652227 => data <= (x"c04d4c965422e992", x"b3332c232dc84ffd", x"c3d51bc2916567be", x"dba3060809c666b7", x"7a689676c30f485f", x"f4bd5eea59ee3205", x"eb805385ead37814", x"0333a1fe7316c281");
            when 16996130 => data <= (x"1545d11d2bad6efb", x"6382dfa486207d7c", x"b29c3d1c9120f154", x"4490b7ac90a93bc4", x"c035925950c143d4", x"3f1da9bcb0b23ba4", x"d11664b54bfa7ad5", x"cba4091b5b9976f8");
            when 23256480 => data <= (x"c6429fcc2027ea59", x"bd11b44a8afc745f", x"c66392183218432c", x"1c54707885d023bb", x"33899d18655d29d7", x"48823abb2798887b", x"abf5ae1ca2e7fe19", x"9193295bc86f787e");
            when 1641757 => data <= (x"a06f9308d9f68d7e", x"a00eeaae9ff6c606", x"343cb7c2d300a35f", x"bdf36cced38cf1b5", x"b15b5f39efdec45f", x"a046590db8681c9b", x"f581f7d179be0787", x"8fa175c03ad61603");
            when 10374150 => data <= (x"b2272927796b40f2", x"6c4cdf89715a81b7", x"e3a3318414fec531", x"e41f86118795f10e", x"8d5789fe63a75f45", x"d07474ed4244973c", x"eb051ac8cbc41957", x"43fbb9c9d6eea2a1");
            when 4469239 => data <= (x"6d3e56b883246634", x"9ba8653fe020e29b", x"e58d7ad9f55e993f", x"6738de7827b01943", x"becf83740201fc20", x"3809b2c5c113eb71", x"c2109d25b1fe7e64", x"d74b930097c72ac2");
            when 15815556 => data <= (x"09da6dc4e95142c1", x"f093bc135642926b", x"aa49dedfda28b13a", x"9a5de8f70eadf099", x"96553b8c7461ed1a", x"61acee9231a1350b", x"b547ce9ed183a756", x"6f283a922c97b8ca");
            when 24475981 => data <= (x"01922db794e4b87c", x"23cf01d622b47de3", x"839c46cd87efba13", x"2acda62b71438c98", x"5ce64e3d62bac47a", x"259a54662e015470", x"efd76480ce6dc93d", x"3a641e0884b6b000");
            when 13430113 => data <= (x"55d05503dfaeee94", x"23ca49a88136ad08", x"fe7f33f730c9cc0d", x"117fe6a2f4d0a618", x"1b677aaa89be0fba", x"f5e487922de17cf9", x"756b3828fa544047", x"99f7a516e84ab3bb");
            when 24044666 => data <= (x"09258737ff809691", x"d214f2ab8c7bdf9d", x"518f60030110bf98", x"104f7e10b03e9ebf", x"b9a44701d76431f4", x"b6bcb950669d1498", x"527ce649f452964c", x"00985c0a19920a7f");
            when 2979777 => data <= (x"3ef64c3968e1edea", x"cb678591705a8197", x"45150adfed0f2954", x"74bd6d148abcebce", x"15a4ea161ab5fd8b", x"d5ff8c9ff4115930", x"fd446413c8277d52", x"481955bac5cc8ed0");
            when 17225409 => data <= (x"0d4e7dacd98e4625", x"0010ccdb667e3383", x"a1705c4d71d00ac5", x"8642a5d1e1a8d2e0", x"f22ec2cbbc56cc3e", x"dfd5dbe2d3a27d86", x"deac8f82341f13e7", x"8c8c8a8c198f1f4c");
            when 32244856 => data <= (x"83f9f18337072bee", x"44c7f0a23ca8dbe0", x"7bec2bcbaa13b670", x"f50e50d604ad8bce", x"c573a09fb93e3499", x"538bd6cbaa2635ca", x"7956be66f709deb8", x"a348bb6f844e38ee");
            when 22106746 => data <= (x"6c32f5f9335190d0", x"84d3b934707a3f42", x"0609013948ef8a35", x"e17090d1702fe4dc", x"26e1a702f82e0174", x"7de63b83eecd92a3", x"5b7ee0e8cf2f3ae5", x"fe026f15d71b3bf5");
            when 29963834 => data <= (x"1ab6753e125010a0", x"2f8d6f7d4a348d03", x"d79953a2ce22790d", x"f58500614c5bd18b", x"729a97a558fb7548", x"1dd43cdd304d5ccb", x"1a39dfa692b045b8", x"a94ea60f2cba33e9");
            when 18952654 => data <= (x"8c90bb6caaac57b3", x"79723fb2f9c85ccb", x"f300a6848aea4657", x"72579dd55db8947b", x"567f5c6aceacc2f4", x"0520e0e090d1efbd", x"dedb38e5183edbae", x"a09313e1da1b3e68");
            when 4269832 => data <= (x"8085c1a6f1af64a9", x"5f92520ff6e781a8", x"7c1abd4718f5e9ad", x"cb5a46955e871e7f", x"64aea27540034868", x"a8a550def4099506", x"aa40c80a1035571a", x"a6cd7c706ea8aeab");
            when 10564763 => data <= (x"a3eb49dfe73cf911", x"3f4b82e5a83cd33e", x"84811555a765f3d8", x"c5a5dcc0e501d550", x"fca31e59ed4ec1fc", x"c594b19f6b8b88db", x"828a63f5fb8b4423", x"21b2ded28f62e8ce");
            when 7695367 => data <= (x"8f049443b4832f1f", x"869afedd3d361b5f", x"f5d6349553eb61c6", x"422d69c0e4b5dac2", x"38e31c5593252f8f", x"993758c741a914ff", x"bd4f7930b792e16e", x"b78fc3be152de7d4");
            when 1219337 => data <= (x"7dc14eb17199cb2b", x"d0fa9bdc7972575d", x"c302046a72c3479c", x"33e6a0edb5d0a051", x"df39258f0113221f", x"4919c9f9e035cc15", x"0857c779e28cb0c7", x"46b79ed1d4f44f79");
            when 22486681 => data <= (x"7eba751968d5028e", x"5509e0dad2e8fa3b", x"236942536329c95c", x"827b4337e84384e0", x"1f8c488ce944db1b", x"0de731e9a2a5d68c", x"016fa1bc284c7521", x"cf176339c3ae5738");
            when 5387573 => data <= (x"d0751ee8baa504bb", x"4284175a8c245a91", x"d6f37d16e63abc9e", x"2f8dc3ba28cd9c16", x"9a473f923799226e", x"79093099e1e4c785", x"ffb75c536cc70e0b", x"7c1f59fab0bcf1e4");
            when 21797363 => data <= (x"75fc4517dcf7b351", x"06de534b2080b121", x"3e1aa4a463a659b5", x"0c246b5776ff739e", x"37c17ef783813451", x"6a2208ec742fc7a3", x"66ced635a7f9ec35", x"eebe48fdcfc5db30");
            when 1002202 => data <= (x"e4dd7fc7b1a7d56d", x"c443f3252bc80d43", x"03138bc8249ddee3", x"3a42c2c85dd70c35", x"86e36c741ba45da8", x"a5892bc08d8d4170", x"bd4be7a3e780dce0", x"e19ba10befc60ecc");
            when 10063842 => data <= (x"92e743edcd486352", x"02f65800a7b52c73", x"78565e8cb8e5cbf4", x"79cd8a401b7cf27d", x"71fc4aaf9b8bb661", x"9bc347c0fd60169c", x"affc15ed97dcfb42", x"22779088687db5d7");
            when 11402630 => data <= (x"3571801a3fc085a5", x"b612ad4c8a6c7a2c", x"214eaf5ffe2bce46", x"1298e8e1f62c8cfb", x"768b27bbab8672f7", x"7519ddd714b03cfe", x"9f9153ca98333844", x"33239c99b9e4c17b");
            when 22920609 => data <= (x"129a19425466d527", x"1c60531fa2a405d9", x"684844a19d10d498", x"4956913be6382bda", x"b7882a22e6e8b9f4", x"e3cc8468d779ea2d", x"ab210feff44f10a8", x"6b2aad243fc7909d");
            when 13086625 => data <= (x"83813856232f9469", x"a56bd4c283be55f7", x"98739995f06165b3", x"685aa7057a7862d2", x"d7a78829db51f05e", x"a8d668ae04bc036b", x"ea520dd42689d054", x"6e209f7fdf1adaa3");
            when 18428816 => data <= (x"a6841b677d5c454b", x"35008ed9394ab305", x"cf2600f75c9d3045", x"1903b40b71a045f4", x"c6270170a5d39b5c", x"73f8a5ce54bd1afa", x"da13493ecd220ab1", x"d5a4bcfef8907230");
            when 33356417 => data <= (x"8c8015cdba3bb50f", x"e32b58a6f7b317a9", x"169e11a773e5f0c6", x"a90af88a9479c527", x"4d82883cf56d674e", x"bd448d7d934949d7", x"b7cd7d6dadf752dd", x"e3451578011c2c55");
            when 9697414 => data <= (x"a9af040a49983e62", x"a917a6777e8c1a45", x"80cfc13a6724cff6", x"ea62e6facbca051e", x"bd847bd88b25aa9c", x"1468ce8ec55ac0d7", x"e3bdd65cf3453c6d", x"be592f3bd308d483");
            when 17634874 => data <= (x"8d017a5337472040", x"e2e6f9bde1119fa2", x"fd6dea273655546c", x"fb1a5a7fe2b5beb0", x"8fb8cd03b53b3fdc", x"ba6ad7d312761a86", x"0b9f1508c3f35fbc", x"7c7500a054782e45");
            when 5386856 => data <= (x"ce48e6c688c25b08", x"2f72178311e4d9fd", x"6fc4d688d084208a", x"769cdb890fc2714f", x"125b9333cd7ae847", x"5ffc499c152bdb2b", x"695714512835cfd9", x"37d3198c44760e1c");
            when 21153858 => data <= (x"b10132d4fef4d8a2", x"df5a4ea6a21f7348", x"4442469886c095d3", x"b4a78e0f6d80b429", x"deb1de7d7388c448", x"a39964cdfbe64f1b", x"a77b449cd1f93c4c", x"0266fb841b229bfa");
            when 7426573 => data <= (x"359890d3fe35c2dc", x"aa3ca8d0a45428a2", x"57d665b30540f600", x"859a68053c90b829", x"70f03e9fa1689cfb", x"a862f406aa66d09e", x"c379ae0ad08c2dc1", x"be9c5310acc38498");
            when 17584598 => data <= (x"3d124c2e64b1f293", x"f09938489179ef3b", x"b4ecfda0eea7def5", x"8afb0da61f19471b", x"74f4d2d8142d9afd", x"bbd00bdb8f7ce856", x"80d705da9bd7f7a0", x"b44180c06660e29e");
            when 9729799 => data <= (x"4cf975186e51c7a5", x"6b100e2613f10dc2", x"24b30202123af217", x"b8b1ab1db3034595", x"a744660b8ec3da22", x"a2e12ff1372521dd", x"75a14d6b7deff879", x"9f9307694886830c");
            when 566626 => data <= (x"be8d31703dab6541", x"9ff0efacfe91c710", x"2ddcc03071ef73d1", x"5e6cdba59cc35c12", x"5b5a39036c5b0ed3", x"7e4c7e22abc5aa3d", x"bc93fd1c41de0db3", x"c52f1822af218560");
            when 25352179 => data <= (x"5690e9cdf31a9be4", x"5a2179c04367f6e1", x"a4ba12c78869481a", x"b79ef8a1ca224eb2", x"7a875a6ce50edf3c", x"697ee542cc6ff9d3", x"aa1493c4b2a19420", x"dfcc3dc93656c1cb");
            when 6453029 => data <= (x"9dee7a01a7b45721", x"4c552b38b22ad063", x"2745e6219dbb3a4d", x"56de0db698ec510d", x"2503b0d91f228210", x"20d0a732406ea558", x"4f38b99feee6584b", x"c6a72839b5239334");
            when 9642528 => data <= (x"9d83410b889a392e", x"7c796211a3690a82", x"dfaefed7a0f423d6", x"c441fc9962eb4ee7", x"d0e886c5ac6ddbeb", x"26426cb2cfc07db4", x"dda9cd176ca86386", x"07c45ad89f1dbf0a");
            when 32894219 => data <= (x"915aa496b04f83d8", x"c63224531cdd1a14", x"b8dbe165355cc2c5", x"625c8c188a786ea8", x"fd107b584356c135", x"d6bf199300ca32d9", x"89f25b214749bad1", x"5737df55aa70eb55");
            when 20562674 => data <= (x"6eaa71f3e215281a", x"f5395be036d95f26", x"081f6a106e50dd0d", x"4ad079693de4d129", x"aa77e9dc3253a71f", x"46ca6d346553df36", x"74fa7ca5af2aef23", x"4ee44da91b3e4e57");
            when 29821649 => data <= (x"f6c535a8b70b8259", x"39bb6ebb4fe5ffa0", x"be5ef8c155d4dec9", x"30d45b0665536aeb", x"63a848d8a75580e6", x"f2667ac4a15f9a95", x"0273a70cb3c76a88", x"ee68bf3f470ed90d");
            when 33408912 => data <= (x"60703c60cf8ae118", x"8e7c0f2ba699fccd", x"efefaddd29ec5fb0", x"812632a6b852a330", x"58869b2809ffe277", x"263c204e23196f5e", x"573a680e5ef2836f", x"6e3eebd4fec808e9");
            when 25980112 => data <= (x"f3e94528400668e3", x"c9a30c7c7d2970f9", x"9703edaed7ae594c", x"b76ca65d42155257", x"919fd1599e199ecb", x"5218471a31ae5f83", x"fe1b9ad46f8704ed", x"438e922a98187f7e");
            when 31053656 => data <= (x"0be85c10e6351c31", x"4eab3814a61d2b52", x"b654b3fca19c8e9a", x"1583e19f9d58f8bd", x"e5cba7f2f5751384", x"bda3117121cc3a6b", x"bbb08e48a14c312d", x"9701771ef86e06d3");
            when 25620255 => data <= (x"6ed6406c36b22283", x"82a2d7119af0cec9", x"0962cc596ff124e1", x"0c20193aa190fd23", x"5e3f1525101be542", x"5901737ca4c70455", x"59887bd6cf64c827", x"f03e09fd6ec3974b");
            when 1686678 => data <= (x"0aeb3bec8ca2b4dc", x"81a3546d111d4a08", x"dc137fd6d747eda0", x"07068327229de6b1", x"9e6a40624d0883d8", x"92fbfbdd78595d64", x"67ba4f52b9c99acf", x"1d1e7c5657685c4e");
            when 19080233 => data <= (x"68e401d8451d798e", x"3b6fe92983a11271", x"3ea7608328b5fd78", x"c9b0679f6f77f619", x"542521d7ecbd682e", x"dbcb9bb4c695ac34", x"6a1cb45ed2a9540f", x"a14f8d3d61e0fde1");
            when 27055284 => data <= (x"c95023d7263cbc0a", x"ff0c755f8245111c", x"627509e119a02b8f", x"15027240424851a3", x"8b769f2d9550f137", x"b1eeb015cda1dab2", x"53afd9f2b4177b65", x"45b79b6cbf17ed07");
            when 19240760 => data <= (x"b17c1146e37454f0", x"5692b0b87c36cb1d", x"2f584945a84e2ad8", x"2146e4d55570fba5", x"ab884cc600d4895f", x"15607100af41606e", x"86b1c2b2d21ff23d", x"52c8002db8176aea");
            when 12861955 => data <= (x"a21b2853caddf15f", x"ea9fc0c948fb2da5", x"48c56bd46a50bb18", x"f8e8b2a16d6597c1", x"dd3b9219eb9c4b33", x"1c130ffbca3b42bb", x"de0ee7d8e6850eaa", x"5fe1b3be33369693");
            when 23301756 => data <= (x"289602dc917a5b97", x"2838746bae5b6b68", x"c89fae9ddc3c5f6c", x"dd0308cf1234a24a", x"8ad0022082c8f442", x"bf9852429e709e0c", x"44b345bca8f4805e", x"b551394f32c3e6f0");
            when 27821979 => data <= (x"129207745be204e2", x"7268b5abb89f4d2f", x"63b234a96592f443", x"7496a2d44f62b27b", x"947a0329d12b30ba", x"47c0f2a018eb8f29", x"ea7efc7debe2d2eb", x"50c8db7e80578a0c");
            when 30545943 => data <= (x"0de573447ec2d550", x"cbac1dbbe60d5ad9", x"503d468814d6686f", x"9fa0a740b48b3ece", x"001bc86c569f240a", x"a413f67695737811", x"f3f3c6325693ed25", x"d506516d438bad72");
            when 12812855 => data <= (x"5a3c00f07e0c75f7", x"f7b5969cb1578183", x"ffab9619e9d2108c", x"457763dd928d48fe", x"961d7b329b11d624", x"ed398e3e7ddc5da5", x"4138c83f2b57bfda", x"35213b823a5b3bc6");
            when 9822177 => data <= (x"6e12667e2ca8eeb6", x"541ae2e479230c56", x"9de5b4cf575ededd", x"cb0f26b16e5155f2", x"ee37c81d9bf770cd", x"1e196a2c6a923744", x"ebbb68c262c53b39", x"c8e78b772506a82e");
            when 7102454 => data <= (x"46f2285ea664bbb4", x"9d51fc38f015f78e", x"80363655473fe0dd", x"45f707e9a5174944", x"787016d6fdf130c1", x"f62628ae67b60fa7", x"007bf92971420303", x"b3eb14681186c430");
            when 18458765 => data <= (x"f0aa1baedbae3a8c", x"c461e60818ea0164", x"4a9b97c067915819", x"2f3166326b28aa5f", x"b58ccefaf79f28b2", x"c90a128428a60c5a", x"85c13de7b6d4f5ab", x"ea344474bbb9d8a2");
            when 864555 => data <= (x"f2252b10a2617217", x"4665102874e23660", x"5f1fae48e82f2ab5", x"759cd6816e20fba7", x"84e8a25195febb63", x"691b0145bd627477", x"eae98101243f137d", x"23f38100cc7cac28");
            when 28504211 => data <= (x"eacaba2850f44ba8", x"37ba811aaa8ce167", x"82d3fb11af7f0d83", x"f556896919393cf1", x"5d2fc4989c6d0ba4", x"76c2334d0d3fee89", x"c2f67396b391786a", x"0a899ee4bf0ad31e");
            when 3793264 => data <= (x"af7714f155b81d58", x"31f2fc814cccf031", x"cd5c064051edbe7d", x"38cad9ffe5dc1953", x"a93a39060c179517", x"2f6b8f1f8c67d869", x"c7c674ef0adf7a57", x"0a8eb1b9f9545df5");
            when 7858594 => data <= (x"a7507386e57968c0", x"73085da9e7565fdb", x"7bcbf683148e6b35", x"2fb179ee25c7d624", x"56601848f7a46f5d", x"1ff46db02728d816", x"fba67fcdb83430ca", x"198f09b01af5bed4");
            when 6734674 => data <= (x"73000297b35288f9", x"6c3522f0bd957c06", x"64d720dd484a49a8", x"cc92e9a8c1e9a158", x"56cbdc22741437f0", x"7931817fd24bf9f2", x"a1496f7423b591c9", x"7eb71dea8c75e518");
            when 790797 => data <= (x"3c80281f7bce63bb", x"fec49ee9406ce714", x"5f206362095f8791", x"f52069ea508852b8", x"0e789b645f37fe86", x"398120ac747f6baf", x"2238645c7ed103b4", x"c1ca3d3cc3aa538f");
            when 26057200 => data <= (x"304a6af96262ae53", x"0e935c1efaf66ac8", x"bca10bb31e27a9a2", x"94dbd87a5b076e5a", x"8c13407e4ff68d4b", x"53940ed3c5de9079", x"87f44bcf323c5eb4", x"0cf4059a24d56ed1");
            when 29790933 => data <= (x"27ab40ef5f837803", x"2e5269e303dace36", x"0f05f46b84af7e60", x"50901b9a8ba2e570", x"61520384be2ded4d", x"864fced456bfb50f", x"06051475a5f8cbe3", x"2ed7866dbe63d928");
            when 23450905 => data <= (x"ba69b20063f8fcd6", x"84c03f8d8b84d853", x"58dbd27ad137c6ba", x"341dae807b68e7fa", x"bf07b9bac65d603c", x"e2a7e94df9935f85", x"4320fc3b0195dc7d", x"b8df0ccac7bc2c58");
            when 18809703 => data <= (x"a641ba770b830aea", x"0b9d6567f381e2a2", x"7dd0c39a26ab728e", x"7ad608d5c443c5c4", x"04c88fd696819a27", x"5622efe001a3c2fd", x"2de3484331629548", x"599f0a6fcd89de57");
            when 11617309 => data <= (x"d2c01a9802f6fdf8", x"cb9d2bbd6005ee2b", x"4b62f15418c69f3d", x"5f3a599020017936", x"572382f1bce32164", x"4fdf39d826d20c32", x"1b215b33cddcbba9", x"a09118f0b4d8588b");
            when 16065196 => data <= (x"8199d65f9b1d7cdd", x"966b88954650364d", x"da6b7a489549e4cb", x"91190dc927aa9bc1", x"dca1c028d5c5e588", x"bd33d2bdecda66e7", x"1a5c8b16fbcbb059", x"4ec01f23e7eea962");
            when 31474634 => data <= (x"287862579e2cdac0", x"8ed027bc367ad1ac", x"19b65642602508fd", x"4c591d4b996b1e76", x"1410883b7d94b543", x"c21dae6730447547", x"30c56f708bfd152e", x"8a8cb3051501b5c6");
            when 18750547 => data <= (x"03ea1d82e5f6b1b7", x"36425c53d1a4d94c", x"d10073f26c225728", x"5ae29ea31ef31847", x"0426f1e62feab33c", x"e2f44b54dc2ab397", x"4bea3ad606281584", x"c1436aa468c90f8b");
            when 21161231 => data <= (x"b01aeb389d917dfc", x"13b66e920065c7b4", x"01be7b22e6f6ab07", x"ea287ab955318847", x"3a47bbd1a09ce88e", x"fb4ff59be81a6986", x"22ce1e1683f2abf9", x"574fade0e274eaa4");
            when 30304302 => data <= (x"217998bc3045104c", x"da57d740718f6b21", x"6d98b49afbbe5014", x"72ad9420e5778984", x"d72f28bb3260c08e", x"3e725ebf1dd44ba3", x"1ed4e6802fe66bfa", x"85cab656ef31cb28");
            when 20936432 => data <= (x"220c887a5bbd8863", x"f48c6d7c0cbcbc87", x"b482b540bf55e09d", x"130cfb931cdb293e", x"443fae59abdfe990", x"6b019d1a3a0f5427", x"f0c414b3dac444c6", x"17f42442eed2cd86");
            when 27789779 => data <= (x"9b86ba387fb8c62d", x"ec438e49ab1d9f0e", x"010f83e8503c3634", x"fabdf30d89bce16f", x"2efad3f76567334c", x"c6b304a59dd3b5e2", x"f22b878116ce45ab", x"bef8bb8ec6e0d0c5");
            when 1219834 => data <= (x"28675134997cc561", x"ef66a3f1c65cf441", x"f609c7c176caff18", x"1c6aa6b39c1d69b5", x"46a7abeac88a6472", x"da48f0399cbced69", x"1f8b226f3c1fd32d", x"29b211b0a4b4e025");
            when 16757007 => data <= (x"fbc8d1dfe923b927", x"e01d24fd90eea494", x"c1e417eb36cdfcf7", x"cace7a87966457b1", x"e3a73492ef1a4aba", x"c92ce40750e0b3e0", x"6de8072ccce784be", x"779b9356f327bb54");
            when 33744300 => data <= (x"2806d1309f1fea0d", x"772f283dcc05842f", x"de234cb8f40ed926", x"f3e82c7fb05babaa", x"fd00a33e1a407216", x"1c249c8da036c46f", x"6953b5edec31299c", x"a3d3858d8f19ceb6");
            when 955127 => data <= (x"bd6cc4c077bde68a", x"474018ba6b57f908", x"e612247da8409e9c", x"28b38978ccdb60e4", x"b7d12bac3600abcc", x"78a239ad310a2c20", x"be13680b86aaf590", x"282bef58b2dfb31f");
            when 23996749 => data <= (x"8efeed0459992d5f", x"38cf70e79e8d0ba5", x"34e29eb420c1d123", x"deeea0d7fee3a574", x"070e477374811e9f", x"e85fd754919ae0fb", x"0328bd0092266271", x"ea273b2a60b88c84");
            when 17658040 => data <= (x"ba41ef8aa7e79225", x"3a73bba5b5ec36f0", x"9703f7282591efe7", x"d77927b2104f7058", x"fba425d2332d8aeb", x"1c349e1c622df218", x"cf2ce4f9526a3cba", x"0a6d8200d70eb8b0");
            when 6696889 => data <= (x"0cd16e6763328234", x"158264cb9a018a4b", x"78b14a38fab5be42", x"9b4966fc336e1e73", x"5a8e391fb0d8383c", x"0311791766b63b4a", x"02f1d7a4ea590811", x"91275ff1d9d01899");
            when 3691036 => data <= (x"9975a5c6c358bd3b", x"e2f9ee91880a9843", x"9f4ff0f2ae042608", x"ec05905b27e5519b", x"1a2d19b151d2eb03", x"facac4480cb5a2d8", x"cc28b78d43b91fce", x"580238fbc1fd0ee5");
            when 10974956 => data <= (x"afe3cb3aa1c8c4af", x"863b6c26081301f2", x"822fef5e4e286661", x"5df9d0debd227f1f", x"b11c5620bcbce7e5", x"939b6a0133d9b0c9", x"e62bb28b11289631", x"1efba81f8e1c4215");
            when 22470755 => data <= (x"449f7c6b83e61715", x"3769dd4cd03f923e", x"3561a730734c76b4", x"388d42d6f2955b71", x"7bca4dfdebc3c279", x"11b37eddf74a711b", x"7188882a7f0bf191", x"a9e98b7eb3ddc9ca");
            when 6294722 => data <= (x"cf407d276f4412f9", x"691aa9d164559854", x"43e8088920aeb613", x"b618c34fea1e67b3", x"132faa9d379f7bbc", x"7eede3273d779ae6", x"405a511ab779d70e", x"052c61c1a07f8e52");
            when 2350852 => data <= (x"a2ff1a24266e3f37", x"28222667dd727f10", x"3b275e0fccc5aac9", x"b0b2b77ef0e5d1cb", x"e9b1dac46c8bdc96", x"f37144d99b7e94ee", x"e575b2f61f4d0e68", x"5e618a5c3785d6f3");
            when 10731103 => data <= (x"e87f006ae1277de6", x"558f9eb78e1afc98", x"57f65be4c27c5d4b", x"0eca5932f82d9954", x"a7a617304d4d2719", x"3c504ef5a76dfaf8", x"1685a0cbda9531e7", x"3485ae9a059e378a");
            when 22985352 => data <= (x"bc7284a80f885b7f", x"e9e99f7ec797f9c2", x"7ce521f86b7de1f5", x"fcc63f6d4bcd0a74", x"148efb9328ccf437", x"3142bd9841bf19d5", x"b71fc3f9ee4b2e08", x"63e7d6f1dbdb5bca");
            when 5902918 => data <= (x"32384583651a0605", x"05585733e4c6838f", x"a9f715e14034d826", x"794e846050fdb9a1", x"b1dfc54207d29038", x"68ef262e5f1fc36b", x"be13e397a68379a5", x"faa2e930d2005314");
            when 18460146 => data <= (x"4d765250e56e0ef0", x"7b178660e607e1f7", x"68e2b817679acbaa", x"0ad420b9b78f13c5", x"8f143704f8c5de0c", x"11813940ffa45431", x"834d8aaf8c3f83b7", x"d347ffd8670d67f1");
            when 31181754 => data <= (x"75a48c45f3615d52", x"f03a6757f2a071d9", x"dc131ae312f52fc3", x"11b07a29359aad18", x"24f0917054495f3b", x"119b79d45347ac7d", x"795ae0ab1a503ba2", x"fd90936ce7167732");
            when 6055808 => data <= (x"1a5bc7df5aac9460", x"7fe17698fe9b6328", x"c5b31e5b2fa59262", x"4ae020daef3db00a", x"ebfd2250fcb00999", x"7bc918d3aa403207", x"8b132c0817ebc3f9", x"6c38a61ec91888b2");
            when 32204390 => data <= (x"55dc44b791a9a919", x"05fea4e3edf6d94d", x"d05006ca88321a8f", x"07f6a0a3813282e8", x"58f87022335133bb", x"a16d9a0737adde3b", x"153b2aea86879448", x"89ff713859a4408e");
            when 25319501 => data <= (x"0661792db9e0abab", x"62b9a23c8f2e0b68", x"887defed8b0e4395", x"34433775141ff4e2", x"dcb4316052459417", x"dc828879d6279ddf", x"451e63c423bab88f", x"5685f1d10b50ba03");
            when 29221254 => data <= (x"ea7281660473e518", x"a6f9f6f0e63f7357", x"6eba75221ea798b1", x"e72138d0d8d99609", x"9d57ed4d4a2f4eff", x"6fd7ce356cf366e3", x"72b2b073457fc904", x"b84c3d1d2ac62feb");
            when 26617604 => data <= (x"7aaa71af636d3fe2", x"b602f14a7a7a435a", x"43890c568144e18e", x"9f40c9d62bca459e", x"00dffe0e1c08459a", x"f3d604fbbd1f9f04", x"583b6031b16dbb5c", x"fb43a51a142a3012");
            when 25909574 => data <= (x"acf4df4dfcce455d", x"fbc13f61aadab60e", x"cbf54d9d63309b7b", x"6f366048a207e22e", x"d496ce1b8523d46d", x"486699af79c013e6", x"03160d8288414297", x"5847fd4c73548e87");
            when 32341611 => data <= (x"00d9b8a4410dd385", x"feb399a24d2d6dd7", x"2ca60cf04b1b45cd", x"297ba16e5664c502", x"e42668db289d6fac", x"cbcbf25613f80263", x"6024d11422544a8f", x"fcd35182b2e53c90");
            when 32522160 => data <= (x"27ecbe66a0d7131e", x"e220c478f420c223", x"dcfcb2ba7a9a2bc2", x"a2eb9492f00d25a7", x"4f4aa959a59f8b9a", x"fb67abe73ed54b18", x"0d89db8a38640388", x"ee7b6d301a3b158d");
            when 3212822 => data <= (x"673bd507da6fbdc4", x"8dd8d95c46665c37", x"ff9cc6435c2a1928", x"7f8f2f80d053af34", x"f8e715c806ab5dea", x"42be2ec5211aa2d1", x"c324b10404291d28", x"4f5cc7a38168bd9b");
            when 19419565 => data <= (x"5c89d07af90de5e2", x"e54a0910eed49636", x"ea7048610ab2dd8b", x"76b8535badc9a0dc", x"80a7e95e63e1c104", x"74c92b3a3fdd648d", x"591dbf79936d972b", x"e519bc4cd02151f4");
            when 29271533 => data <= (x"f7cdb074afc561f9", x"f79b6acacde1aefa", x"0ef633910769e895", x"da00d3c31e79f83d", x"b63644dab916b7d3", x"d362f408a2feb5db", x"61abe17ff2043bfa", x"b4ab21b79035f32f");
            when 21751851 => data <= (x"21ba76334a74d749", x"8b373d34e99481ba", x"e4969f0d02bcaf74", x"cd9e0596ea200852", x"e4f9974c8433b96b", x"fb0de547c307d57b", x"3bd51f9823f821c2", x"42a022122977b68f");
            when 31882098 => data <= (x"e62a23745b7a2372", x"cba0f5eaf28e2e7f", x"8e7f82b689ef42e5", x"7499fb2e833d545d", x"b3bc926a6c18a4a1", x"79c58b9cfed1dfef", x"d89698383dcb2b1f", x"fa85c0e783ec8b2b");
            when 21677605 => data <= (x"afa6438cbc0481cd", x"48f5f355f02f50ce", x"33408344c6f18a20", x"13d2f4cef34bb36e", x"05e419447a223f49", x"8b73885c671566c9", x"4e2eef4c61758d25", x"11f19de3741277bc");
            when 3964589 => data <= (x"462d85c998fa111c", x"d782b1f8adfb431b", x"ce06223d2687a694", x"24960d6a8e450039", x"4f7d8e4771f996dc", x"f4176a280e33a396", x"25172237d88aaa1c", x"461d4343ed10e980");
            when 24153329 => data <= (x"e70ce9099cd08f00", x"5ce515ca0792773d", x"f181a95806a75127", x"e0533db94901770b", x"492ae1ed19fd1ab6", x"5b9d3da0ac4f5554", x"fd3e3c598940a0c5", x"0c72e9ca41a17c50");
            when 29464814 => data <= (x"d692c827c27f7368", x"d6c1fad8fbaffee4", x"f668c2204cfe242a", x"435f224224126fd2", x"3e16c24b4bdf3ccc", x"631b73cfbb812083", x"096d45be773b6335", x"354fdf664949d7d2");
            when 17040150 => data <= (x"dbd0a1d7d9c52a39", x"f6658c7dc45227dc", x"ac51f6c9e5906b9a", x"888bd525cf9a203e", x"6356e8233d74823d", x"e4eead2e59890faa", x"4203d65e4dce71b9", x"35e1ef30b278fa65");
            when 8041873 => data <= (x"e689fd8cb76a4ce3", x"c003ee24bfb32ff9", x"5a7138f4e1958f77", x"f0c07b792b225b4a", x"0ad2484aead19892", x"35771f02000c4314", x"be7c95c961864e8f", x"a55cc464221d79e7");
            when 12531970 => data <= (x"2d5d1791d5a5eb40", x"d5d6be1bb21452d7", x"a80b211a88324808", x"7c1d437064af89b5", x"1dc19c693ef1ebd0", x"1b715b9fc6ca186d", x"cb4a93e5a9116829", x"61bc13e31b701242");
            when 26515586 => data <= (x"29b8e5870582d295", x"f2c8e8e43e9813f0", x"5af1dddf12b54261", x"64cd80a42d0099c5", x"6b88a68d74bbbc03", x"fd9075a0cdeb50ae", x"22e0a74ecf626481", x"5446b6ed7ce0b076");
            when 9365672 => data <= (x"3d1f4b7717ed84a4", x"042207ea6333e1ae", x"eff943933c486661", x"ab4220d2f9491bf4", x"79049e52ac54977e", x"0fc9bcf3bcc62533", x"01d25eacd10a972d", x"6475be5b2c175703");
            when 15464338 => data <= (x"8fd6da7d0855d609", x"66e513f75a62adb3", x"45ef5f667210e629", x"f9a5fd8848511fbb", x"0c939841ae0c9b3e", x"49f03069e1c6f579", x"ad472cbd89d2c76d", x"3f42174c5a7c2a9d");
            when 25263723 => data <= (x"c165414daea8b4b9", x"c1fd524ed24dff0a", x"9518b42de6752108", x"6cfc32f31a08286e", x"aca89f29d76f7051", x"8f39d83d9d06b1b0", x"91ce6fc7fd25d595", x"dedc03167929d376");
            when 13327481 => data <= (x"22d5b6d43d4c4a9a", x"834d8038084f0cda", x"b35fa39585737e23", x"3d4ce0bd09e456be", x"290a19c1ad8bf29c", x"40bf4b1d755cd66f", x"9554fb5927a6d23e", x"dc35ee0ba2d1d3fc");
            when 33316486 => data <= (x"cdafb5455d918768", x"24ca18b3254cb66d", x"d0fb4d98a6c791c9", x"d5db846a881faeb9", x"70f200c4f822924e", x"287a8cb3285595f3", x"6aef7603b75db162", x"c034c1958aa4a52f");
            when 32481660 => data <= (x"ddfe5bc4cd3ca9e5", x"7c271cc4cd1de224", x"7b7a9e7bd7f806f8", x"ff8fc98f8c78801d", x"a2320a6d88e6caef", x"405089769a4274a4", x"1f7009d8e68ba3bb", x"a0678acd6f227cba");
            when 26706043 => data <= (x"00593041737b6760", x"c88e4880a45a2c23", x"860af33a7d72a645", x"252356bdd8fc60a6", x"2849e485409f1abf", x"0c6a3aa0ef367526", x"24f361aebfbd4086", x"a70e18cc426d28f6");
            when 12680426 => data <= (x"eebc2c005aecd9ac", x"1219286e68e95100", x"c40526aa15ca23bb", x"0501ac19d76c4a3e", x"ecba911a1166f79e", x"dd93ee333907a382", x"f36ef0e4a32d23bf", x"f4909a4ba5cda863");
            when 23788447 => data <= (x"475a66a85e29c106", x"255fcc904c354b22", x"5000e3496cc3d570", x"09ac4fc102900e18", x"372109e877249b47", x"72dadd25352783e7", x"56ee4f37de6b5bfe", x"b7cc65f9ed5470e8");
            when 22587295 => data <= (x"a55b4e6a6bf17ec1", x"dbca5091b619bda7", x"dc1110d0c378771a", x"c8d61dfb73b55201", x"c60af2133d0731d8", x"ffa6dcb66226c992", x"023cd3f798a0fbbf", x"36e705a6d2b0b614");
            when 32812688 => data <= (x"d369384bf57d3615", x"e8e55e5c42bb72f8", x"20107c6ee628a11c", x"a88b1fac27145d54", x"789bd4bd5a89cc80", x"e977901dd2e2d943", x"13d13b9eebe8dd9d", x"8dd65fcfc9e7430a");
            when 5331943 => data <= (x"f6c10712beac6a9d", x"e8915c93ad07a520", x"fd0ba7a8d1936a41", x"81a4c5a58e97f1fb", x"1914d0dd905a677c", x"a1a4e7d1f4f16f9c", x"1449ba0b56cbed11", x"ca45f31115af8f5d");
            when 3029484 => data <= (x"419ba2489deb217f", x"0cb547b0b48735ee", x"f0375d0698b2acb3", x"4848d370a3ed8272", x"e46793c97d56306b", x"9f79b1e8564342e0", x"2f6ff04b31267a64", x"07daea359d4ba116");
            when 33445194 => data <= (x"8831c1c339080fb1", x"7095648e83507a26", x"51e7992605bd096e", x"f0321bdc800b62ac", x"b4fbb5dbc4d36b85", x"10d2f2a859dfd834", x"ab87d1a92dc8e3b3", x"34e3dabae2430a27");
            when 16219972 => data <= (x"691951b7274994f4", x"ecfe384e66418c26", x"1987cd7d02f0c5e2", x"a50ac8e9b35cef22", x"c7acfdfd71cb1f5b", x"57824b66e6028149", x"f316b9872297c0dd", x"e31832b50c9101f7");
            when 11600945 => data <= (x"4e8a3deef96a0abc", x"e9172f14f2538eed", x"aa5b0fa6de25fa96", x"808ec67ec664763b", x"b1f1f575c11258ec", x"ff4a66eb2506fbdc", x"4127208616a3cb98", x"2491f32654721bc1");
            when 19291059 => data <= (x"cf525add2012a41c", x"f3d973e180ebeee0", x"f1e2b186a8b0389a", x"0f8235a15dc9644a", x"983ad67f33b87c50", x"50ef23a93d074b1d", x"64f98ef21b9df305", x"7ab4ac92afa42717");
            when 24829575 => data <= (x"709adaa150ca4cda", x"b4927b771c2c9227", x"9a9be22a496ac016", x"abaf706003fcb04a", x"9b2814b7642b544f", x"e5387a63ff4a17c9", x"d644a9c7110c0af3", x"28868273ef6ae261");
            when 20789458 => data <= (x"b5f8443e269f17c9", x"58f32bd1013a66da", x"c5cb252d7c532939", x"a3eae5659e39be90", x"f8c6bff60448c524", x"33eb6577d6380dcb", x"c3d0d979389af873", x"1f6676cd9b8a2b96");
            when 5511566 => data <= (x"5891b5fb90edd595", x"9508b8d145b18d7f", x"cf0aa7321b9b6dc5", x"ad839272d1f1ba91", x"eee237ef2790ed73", x"f48a7132fe6b2d17", x"d0a81730192cd453", x"351d4e369152654d");
            when 27663273 => data <= (x"4b1eb317d6d38bb4", x"6cbc103609c2a4ad", x"c0d3db936320c7f1", x"3662f8d6b917a332", x"8fe8e9cbc5ee1415", x"595731b393b18c65", x"74384db982206d46", x"b2b7db5c58d1446d");
            when 5691890 => data <= (x"3dd3d7b19fa29805", x"34e953b8c56d6611", x"8dbe9a0517f68c84", x"80e538cc3f657f6f", x"c8a461969476369b", x"24e8b1dab4a62479", x"0de84181370fc73d", x"1875adec4d98bf9a");
            when 8735834 => data <= (x"8ab25e5742d118f1", x"1667bd3798a1dfff", x"4b6cc28a046c9332", x"9f7f816a517fded9", x"a03f425e201f7952", x"b8d9bbfa809e4d9e", x"599aafd2d2d9371a", x"308c7707cc5ba263");
            when 14404947 => data <= (x"7e42997f85cc5084", x"dcc1afbeb866a629", x"d4a8e77b00f09d80", x"337df2e6900d9229", x"1e061b2d0caee0dc", x"32c11ceeb2c3e6fa", x"5d625f14a6912f3b", x"36fa22c9143fdea5");
            when 5290503 => data <= (x"ce08a05053512e6a", x"d5579c5e4c8f0834", x"5ebea69906f8bd7c", x"053b83c9dd78d03a", x"d17f11a5681bb127", x"e6b5a34c3f974f78", x"f8260b165dfb7ebb", x"235904ff8b9393dd");
            when 23629449 => data <= (x"aa37a4091253aece", x"d31df0bae62ae292", x"fa4350dd3d2fa703", x"86033bf0db857e7a", x"8834933812868585", x"cf541584c10a798b", x"0ab9df5b92c59b97", x"6ae13600188740a7");
            when 3145755 => data <= (x"17ecc8240c4eabb0", x"6ddcb9b256493673", x"db910ae50c8815ab", x"15d76ccda2e46011", x"5c4a66f7a6981447", x"8b85ed377aef0c0c", x"916b3118ed3e4661", x"5f125ff2ab1f7ec8");
            when 23540623 => data <= (x"d0b8205994a7b388", x"9840c58379d6a860", x"164e9beb126e19ca", x"3a5416b3347055a6", x"961e91a619797568", x"cef4094accb6be5f", x"2fd907c2332a1a87", x"814ea053386bd4a2");
            when 2709207 => data <= (x"32a4399fd60eb3b9", x"d262e5bb317b8431", x"2adb1e649693359e", x"9c841af1ea6811a4", x"c52ea7fa4183056c", x"fb4badef865a532d", x"c122a68adcf497d9", x"c4d6e41557f0f966");
            when 17249306 => data <= (x"435e2c1e87be4280", x"2f4d6b1f34993614", x"61790cb81be6d458", x"8248680bc7c0b24d", x"99fc802f37a473e5", x"e4eedba4b756f904", x"378c776d69b11932", x"5079ed267d9d2342");
            when 14779135 => data <= (x"e69d7272bc74b302", x"e420dcc56a2792c5", x"1a2f62c9f9566fa5", x"8f9223e87982c13e", x"88c2da210b1d0be2", x"8d531879a6e3a155", x"89cb1f0177b8f6d7", x"8d23a66876946fb1");
            when 30312386 => data <= (x"9d72a9a53531f111", x"e7d70b84ab519643", x"aabe1bd5b2ffd4ca", x"014cbfb522e8f3b5", x"91871c25d10a8e9d", x"7f5811478365ff75", x"3b64ea28fe723bf8", x"a02155196ac6cea7");
            when 24076406 => data <= (x"87c2a9677ee6dbcf", x"7fe95e69a648312e", x"df9aada646a2cba9", x"4b09f03ad918d3d2", x"f19ad60abe709560", x"5803fb54d39cb503", x"d51e532d5e52f6e0", x"090b7e608b25e229");
            when 25880298 => data <= (x"9a5242957941bcd1", x"49d4ac3177cc2439", x"16ca6a26d683806d", x"4c2143b7e2141018", x"3f41b668e3b6babf", x"e189abacf56e3cb5", x"7419440fadf15ccf", x"c187cc33d7a592dc");
            when 16037227 => data <= (x"1c4550b9cbb1614b", x"433a81e52b25f345", x"b4d660d687011cf5", x"8c0296fdd15235d2", x"acac85650da0ff63", x"2d5ccfa45e780309", x"8f6b096711918df5", x"b83b85c0ecb2c8b0");
            when 13004935 => data <= (x"6ebc10075cbffe4d", x"4b985398a6c2ea06", x"977fdfce797bac5a", x"991e0cd49d87e2b6", x"ab20f5105d81b792", x"acfbdad9f29fa149", x"af89f1a3ec854788", x"7da2078125623915");
            when 6346472 => data <= (x"3a04a1004ff90469", x"49de67b31f7167ce", x"e57c69d0f27d18c3", x"4b00eb855c016504", x"e83dce7f6a66db33", x"b29ea6aeb89b033d", x"9ec6abefcde69b4b", x"6b1eb36b4853bf34");
            when 23899121 => data <= (x"0d9af927c1308a29", x"26691cbe08b42110", x"bf48dedaa94c1cae", x"cd18fd70d678ef2b", x"085c5b07244d457b", x"f6ce64e9dc35e929", x"8d9c07a46dd96918", x"0e2720587f9d336b");
            when 9844168 => data <= (x"5496009561ba637f", x"2cb23c3f4a88b697", x"b40189e2f8970c81", x"5deb100b336623f1", x"f3f86b16986cbd4d", x"5a4e5e965ac4ca1e", x"a31a93bf4c15e588", x"6e976a3e835b5e57");
            when 12783603 => data <= (x"97427bce3510b973", x"2c4545366256c684", x"f11348a0d3413a24", x"f01eb8b480856cef", x"ad56e24003ef88af", x"568d1181924d1ad1", x"e637f1167d737a24", x"02b44b18bc526478");
            when 26747708 => data <= (x"2f20b814fe577a1d", x"730346cbaa65cd02", x"edd8f97a7646dad8", x"f1d9a5b1b20720e5", x"41aee5eefd91a7ef", x"f86ecd8413ed02bb", x"8a6cf78ab8214519", x"3b0583fd623452b3");
            when 21017904 => data <= (x"7456daa54ef5d293", x"162927a0773961b1", x"c65a4d095bcf87aa", x"cb34d105954cebf1", x"52afe0cd6149942b", x"d61f980a5073367c", x"4ab6bdf0f3639c2b", x"72f4edc9fe83e098");
            when 17700577 => data <= (x"4eb45241bb177c68", x"583e254310ede74e", x"c7f7ef63a68ec7d4", x"4a03054d74edae9e", x"9858e12ad9cb971d", x"b3c6a1e03da24b26", x"10007a23c2a2e4f7", x"020f2108b37928bf");
            when 6174913 => data <= (x"a746263cfecd341c", x"31c960b0d5b22d8a", x"772026d2221acd22", x"93b8ecdfbb4e0269", x"d05ffb5ed2c693f8", x"8f153c4010124a5e", x"716892a7dbb3c149", x"44f41ecc5f7e699f");
            when 2541596 => data <= (x"f4b7fd4ba438838b", x"a239425934a111d3", x"8736e7b4a5031b29", x"17dbfcc8214d2e09", x"47754938e9fe523a", x"0aaeee0b38a23cfa", x"e51961ef827d90a9", x"df9bdd0fed87ff13");
            when 25682067 => data <= (x"6637e5bca9b3298e", x"2af67a22aebf2e59", x"012431d269e57c8a", x"82c0e171cc051f62", x"6f08d24352e9a3c6", x"867c87d41b249e32", x"17e603c0fc191570", x"ac3873e1d3ebcb7a");
            when 8419058 => data <= (x"faf5515ad1e84ce3", x"9d4dc708fce22a45", x"4a1e26d15a1c6f4e", x"01a7a2a0638c2d3e", x"5ca6566f99213d93", x"4fc166113f40ff34", x"e31252941bb84254", x"4363de35d1960a3d");
            when 23486946 => data <= (x"8a7df9011071379e", x"0632a21ae7c63852", x"3815033f8b7ff0a9", x"a54776ca3fc430cc", x"15af8c476f67d326", x"52cae64b00ccb4fe", x"d3ef10ea84e098ec", x"ba7ce44bb3e4ba3a");
            when 24048403 => data <= (x"c0dd8d532399fdfb", x"82a38e96c7c75c61", x"40ffa807c94ca1cd", x"8d5aaaa97009685a", x"ebd23ad922ee1422", x"5395214fb7b06e4b", x"231b40c8274505a4", x"275cbadde8c40565");
            when 27030979 => data <= (x"dc278263a9847d98", x"3193bdb8d8d2f555", x"57361ed68a912d58", x"75202886e41bc01f", x"1cb80a94c26750f7", x"cbe8544cb2cba0b5", x"8ae2ce5baca86e73", x"52c79204870b9c34");
            when 11429891 => data <= (x"91970cde72833c28", x"c0423e7c69c91f5a", x"88772c45ffa51aa2", x"907568e833519e3c", x"7c7bb66d61b7c2cc", x"f93b3c2b47c3dcde", x"af57bdaaaf0205e8", x"f036650028ef3f90");
            when 10547944 => data <= (x"705da01467006fdc", x"b269c09641248257", x"2ff07f8d6e3387df", x"d5c6767c69249788", x"b055525c7339f534", x"74a493863d90f558", x"70359e48063d1e2c", x"daf70ea8ea5f3874");
            when 5473306 => data <= (x"e19d18d0fcde2f39", x"28f6a6690284d0fd", x"11d144c221496f5d", x"5b4609dc7c7031ad", x"b3f66c1bc4dab6ba", x"4b2b3878a3573c82", x"50cad2896ef11b96", x"f49075b990522043");
            when 19597822 => data <= (x"00eff2f983824450", x"37686743130450c1", x"6452f72b7f4f731d", x"5de0bdc8680474a4", x"0e76861f5578a7f5", x"0071041a760104ea", x"ed267d565acffec4", x"e775c069eff36bb1");
            when 18747332 => data <= (x"1e3430580318d019", x"f1b32c8e40650d46", x"0aae390a331ea88d", x"702def238543acbb", x"fd9d6358b998af45", x"444ec7e0eed67d7c", x"9318e2921b460b36", x"f2be4d898e9c3e51");
            when 7449224 => data <= (x"6ab326a5ddf24f6a", x"980c9696042252ca", x"986fcabf44054ec8", x"dcbe757fc2155af0", x"a0979efe8b872421", x"92bda76ce9a942f6", x"c2ad50226be2932c", x"33a5475994cfc867");
            when 25717126 => data <= (x"e4f0d9ace393213a", x"5dad73f32de57aa8", x"5c3af6558c8cbab3", x"90ab54c30a074d95", x"91e51c0bbe77c137", x"8e1e830b95cd3cb9", x"64fa29660c58fdba", x"ee4fc4909ac434ae");
            when 15762388 => data <= (x"37f9e86425429a7e", x"6e2542c070c1eaae", x"4ca2ca4a52e28552", x"5e7621cff6fc8e58", x"74f69853c58b73ed", x"ea0ff03dcfd8a512", x"c456698bd2fb8097", x"03c6c1c2cf4c009c");
            when 28006262 => data <= (x"1fe3ed9fb63d18c3", x"1f4b855521fb41da", x"127f1192de649693", x"0e0a26a5f018f3ae", x"8c3b9fdf87f3cca9", x"3f130d69b1116433", x"83a2447bbbbecc2f", x"01f264d40c453412");
            when 27966502 => data <= (x"71856502daab2b69", x"468bbb9ad8299431", x"56f98c19feb6afed", x"af26681d19b3aac3", x"2e319f342030628a", x"520458566bdd401e", x"3f9bb2cd1e6fc063", x"7e9bbcb433dde2fc");
            when 33873449 => data <= (x"3e92a5542551f990", x"e5840ac9418c41a6", x"5dd20a82937557e4", x"d833af6c60bfe95e", x"4d96cd6174228e14", x"fe232c1bb344c65b", x"6b48afe48fb0b289", x"b7abeed483acc317");
            when 31758555 => data <= (x"e04f00921f858c05", x"afa299fd13193fe7", x"3a0638a8d29d1161", x"2f2986deae1e57f1", x"876574434b7995cf", x"2ce3bf5f5d5ae103", x"e52a1c6297fb5d4d", x"ef456a7bdf51cad1");
            when 32930894 => data <= (x"894418afdb9f7cd1", x"8d54c6f3b0be49de", x"614b5ee778348db7", x"68b8bf71ea25dbba", x"0fef653a743fe452", x"fa517c87d2645315", x"63edd80817b024ea", x"a760dd5675890a6c");
            when 29222090 => data <= (x"f7e07c7cfd24a8c3", x"eaeedec95e7cfd5e", x"93e959b3cf4957c4", x"0a5ea7a87440c753", x"d49c27c8cee50f83", x"c8ea6f0160c0e943", x"4455649256050ea7", x"5f4826bc3c397bd2");
            when 27916012 => data <= (x"a0c0087473e7e077", x"cf2dc105ba3d8d60", x"7f0a62f482398cdb", x"8fb44fa136f700e1", x"07d9cf5163b2f41c", x"22320f0c46d3f95c", x"c576c296c0d0b36f", x"72028af3bac8bebf");
            when 5162390 => data <= (x"761f1aad9cee962c", x"778808a53369411a", x"b29c47d9869100f3", x"1d5fc0b2c7d77967", x"0274fac97dfa8426", x"b792eadb36c0deed", x"31e237ed1f954451", x"9f0f7303fed8d45d");
            when 14362837 => data <= (x"948ec23ce788851f", x"15861a12bc03322d", x"f28418c6a33d279c", x"67a9fbd76a8c9598", x"2c2e8efbf6e354b2", x"d9bd08dbf33f8e9a", x"a02bdd18bd382f12", x"9a069f55f5b55cc3");
            when 32839893 => data <= (x"09427ca6ee8f600d", x"1443ea1b84808367", x"7870067d5d61fcd3", x"16843847dc420e8e", x"999dbb0ebec075c4", x"92e46b8208330ee4", x"b68dbf6aef975703", x"b95dd9ef63eaf85b");
            when 29639079 => data <= (x"f4d844fed2378ecb", x"57b184b1b578bc03", x"73274cffc3f69467", x"0343cc19aa8a8605", x"39c9551c5f1248f7", x"53f19672df834eb8", x"193a198d41b2dfbe", x"636a6ce9648efc27");
            when 28194766 => data <= (x"3491a84575536993", x"e68b01689af8f62e", x"71a86b0492fa9688", x"c3f4c88601f9685b", x"a148671b3f090075", x"61e5b2010332fad6", x"5396fc9e5cdd6eb0", x"b0dddb7c45d274cf");
            when 21832874 => data <= (x"fb3412117ae05a6e", x"9bdeb3059a6e04a5", x"4f927ec36c4bd948", x"cd8fd4866ac481c7", x"6ce614aa0906925a", x"e29dd3cdfc08a227", x"b9bbf99a4adf2764", x"a04ef47a2406c0b7");
            when 27361645 => data <= (x"e138b05db8e9760c", x"b84895f32a0ff257", x"9ad4b05761e5ea7e", x"e3895834c4ed7b12", x"e666e1c60d051513", x"b522caff75352d16", x"696d4e0cf76cca4b", x"1c49dbf7c36284d6");
            when 23740324 => data <= (x"659b91df22731378", x"102ab80da2566178", x"cfe9beebd2023d71", x"540768186422db7e", x"ebf665018344809c", x"c55c9099955ddb94", x"c4eb818bb6bebc93", x"cd66c7dec7b8dc22");
            when 29041251 => data <= (x"fece076b12fadb3e", x"0241802f63818913", x"f3d268ca979cfd78", x"cc08cec9ec0b4020", x"b5f30d36f8496b32", x"225f89903a2f1264", x"a12d4e36fe60e71b", x"c60abcfb0cc17b46");
            when 23990923 => data <= (x"addcb9e6672c1b89", x"522e536fc7336422", x"8cc0922720bc1848", x"09b15610a9fc01c1", x"1880485444547996", x"318eeffdb5b37151", x"fa650a6df6cb2131", x"2d2b624b41106a36");
            when 27437042 => data <= (x"7ad377675e97f889", x"00f2a954cd7139b5", x"23b94fe2cc640c60", x"a39c20e8a04fc97f", x"1464109689311a2e", x"ba1300df3f85e45a", x"9a9d938f7e63b7e6", x"9b53a656047891c2");
            when 4526386 => data <= (x"1d1e1bbb3a03d134", x"21f72c73807028f7", x"93b320c9f10b8a64", x"f649cf71bde6ad7c", x"698b02796958b318", x"3ff8e38df35c49b1", x"8134ebde405c178b", x"f61de777e332686a");
            when 27559693 => data <= (x"f90d0acf85abe517", x"4584585473173b0e", x"2f5d9b41e42b9b71", x"cd70b6c2b6e6c00c", x"c149362f349be3d5", x"053d5b2bfb9f931a", x"2a79bf1ffc4a62d5", x"7a1a201ef72e5c19");
            when 29884365 => data <= (x"e6db154671654aac", x"923ebf9ecb9a75c2", x"b9c7a07505697fa3", x"0fa9c26928d945d4", x"a8d459549a934ccc", x"845e86f1fb2b330c", x"0b395f9ed137e1c5", x"38a0293da46d5ce9");
            when 931354 => data <= (x"ffc015830c92f791", x"718bea7a12e42ff1", x"7251f5291a2f0f19", x"a38515cf50745931", x"511f1ed5e604f24f", x"1c2a43162004a6de", x"9fcafafb43a519a0", x"53b8e9ea419fe0f3");
            when 3860158 => data <= (x"1dfc75964d533c08", x"6cf21ad714885e0e", x"2d4bd4997ee9dc62", x"c0c1b28e584db0ce", x"2cda6352d39324c6", x"ca27fa1cf5f8e3f9", x"3b9854749516dc78", x"8be6d22276bc2716");
            when 28886817 => data <= (x"f3746cdeaf6183f5", x"af7d97e9d478d3ee", x"2a5f25a341f62c94", x"969897fd97ee78f0", x"8d706625ea61b351", x"621fb6f89f020cd8", x"fa114ffd1f356cd3", x"7a1795b40b11aea1");
            when 621682 => data <= (x"a9d8b9535e3c2bf7", x"475075366be8f5c2", x"95fea4260d0ad1b8", x"aac75020facf000a", x"752d2a8fc0983f1f", x"89933c1ddc5ba300", x"9965daa35ef8f0c3", x"dd5d887fe6e409cb");
            when 20648900 => data <= (x"6a3796e5e43f3d80", x"7d2c89e91cc0235e", x"9bfeaec7fdfd5905", x"f4574e4edc28d389", x"375b8d63cfa50a87", x"18916b39c1f09c32", x"27f1bb4ba9164c74", x"0473f2a3e94b1dc0");
            when 17768112 => data <= (x"a6d0f7c2d28200b3", x"e957daf65542e2b3", x"3c2137fe78341cf8", x"e4011a3c42a17ea8", x"039b28b9d00dd16f", x"65937db43b7659d3", x"e9adcf2f58cf66b2", x"e8712726c3049b23");
            when 7456421 => data <= (x"7d3ce68b1e39eea3", x"5f8abf75f83a370f", x"2f47b4ec2c15d459", x"663a0e070a934457", x"48879389deb2ad14", x"787e8c6785408d0e", x"89b35a274f2927e5", x"fdb0497b54155520");
            when 3341540 => data <= (x"c63a09cb89f780dd", x"ecec74a45cb4925c", x"6d88d16319e1e548", x"804ba1863d065500", x"229ab4399efa561b", x"0f004dfe587cea50", x"f346c09b1c73d606", x"26132ba0c8a15641");
            when 623598 => data <= (x"bb3962537236d381", x"dd9ea69eb13b2a30", x"61e964b713907839", x"2758c2e09ad0da0e", x"3660c08191d9389e", x"8ab221ea2835ead5", x"d0c250209fa43699", x"1d9deee9cff33488");
            when 7448355 => data <= (x"a81324295bfdcebe", x"226664d6a305c59a", x"fd4858d3f4109056", x"65e9691ccd9fe5c8", x"02cc7bd45b17496f", x"28d4638f5feb8340", x"6ecee67fe56c43bf", x"f0911997d6642e98");
            when 8420705 => data <= (x"90af9e50a57c9979", x"22685cd83282f33d", x"f5431f05ff68eb72", x"18056aaaa35ae972", x"18e7aa82ed48e2b2", x"c062243a21da7d05", x"43f40f1724a3f0e9", x"6010c553117c855e");
            when 10534573 => data <= (x"69af0bd255227e3b", x"d517ef5b40e6615e", x"6bfc0cb01945c31c", x"ff9943ff105a8da5", x"fafe2c81e09a7465", x"7c9236c1d046b3f7", x"af39bf334c7cc96a", x"fd49d0e7913d37bb");
            when 31166036 => data <= (x"32c2ddc4ce70072d", x"ead16f581a4a263e", x"d8f99c5afdb45583", x"e2f40365e1d0bb44", x"4094b791218b68f5", x"a3bc589543d22c89", x"b4edde8bd3fd2504", x"2dae67e3495346cb");
            when 4386405 => data <= (x"0fb87075aff08b68", x"1d77f54cd543b37d", x"4af2abdc6d8ceee8", x"0af325bcfc15b897", x"cc9fe5ef0cbeb68b", x"2c8a7b44ec42ba8a", x"8ba59785d5c292bd", x"60483a53b2c1c566");
            when 16048829 => data <= (x"35b0426203559dfd", x"6529249a2343c677", x"604cb03c94cadb7a", x"94c8468543a4e7df", x"58dd4c42568d108f", x"2fa4b48b79cd1130", x"51e0a087094f25e4", x"8cc2fff467abcfe0");
            when 2936997 => data <= (x"c9ef2c3cb5d38c49", x"ed6f0319ee3d1bba", x"85884b49815c6c8a", x"11098d357537a9a7", x"62b8e11e39050ab5", x"9062235cb6993cac", x"ba1031f1d32fe3a1", x"8c51faaef8a8fcfe");
            when 8824365 => data <= (x"9ef1f00177cfebed", x"d3989ca9b8928f92", x"d758add55bce4de7", x"332567d2940cd82f", x"f4d67c9c9750bd5e", x"e25a438407aac8dd", x"1bfcacdafff546ff", x"623887556b3988f0");
            when 10765492 => data <= (x"bcd05e71a74d4f7e", x"0cc342dc010d1dc4", x"a5b1be599e2ad79b", x"dadfc7e6b60a0390", x"8beab7a005418ced", x"bf0443f2821f5c7e", x"cfd91f718409c8ce", x"827ebbce6e567d7e");
            when 14271299 => data <= (x"3aee94fcf78fe33a", x"4cc16ef6e2840fce", x"54c50f989ae1e2df", x"548769618ca60546", x"27b0e4c1880c5aef", x"34df740800de524e", x"f8a797ac44ee4c60", x"1d113aae694c824e");
            when 22454877 => data <= (x"c58453a82e60ced9", x"49432a05b8b36320", x"43163f1c8fac9397", x"469f7d45fe969b16", x"52e4cc0d14feb7a8", x"64e8042a23796289", x"26a19e1a821f82f1", x"fb20415d58b3b711");
            when 14655813 => data <= (x"cdcf02126c8a5a1f", x"1827b7d7f51a6471", x"263157cdb62ac581", x"708433037c2f59fd", x"e079ad38abc876ef", x"085d2a2d941df1ef", x"bb42a413352abde2", x"c2b9377253b52793");
            when 9905827 => data <= (x"f643c65d715801d6", x"67fe3b63088b79c6", x"b20491c5989a9d64", x"e1db52c9b4b957bb", x"e862b26fbca770a4", x"ccb04c5940eb4de1", x"5e17c2eadef224e6", x"2e3c6b74165bc426");
            when 26037631 => data <= (x"b177a5dbbf47ebc5", x"9340375aefc6695e", x"a97c4df565ba518f", x"5cfcdbb5c40c83ee", x"031142836067dee9", x"928293da7cadfcd2", x"63b49ed40e32cd23", x"bf57128631c2c755");
            when 28338227 => data <= (x"b155c778ae36f887", x"bb846435c736fa22", x"1a61c591eb23bb96", x"1ec9433e39da0c39", x"0f37ce2b8e4bec7e", x"c9546e15b30e3e14", x"de421025cead1f46", x"1421c8567c9d5fca");
            when 3272460 => data <= (x"46acb50753c195f3", x"13934db80ba053f6", x"2fb4cde3a56a0021", x"20bd096ca1ac7a2e", x"08d50bc308c6de8f", x"9afdffc9ceb02d12", x"ce98c6864b0fd2a5", x"48994695bb7b7ce8");
            when 33505635 => data <= (x"c5a476297d62c668", x"50734a9f54a3484d", x"ba9c97f982b965d9", x"37d782d198186d3c", x"13dfab89c1c406fd", x"08f0fa7735cc105c", x"9454b458ffe463e8", x"e89e62f074bedb9d");
            when 7342416 => data <= (x"11b04c9af7eeab1c", x"e04bf44778910565", x"1a4d9cde0e275e54", x"692ba91a9ec2139c", x"75586b56d41ef5b0", x"85007e56c8001895", x"d04a0d3d7855af13", x"333f703a4585c936");
            when 5359157 => data <= (x"d5769b92ea187510", x"5be6c22eee8c025c", x"1ef341e58a785a6d", x"8ec0e5c0004b46a7", x"d71f9c4878aa1a78", x"7c6c94ba4968a789", x"144b775e4ee19ea6", x"9cd4ae5707969d30");
            when 9664728 => data <= (x"863dc2d8c4ae30a2", x"9878c0d6ac1758d9", x"c4e8570742f97887", x"811d6e594ceac513", x"1f405df56f38512d", x"78b7b2f97bd78771", x"1692f7a7feff0ec4", x"32b4a7266419e442");
            when 2890216 => data <= (x"c9dac40a8e6f4b16", x"275d11bc064b04e6", x"fc7d7eabd525261b", x"2f5867b0e6895679", x"e3b3be39e32555b9", x"3b503eb042b02692", x"00668807f07772a0", x"15f8a23a4c0b0bf2");
            when 22128729 => data <= (x"203b43ec3acb86dc", x"1af47579fd8656e4", x"73522a7a9c397772", x"c2ff579974c620cf", x"a49a075d1a5d0d83", x"0eb9c5c1686825f6", x"4639950c71e03d2f", x"756b73593345d897");
            when 27773924 => data <= (x"5b0797ba6d29cc97", x"ce6fd5ce09283db3", x"d6c1deeaf994a6eb", x"74264ba3ff26f850", x"e6950ba81c083d08", x"632b956db2a33520", x"2ae38bbea91fe7a8", x"eec4dbe1e87692e6");
            when 14529329 => data <= (x"dfda3cffca0fe958", x"c560a0cc90036363", x"a24b8effe610e208", x"8bc6fcd043906adc", x"7a7ccc1e521fea0c", x"4355587ea89b6163", x"db1791235222722c", x"0f49a9ea8d9cc443");
            when 24692107 => data <= (x"3d3a6f9227d1a0c4", x"40dd3c7eac14b58e", x"f9682bd80b7b76b1", x"952f1e23b4fa46e3", x"f83b5a07cb95108f", x"9ff0a51f94fb9bb8", x"c93c21b1adce268d", x"0d724f2b87fd8779");
            when 15301824 => data <= (x"604f38099eefdf8d", x"68685814b7e61632", x"9e97b8d0ed834cc4", x"b414d61669cc4339", x"9fb9e7435f0ad9e0", x"48e14b0c1ddd1753", x"027fe27540c96be9", x"0aba0bb21be8e32f");
            when 16790488 => data <= (x"39bf78af43738f91", x"58fb3b44c4a43d29", x"1dac0d3954ebd37b", x"f4316a343dada65a", x"93df7f026953f36e", x"cdf83fbd3bc4bc74", x"d053c019a1395acd", x"5fc6a3c0b6444b00");
            when 33587264 => data <= (x"1bf8d9554b1b4d21", x"d94871d450d07757", x"7a8414c9b5ffa5ec", x"83a3b480284dbd7f", x"eab68b9d49143e82", x"789efe40492ba9dd", x"329c94a108a9ece5", x"6a80f4a84bd0082b");
            when 7354874 => data <= (x"cfd04c421949d8ee", x"e7a2b3fdf67250c5", x"1495d416ae567301", x"9c5e7fe674aeb834", x"d0531ac10a02bd37", x"a759d4c1365ebf43", x"598b96cbf363c7df", x"91516df8820d08c5");
            when 28797059 => data <= (x"c9027e640a310b18", x"0489c470dd10da89", x"298acbe7e3e639d7", x"100f4f28b0c74401", x"170536cac9b299d4", x"5fc2588426061118", x"24cd4498ddf5bc48", x"a54d6f28c394db1c");
            when 6171400 => data <= (x"2c7adb50cfa1ec8b", x"1b85f214c6aad775", x"017de81892a8017b", x"cbaba078f56a8690", x"43244503ce60e28d", x"8656b4d894d565b0", x"95dd5f997edbae8e", x"2ffaabd015cba205");
            when 12270361 => data <= (x"652fa769d3a911b5", x"a1f9643345472fa2", x"32b04904361b9502", x"945be4daf209047b", x"9afaacf8cf5ad876", x"6ec384f6aca545b8", x"815eebb9305ea7a2", x"9808c8d7143bda5c");
            when 30294212 => data <= (x"c06433b073a8384c", x"b633c14a64eaed54", x"9c400471f6911282", x"4e3df051f23eca32", x"5091012a4a4e40e8", x"a84e4ef14ebfec1e", x"9b5e709c5ce5b3f8", x"b62f94e82e4706eb");
            when 6421603 => data <= (x"0ec72f686491ae42", x"ff9d743894918293", x"be6c31ee58e64fc3", x"91384f84b801368e", x"3086130b295e64d7", x"687ffa3e23b2c9fc", x"2edb0a245c5ed324", x"42ad742d978fca0f");
            when 3401070 => data <= (x"259e2d1039236263", x"0056a906d0da0bed", x"c867086e41403915", x"1730b85af0bf293c", x"c1bac722d58f437a", x"6d872ff6e8994e41", x"48e5f7a349528162", x"0e03dd35e443517f");
            when 2076107 => data <= (x"0ecc8c8d34856a98", x"bf64394c51b17457", x"dca3d8f28aeab8c2", x"52e16e5da266ec4e", x"871cbd742683da7d", x"2c7f868523a3a827", x"e1818437f7dd99df", x"aeb2895adc94d849");
            when 14327498 => data <= (x"41bb949a1d935f4c", x"e0b003aa5a4445b1", x"76c8b0dc549bb657", x"a96081347235c9d3", x"ec02345082030ed2", x"63640d432dde01d6", x"ccacf3df652af93c", x"27250f4921f312b1");
            when 17738755 => data <= (x"eda7883000f2f3a5", x"18d482ab40acae69", x"9e0f367830c66b51", x"5467aa2c5701a291", x"530c38b5b82b3a4b", x"a500c9688de1a930", x"0ea8425fcdcac039", x"696cb6078c50c6a9");
            when 2115121 => data <= (x"5a4cb2f0402c882e", x"396ee176cde159b8", x"c3631b31733bcc8a", x"48e87bbff22a14d9", x"31035161b36b02d0", x"b4589b413e4fd8f6", x"4abecc94856b07ec", x"ebcf14b7a24b8ec5");
            when 24617151 => data <= (x"3e1bffc58e0040e4", x"84a46ce9a43b3ced", x"461be917297eb019", x"8017d7870cfc3331", x"ea381990b500fedb", x"5f8af6001f266e78", x"0e988a337f2a6454", x"191efa1e6104e8cb");
            when 21019203 => data <= (x"5411463052628082", x"34f09e9175530603", x"fa3e759dc0e90148", x"c49cd34f63dfed35", x"11011f6f739d78b6", x"221924367c303f0e", x"a13b624baa5fcf0a", x"a832456197800bf4");
            when 15401353 => data <= (x"410f92da28630a66", x"b583e1246c030311", x"9c0f8849ec4b8c36", x"dc2fb5c9a3ab9a61", x"3b46194bb41c0b46", x"7f68ff1734add07b", x"3e2a0f643cc5dd1b", x"350e66885b4b0a8c");
            when 10098640 => data <= (x"bb43946efd900a7c", x"4cca9d0cc3b62380", x"e7f3bdb17db5fd46", x"a4db1fe103810293", x"c71094422f4e3cf1", x"643b7828a0a773ee", x"61aa532d8c872c58", x"65d740ca031cbe13");
            when 20350267 => data <= (x"4079bd7263dc33dd", x"8a5a74d45fca33f7", x"fc18f8df0c28aee6", x"573a722147f09f71", x"17175cde910f8078", x"bbe80f296a6ba255", x"410ee8452add2a55", x"7b6242ca930968cf");
            when 4920024 => data <= (x"98e4b6ea9f28042c", x"25b55c320c528d6f", x"e580ae88884ba6a2", x"a92cde94de59314d", x"446aa8fb9419a31d", x"4b5fc20b95416027", x"4e89958e2885b0c5", x"ab8ca165a1e62c9d");
            when 13480773 => data <= (x"b1a42851b8b4c66a", x"3caa32508db76331", x"1c1b79c667624b56", x"8c1a92c2a03ccb8d", x"1a459b010427be3c", x"66d2f148fdc3d33d", x"f77fb67b1ab861cb", x"f56746c65532b96b");
            when 13260551 => data <= (x"0282075af7ae1d5b", x"2a353dd4e4f63799", x"fa0925656db54c25", x"3bcde29a61cfef98", x"cd19e423922f5823", x"abd572d4d2d61612", x"e4a10981394c7896", x"3fba0cf695b580bd");
            when 7864944 => data <= (x"ffdacdffe54bcd08", x"e8c7434b6f09dd11", x"4778c041644fecf7", x"7039ec9f219330ab", x"fe3603ba5cfa511a", x"d34baa2040d66313", x"f2c4ec7085d5c68f", x"678ef47d05368a6a");
            when 12813963 => data <= (x"9c2c0ba477dd1746", x"e080490a2b15717b", x"8f21f22faf44036c", x"480a0b7e58ef9b5f", x"3b7a59896fe139df", x"df11ef35cd517df7", x"24c5325dd3e66e0d", x"903781e16a85c2f3");
            when 11878463 => data <= (x"ca49c4242b719849", x"4fff4265760258be", x"7b780b200e5dcc90", x"7c960f9baf789edd", x"feff01e97cf8bbc9", x"21d5963f5d5d101b", x"0da5d71f8c0b6f6c", x"07ebc51ec29053e7");
            when 28888602 => data <= (x"c58ac484791dff91", x"2d37c0a1628b979a", x"0f5bd88f391d9ae5", x"bebee08e31aaf6cd", x"aaceddc572c8b833", x"dc48c5d6ed74f22d", x"4e66623734a55015", x"5ad525b2002155e1");
            when 20967116 => data <= (x"f7cbe9023b6f2922", x"e09e9d7c6c08a503", x"061caebd3f58c18c", x"871de70508eefe0d", x"43f465f95f21b67d", x"97fd5be7bbb690c5", x"c1f10b1e27f48516", x"ec650905fad0f800");
            when 26693122 => data <= (x"1fd107646d31d0c8", x"437737de4272b4cf", x"2dc07c5cb87debbe", x"dfec29f5edd98b78", x"99cf4ab6937be499", x"a60194ce42503048", x"6f70a5d798b50213", x"d520338a11453d67");
            when 16481528 => data <= (x"52a63427141e5fc7", x"01016819b4cc7462", x"bb85f4afafefb0db", x"a326422f9cd1118f", x"b1528665dc7a9efc", x"4300a63cb5bd567e", x"f319c664b5794776", x"9d235601cbea8b68");
            when 28780363 => data <= (x"365bfea8c06697a4", x"4da4c8e1218fad40", x"c18845529e1523ad", x"53403a44b9f66879", x"8b2757335031a954", x"4ab5c17a96556a97", x"01134c9651e46a56", x"b98435784b385855");
            when 9857851 => data <= (x"8b757b22fc234e57", x"62fe1ba290f7acdf", x"08c7286b61a050c8", x"76173a72837e308a", x"d620d705e39eab10", x"9ddecae5a20b727e", x"b023eaf82922d06d", x"aed269f5003290db");
            when 14143708 => data <= (x"b77d4838a05dd9c3", x"efe0a04c63b34cb2", x"ec8f942936a3e136", x"c5128f3f7af085a3", x"33aee42175ff6a07", x"62594f3fd9d9df65", x"a9b2caecd945671d", x"43c4af398762b226");
            when 11696176 => data <= (x"36b4e73e86880859", x"ba768e038d850619", x"4f75710f9a9e6f1f", x"78ebd6d0295d4ade", x"b49897cee3fde040", x"358e402b8715129c", x"dd35c3b081fa5de9", x"0b10c22d9df7130d");
            when 27824468 => data <= (x"ca0069361108343b", x"1be8b2e9cfa1aa44", x"f9cdd504e2e2898b", x"897c8a7f1df265ea", x"785510ae260c5f31", x"9cd105fcd5fd95e9", x"0cd6ff019f66dac2", x"e13140de12c44542");
            when 33085148 => data <= (x"a1151dff3dfea81c", x"094adfa6d72c280f", x"e0b1b12eede4f752", x"80e160e0bab8d780", x"e4020caea69734dd", x"c14779bca46afcce", x"900e31d81c908ff5", x"397a9371ca946d7e");
            when 21073995 => data <= (x"6b228f29073ff014", x"45668b53a941ddf1", x"6a0f081fe677fb80", x"369877810df59f05", x"877dfe7f7a56bf0a", x"aee8fbc98a8dfb85", x"1b1416bd33367f0e", x"917471306ad1b262");
            when 1555412 => data <= (x"14827234083167cf", x"739860570760d8af", x"0f14f2346d1e5af5", x"d0f92f5008c1ecc6", x"455d18e49357f5df", x"9c4b93e1e75525de", x"d34b954fc81b71d8", x"61f632cb2b426ac6");
            when 12678660 => data <= (x"70d1646bdbddde54", x"9be391225117cdad", x"9c6ba3c0af61f9ab", x"7ea81ce0608c5383", x"31a1c4c0db34b713", x"9ccac09d63fd6885", x"6b07d3ad2500c341", x"33937da47d36951b");
            when 16458147 => data <= (x"69a9c07d127e4f28", x"31e9986bacebde85", x"9121c49724508c01", x"64f806b974e03c4f", x"9fd3fb67f6217542", x"a6a25fbc9ea27c16", x"a10a1d64e6af5c31", x"204d76e776d85128");
            when 8972796 => data <= (x"f89154a37048660e", x"d81616a0dec56bb3", x"bef2994c69ab229d", x"37054f7c8bfe5527", x"687f177146bfc1d4", x"4b022f9a6a7c646c", x"8366fb3817495e3b", x"d0d77bc92088379b");
            when 12843681 => data <= (x"4b79b76ff132c381", x"79c636ef14eb8b05", x"2f23a4f30f4f368e", x"eeeca977711ce721", x"988111b92fa3c980", x"f89e588989943802", x"69a08778cebcbb53", x"6d3ed3c5ee3dc218");
            when 7439734 => data <= (x"0dd26d2747d6bf12", x"d255fb4158a6f1d0", x"19adf8cee227a3b4", x"b05a96dde13c10f7", x"2c8a56e4910e92d6", x"739c9302c98fdd24", x"f7d1428483e0e800", x"2b0f7b0942395b9f");
            when 22009797 => data <= (x"4633dfc24b060230", x"990dc53cb978e4dd", x"c67d26e97b622c05", x"e7e2f85d94296167", x"f939b05a50608ca3", x"075f64d2b621c6d1", x"35a80a5d95b2d153", x"4336d9dee6d75845");
            when 28200155 => data <= (x"8a997e893de1fe87", x"5d2e27cf8316920d", x"a05db4bd0d63c120", x"5cfe628f686e692c", x"cfc824f12ff17e48", x"39ac0ab2bbd86ceb", x"5307184f1454a5cc", x"8e40b10b2038a0d0");
            when 21630270 => data <= (x"f9ffae31e1496044", x"9f96e1af1ea7ed53", x"bc3cf09e4932923f", x"d941c46c2213a916", x"dd5d0d80427e1eda", x"81bf578504d03b96", x"5e75b7420b4ce3bc", x"6f074e507f158279");
            when 13387162 => data <= (x"468e4d04f92ca873", x"081cb2684309659b", x"b906564bfe207222", x"1ca9afa5f8a32b6c", x"1baf173753482276", x"97f8127f9d223f12", x"5e386b4db71d0a99", x"a5a25d8a7fc542bb");
            when 19058401 => data <= (x"1f871100ce93d18f", x"c41cd39632979030", x"1562919b893d4314", x"1481a8002ca2b51a", x"67d02b1b6ef2f45e", x"1bbe1ff8d0dfb2a6", x"6246bdba0bfba321", x"1b8840af7291968f");
            when 16367745 => data <= (x"c74cc53ecac63e20", x"a1d91b7009a12bc3", x"7b7ae63ba09493c9", x"4aa6c8db94836dfd", x"123d86cd8db0c1ef", x"921b2fa9b0f0800a", x"a557f5bb4d9f2d00", x"6eaeccaca67e7f66");
            when 5084368 => data <= (x"67da1f5c9ad80e5f", x"656592a223c32538", x"ab2c639fba27b9eb", x"1e52317f06c9453b", x"8e2827a047d69d5a", x"859fc75f0c3e0ade", x"8520eba84276c2b7", x"227dbda4831f1bb4");
            when 8564377 => data <= (x"87588b5cce2f6d6b", x"75cc07c1f0cf7aac", x"22eb8fed34e14aa2", x"6a3957e7d997d7bb", x"721c1f93fc86c7b7", x"bd7da6eb137270fa", x"d5cd229610df1160", x"26a86b1f03aa1648");
            when 25239913 => data <= (x"8a015618b3cc8894", x"3dc55c525021c3bd", x"eefd411c6f2bc77e", x"ed646390cbbc1d36", x"cf448cf0c24daa06", x"d1e807a722c35f61", x"518797c436161c49", x"429850951e8b37a2");
            when 33983141 => data <= (x"6e306760b3586774", x"6ac298b908e68009", x"1f5267f90c896406", x"1d4099544d9535fa", x"2cef0349f82e10e8", x"9ca1ab7e05891f30", x"2cf6a5497e4769c4", x"4a1445936649f910");
            when 4434088 => data <= (x"63f80b262402410d", x"3b32cc0d25436341", x"c3fa4a0e7802bd0b", x"c36e3f6ddae11d63", x"0a529abe57b7197b", x"80c9050bd7209771", x"d017f8ff5c82c282", x"627bfb201d7f051e");
            when 24715138 => data <= (x"25c23dd011fb81a5", x"cabf346bb6428547", x"2a9a2d38e4abb3d9", x"5f1d6c476f0e1f81", x"3c73ecbcb928a132", x"09e804804137afb0", x"74b597fe1781fd79", x"a65a12b911d998d2");
            when 31443051 => data <= (x"afe08a5908d87ef2", x"2306d5779837bbb9", x"a1b658fa81871d68", x"04c079001c9b9293", x"4bd37b5b92f4c518", x"4642ab0d18b8b0f1", x"be1f6a32bfd77482", x"8c0cfeb388450cf5");
            when 32065619 => data <= (x"b8d9a88f02e340c4", x"6c5cc272694431f5", x"d74767e5644e5196", x"ce8108729036788b", x"ffcf8edec3c3eaab", x"fac046b665661cb5", x"44950e30f0bad18f", x"5abc8aa975f8939c");
            when 30928606 => data <= (x"c03eb1a149d80268", x"f4a208175baaedd8", x"dfc43f59217d3b88", x"dbdf68d3abae4d1c", x"cb95fdcf31fc639a", x"6b13d660116155af", x"1511524f1fc04a54", x"0c2bbe22b035d768");
            when 2164222 => data <= (x"035f9c24b37c3d7e", x"9f09618b2dada083", x"59514391ce48fe76", x"e8d63b3da5981061", x"2d52148c80151b75", x"476d8a27d817476d", x"ebbdd90fa5b3a931", x"b51e9c37e100a7ba");
            when 24836775 => data <= (x"8afff16ce0b0e526", x"944acb194124b9e1", x"57770c99a8f5feea", x"3d7adbfaaa7dc159", x"cfb076c9ae23a22a", x"4a9754c8b72150ce", x"aa16231f57df09ee", x"a8958fd8d663b3d7");
            when 31469790 => data <= (x"c35af6fa3e137524", x"1f9c0b70c9281219", x"fb501a182e009da9", x"657b0452044c69fa", x"af3022239f59284a", x"c0ed1a35559b78d0", x"fb411eee3e6ed826", x"ef87bb7abfc4671a");
            when 31818104 => data <= (x"038c5cf82f8c72ee", x"2461d75877c70e7b", x"9b96a75fb76a5f09", x"e5fce15349f6728c", x"f88e2bb24b0882bb", x"574a3a14ffc61ac8", x"dec54b639577185c", x"cc9e1489bab849b5");
            when 14632306 => data <= (x"16aea94fd22e5d8a", x"7e066ac7ba2d7395", x"c734e35f23eaa199", x"6ec53d10b160f34e", x"b2eb666711ab58cb", x"4f0f21693ba81385", x"1507345d05842851", x"6c7d9be91c98404e");
            when 15974701 => data <= (x"d0adc99718a1449f", x"6236a2f4704b5a9d", x"450810faa381993b", x"cabfacd2ce2ed242", x"4be1dfad19bf213a", x"09d6db3f7b02a782", x"605bd5c4d11c3e53", x"2ee6e7778333acac");
            when 22733305 => data <= (x"e9ba527a0654dd42", x"abc4f5aca9178407", x"dd82ddf10d36d91a", x"6d91bf44884a78a8", x"c447d0550a0ab13a", x"ef8e8c00ede63670", x"16a16ca8f7c0bcd2", x"73be509de46b19dc");
            when 24798296 => data <= (x"2b08e201bf10ce99", x"39db5870df5de702", x"2d10b2d974e6de39", x"8671af42dccc9f84", x"3a72785e2f7395fe", x"604b6500c8d46535", x"0e0cbbe649123720", x"07b5b6d1c7e32c53");
            when 30906410 => data <= (x"a030c666ec06f784", x"387cea5e167d2789", x"c47b01391b532dd9", x"4f52350f2c79ab26", x"4c38bc55c6e8880c", x"821f77d2b313dcc5", x"d12152a64f7fd225", x"49ffb059f88ea411");
            when 16503517 => data <= (x"181e9149ece5dd6c", x"a4f1aa8c6acf5ab4", x"d1491d0458756a39", x"5faccdfcc12fa381", x"e1cac61bfb19c36f", x"d40ac21bcdd6ac6c", x"4e9d4098d7636248", x"a84fb96f51ec83d2");
            when 31660190 => data <= (x"965eab974e53a1b2", x"0ad21eb4ded9f727", x"13734073f1f0950c", x"1eb67abc3f54ab00", x"f815ab71a0e2cd4c", x"3d7f0ac1d48457a4", x"1a6079af0607bd39", x"bede2cf3378c1e68");
            when 30673287 => data <= (x"1bb258d30f34db4b", x"22f6b2201d46c2f7", x"9ba1062a649f2377", x"26e8987192d96f0b", x"e9f2a9550c8c4d42", x"49706220f27e6086", x"e92151394d5f8ee3", x"aa4b5ca288107026");
            when 12006613 => data <= (x"014c6ffefe2041ac", x"8649c03da539e753", x"93086d2cfae6691d", x"31e0219a48fa50af", x"e64024592f66ff27", x"0fcaa30eaea365c1", x"f493419d5e5389b4", x"9d13db3b34a927f6");
            when 21111659 => data <= (x"1197648fa96a2ab6", x"f1e7ae9e724a1f7c", x"9b1628abd70d000f", x"c8439cf64d273ac2", x"4cee31a547cbfcd9", x"93432cc33702c782", x"a224b72274406243", x"52b200db460d4183");
            when 31263773 => data <= (x"b895a9b92a5efe85", x"8e0e7db19df6254e", x"173ea3653cf01ada", x"e946959d53a5dd25", x"67f9487b79dac2dd", x"405ed2d0d0e90e07", x"52385024b41f2829", x"4cb71c8f7bf425f3");
            when 23618171 => data <= (x"373f468c5297530c", x"9c50e523946a366f", x"6c4bbd7c8d3070d1", x"875c59dc2d2e87d6", x"8dbc9de2c9a97d38", x"df6ca4dc32dbacc1", x"76f293e21d6fe20e", x"e85b5a330ff40409");
            when 18039808 => data <= (x"8ffc9d2aa5ea5b72", x"5042f087a4e7518e", x"0d40563d91d3280e", x"765eb2af3a8365e2", x"d4d44acdfd21cf3d", x"551855749274ed87", x"6d04ff0021a7ab21", x"ddba312fa9312882");
            when 11070939 => data <= (x"696c262634050898", x"2d4a09be2276bdd5", x"d3fd8cecc29383d0", x"195da8655a0aa871", x"c684937e77910e38", x"773c0255ef810c9d", x"f07d52f177daa6d5", x"268eb35ec3057c02");
            when 11109178 => data <= (x"9c73646004811764", x"4bc56904c66250af", x"a42cd625093c4a62", x"2e4526140f3f96b9", x"a1bf8b09f6219886", x"1529a2469acebfa6", x"4efa4b055d59664c", x"c008a905f3cbd91a");
            when 20382768 => data <= (x"7e231dea041e9473", x"1775370dfbd5c268", x"fd225465b46718b5", x"13b18b342801b1c8", x"3bc00c6073fe0752", x"910db2c6000ef2d9", x"a9d72791d22e2eb7", x"88551d3bff52e149");
            when 26742418 => data <= (x"9e8f6d215467e59b", x"71ff8156b1dc03ab", x"eb7de23ba31cb0b9", x"452d40e5dd7d2ab3", x"b85d6004daf8c827", x"e1db05ab5cafa349", x"6b6026b54ffb52c9", x"0b068a2a24253b04");
            when 6314328 => data <= (x"b3495b6e172d2731", x"21c8c29d225fcf77", x"9ffd39260e44b5c1", x"fe65f6fab49453dd", x"de188e3ecfb122bc", x"559d44eb6b70b400", x"67e8b95f1a799d87", x"462968e49e4cdbb6");
            when 25370360 => data <= (x"ae6a29e5109dc634", x"1e8f7fd25aea7784", x"e47b39d97f2755cd", x"7fcf5068c18918bc", x"68db5d8e71302068", x"bab0ee62851c193a", x"13e08229568022cb", x"d42c3edba3a44ff6");
            when 17193027 => data <= (x"3bc1d06cee610077", x"32788f7f9a8e8442", x"ee893eec57590f9e", x"fe3a35dce7123f55", x"59bcbfe370683156", x"0e93f46fd422b9dc", x"ba17ee186ff9ada2", x"5c9d4cf3c1d45bfb");
            when 13101914 => data <= (x"2cf8e425f32617cf", x"9da022e02f166694", x"9326f9c3249e818f", x"167b8d33b1b3f7a5", x"1677f16fa53ca9e3", x"9d036b9fd4a84bf6", x"360388fec70b37e4", x"258bc3be1f8feeb2");
            when 10364951 => data <= (x"aef066571047f2b0", x"dc4d817afbdbea0c", x"01bc05e50f0a6d11", x"0e77aca88ed4c57c", x"26a66488584a3b84", x"7a14bf7e75088811", x"2832936e8c317bdc", x"43701b19152697c7");
            when 18637743 => data <= (x"3288e5ed24d0f110", x"03811d6311301921", x"e2eb7d5c08b77a72", x"c60173197d288963", x"a8ef941524912b3f", x"d3a07e67ad75c50a", x"3ba42f1499c8bf3e", x"5b8202a68be108a7");
            when 22679698 => data <= (x"8cb40b0866e315ac", x"f6055aede34b0c6d", x"abbf83be90d964d2", x"9fd6f4ed67128d56", x"355a1abf1d682746", x"9f1ae001eeafc92e", x"5a7684b48e089685", x"dfcfff4f433ff0e9");
            when 11952361 => data <= (x"2fb5c3fe36d3114d", x"9886ba6e7b108a85", x"38533899c702ae8b", x"d3e782bbf19fb1e4", x"4b8a8feb345e0d74", x"35a85e3bee63a634", x"9c33a8bcbe22626a", x"df5c45d20440c7c0");
            when 22609912 => data <= (x"e520a4de9f0e773d", x"67cc0c1899054d8c", x"86207ed9e503a448", x"e3630782938ccbed", x"eb42bc34e72d6913", x"dbee9a21153764a7", x"ac9b5b865b4901ca", x"423cc1b6b68fde8b");
            when 33348801 => data <= (x"011fce9826148cca", x"4834b99046046636", x"a11b17cb89bcfaae", x"9a78f5cd0c89e4e3", x"0f26792fe24db336", x"e0c5caa77f9a509c", x"fbd8261ea8d81d1c", x"f758342d3a55aa54");
            when 13129127 => data <= (x"8fab6fe0cdafe618", x"565aba08c2dbcf5e", x"c20e97232bab99d9", x"e75697f21ff91d5e", x"b5f4c8bc30319d17", x"728897a1a105980c", x"1be83690452fc904", x"2e1c095036516051");
            when 7287910 => data <= (x"162d9945cdbbaee1", x"6db0a1c4b07b45db", x"6f583825a3ff51dc", x"6c527f3de6326d3a", x"13c10ad18b210006", x"85ac669dc1559d32", x"1807ffe764cfdb76", x"0ca80d5dc0e43c91");
            when 27179684 => data <= (x"ca35f6aaa8dd05f0", x"6b37403268f92e2d", x"220c6fa783fd4ecc", x"6443b289e1b9e58b", x"51ef0b3cb1acb633", x"a803d540b998d448", x"c909fa66be4355fe", x"fc3be7e3716296d9");
            when 8173752 => data <= (x"6eaa1ec70d045fb1", x"114d8832ecc7f8f7", x"f7a5ec7df5c94acc", x"fc0cdf664100de6c", x"097d72e07cc134db", x"8350a7c4b60e37f5", x"b5c5d232e46f9db4", x"ffaa061d17ecebb0");
            when 22752854 => data <= (x"e9fac0eb688945d1", x"6b352b5416c05009", x"ab819c0d7ac2c94f", x"dfedc246a3f8de16", x"c9ddfaea12228b84", x"1d6143da476cb776", x"c4c61bf21f9d0601", x"022ead9cddadae67");
            when 19271597 => data <= (x"05b21d318b6f771c", x"ccff80b4e7ee3990", x"a060abcf5e17e0e7", x"fe3f8a9f0dbe577a", x"95d65910e2add495", x"90f93bd935d38899", x"d750e434c80b0406", x"56b1bde762292636");
            when 31504256 => data <= (x"a5c3f7c23396dc82", x"1e751ceb110e5a71", x"becc2d7c900b521e", x"2716786e383c0e88", x"fce3ab3aa8ff6b5d", x"7f2ad152805ba0de", x"9ace3c22f916ca7b", x"507bae0c35db7d79");
            when 30850357 => data <= (x"9fd56685b52c889f", x"41d3488f48ffa5f2", x"f5b14df271f3c45b", x"94e3d0c6c4c30475", x"e2a9f9489ae4b70d", x"4d320336be2c0889", x"eafe6d7febc80f96", x"3a807085c332d45a");
            when 3490453 => data <= (x"46b09601467e78e4", x"51c952a96a3a2e81", x"be670ed2ec4f2179", x"94e85941ab4dbe50", x"18f82c595128ad1a", x"74557c6f5374a214", x"27949dd478b0d8da", x"6f6d89c1b5fcf106");
            when 31844522 => data <= (x"008abe9d9dd97983", x"b7e65fece24586ad", x"5afa4f074c8b8118", x"d9b67d52e0f4c26e", x"07a1f23a45f3b8a6", x"205eb5cfdfba27c1", x"0fe21b93ea1bec02", x"51df4951e660b7e8");
            when 6265487 => data <= (x"b84b33b4de0f45c2", x"db1e17fcf155d190", x"1a00cffefb4ae90c", x"3f5da5c39e012bd0", x"59cd1255c8cc514a", x"f317c0f126721d03", x"0a655b0413812ffd", x"fd458315a91c69c9");
            when 10661319 => data <= (x"d61364f79530fdc1", x"41bd4aec466d3092", x"58a626e7a832e541", x"9e34b87186236ddf", x"60e63d5ea1e7f6f5", x"2bcd78b7da9433d7", x"149a704961a2cdd2", x"0eac77d6002b04fd");
            when 32853738 => data <= (x"f07c94835fe92792", x"a320bb66d624609f", x"25c80f925106acfb", x"6311590068828b76", x"e0d776edde033db2", x"4e501c4cbf81b395", x"2da60a7bccb590b5", x"464eb60ab8eecba4");
            when 21411334 => data <= (x"a998c4b777ceb383", x"3d16e739a7199a1b", x"f1057001898ef0ba", x"ecb8d57f51ec331d", x"477cea502e4c5151", x"8f38e158aa359493", x"15d146e657e3cf70", x"02a2ba901f1b501b");
            when 777383 => data <= (x"179293ab13d04665", x"30dc0a6b5101f6c8", x"a46488b2a96d7744", x"39dbbb5e620d83b0", x"a59952878e83f271", x"fb615a58a54dcca3", x"b11a65fa8dae2dd1", x"8c4484874f23e8c4");
            when 6601382 => data <= (x"bf229ea0e61bc4d1", x"bae7a01a4b409444", x"b83e7cac81c7d43d", x"22cbd16e6d8429cc", x"fcf08c293763412f", x"00fe2c999543e6e0", x"301eed69caf0be2f", x"d0cca923df5df4a8");
            when 7123204 => data <= (x"f7affa8e9ac4895f", x"c784878a22f44a55", x"4359666bf41ba9b4", x"2de5d612057d7fca", x"9f3f1fd94c80e4f4", x"ac22bde584a1b69a", x"f61815c9248b7c57", x"01bef19fc3dd551d");
            when 1575025 => data <= (x"6f216aff90afdb19", x"a52c61119e7a0949", x"01056589d00d99ec", x"dcde7f730426a9a2", x"c1f0d28e5823c03d", x"1413550a8a1ac656", x"fdecd4b526919345", x"b8e1ed6c573533c5");
            when 6285834 => data <= (x"06102c221b260a27", x"16f13a1a0c819a2f", x"2a808d7085d58643", x"03d4a1d65a3e8d5d", x"12596405019a7ec5", x"ae7d54cf000043c6", x"a9362aa47414ad8a", x"4a34618d321adff6");
            when 21730937 => data <= (x"355f595482df541c", x"41858c08bedc69fb", x"43652e6db075116c", x"3c355d76077e844e", x"518ff7759cf409da", x"7d1afa9bcd1162da", x"bb64b4cf50e755c1", x"f4fb44832caeac94");
            when 29831261 => data <= (x"b57337cd46089d51", x"bc2aa700ae6e93ba", x"196c53f64e3b0926", x"ddbca0db812cef35", x"3bef9d5db4aa8c06", x"e875acef9da8283f", x"a3c5ddceb85682a0", x"645b5b9695cb6d75");
            when 4966434 => data <= (x"cdbcdc57c32c7a73", x"b478acb7d610f8c6", x"81cb6d2b2d937949", x"1ec5be4f01499d31", x"12560735d83c8a75", x"87d905ec583456ff", x"2542a6784289e73e", x"d7c106adb8ecce78");
            when 4628484 => data <= (x"7a476021bc1a4e5c", x"3407beade8fc398d", x"34468d5908618b6c", x"a499f39e811fc95d", x"02ba8cfa0bce22da", x"ed96018e237467db", x"38675447cda02fbb", x"24ca94a3c8ec9a7d");
            when 12490857 => data <= (x"dea62a1af7d84923", x"98e36a4bf91a0472", x"599925f2ba10903f", x"3912e04db4a80f8e", x"3505c6e25bce1cef", x"0bb9a0be2d242d64", x"583a6b8ddd331946", x"dc88d6781899b731");
            when 20049691 => data <= (x"539632e00279598a", x"4e3663a413cf08b6", x"6cb431ba65df8455", x"58658bb53bb72319", x"400581e9cd64cf01", x"e96d4662d2c9b9d4", x"2489bc0afde93cd8", x"ad1e64099bb9c6e4");
            when 18486452 => data <= (x"0f4aedb4a55ff8eb", x"58326c5e8b462305", x"48c2ed123b8cf234", x"9812a229d5dabc47", x"f786001cf3f044ce", x"b59982796d3739b8", x"93e34ad5597c5112", x"a9d0d51ac1a716e0");
            when 955975 => data <= (x"8cf811c70cab00cd", x"ff84a0a99f97f62a", x"e5930693c908ac67", x"4015096ff8277360", x"05e42707cb8fdb5b", x"30768a3b8b0ca5a1", x"732b1f8409d67e10", x"8c15f3d033b56e87");
            when 16658802 => data <= (x"802d5c62fc0b6cad", x"90e690952b4ac0de", x"d20e0420fe8a5219", x"7ae8dc03c0924465", x"6691fce05ebe474c", x"bb686db3d9fbccef", x"e134c9a785518aca", x"1d78c32bc7994bed");
            when 16032159 => data <= (x"6fe7260f10390c6a", x"adc07e06d5381a21", x"e4484fb0944445df", x"ca3d762e9b253679", x"fb973490b47b8f80", x"8c11b49a181e5d25", x"5ee433b92bfb562a", x"2e416b8d9f76c266");
            when 27485268 => data <= (x"8ddf894c0fc05ab9", x"d9f41d13ef2ae7fc", x"31548ae595f29959", x"337faf3313cf6e92", x"9c622813762a34d8", x"7c3ba12b2285b443", x"9304495e8300489e", x"f5c87f455e4d4f32");
            when 30308157 => data <= (x"6dde42cd194a42f3", x"1192e65081f4cb14", x"5f0e1405cfdecdc0", x"f5570d9283682e9a", x"76eda2654f692a76", x"af7007f31a69ce4a", x"8f88bdc0f731fd1e", x"35d51c6f5d581c51");
            when 18308297 => data <= (x"b0d8155a4efaa274", x"9534430d2b805360", x"e196cbc3b43911d5", x"f5e03126b726c1da", x"02b641d8161b0a3a", x"1133f344c07d007d", x"756bad4b40eb7844", x"ded04887159ef388");
            when 5417761 => data <= (x"5030a3c13b0f0e17", x"a31ae4025ee64f59", x"39c3ddc35b1858dc", x"c5eeb64f4433920a", x"ab7af9fcb3c69d3f", x"0d7c3ad96e60e1e6", x"09a3f01baf431b69", x"698591f8329e0819");
            when 10784558 => data <= (x"d2094c700a18b4f9", x"58e12c106b9a02c9", x"edec36ed1b74bd02", x"1c3100de899e3711", x"2987449e75257ddb", x"1c0a04eb8d82fcbb", x"7503f54b0cffc961", x"c71a1c0f0fd578a1");
            when 4711116 => data <= (x"88555aef731417c5", x"b208994f47bcf322", x"1295a32a07486e31", x"aa9cad9fa1cdd75b", x"09c1e7ad4d649862", x"80027756715188f6", x"f646309cabcb8844", x"6aeeddce869572f8");
            when 15741316 => data <= (x"4e0677d9a129cc70", x"243a41f03c89248b", x"e9577919cc915d91", x"b83e6c48e89ede7c", x"2543590b7d4545a3", x"dfc0562986f2115a", x"2194d8ff1f05a142", x"d28c840ba6a1583e");
            when 16095327 => data <= (x"7e29ca9de370076a", x"0a6ee69bfa64bf9f", x"0e76fa45b175b8e9", x"9a26d82602c715b3", x"8025b7239e03dc11", x"0b20ea420f4f394d", x"f7e8641e93332113", x"260e5da94a2574a0");
            when 5134512 => data <= (x"4a6c79f9f8b161db", x"950cf58aa7448bb5", x"ee195ecea91c2cff", x"65cef39d0f7e0069", x"74f11ac29647ba9c", x"d0876e08a6ee0fa6", x"814b5400fcfc2c2f", x"849172a9334af7e9");
            when 8821820 => data <= (x"266e248f5923ab79", x"3d5340045272fcd1", x"92159b3e8d9c4266", x"bb40c905a97f0373", x"544aedd4bf97d9e8", x"f3a169b5498e351a", x"0a240155064570ae", x"c02ed13d48988ae3");
            when 22092788 => data <= (x"247e24cb8d794cff", x"d571aff53454da17", x"0159206b4b4c684c", x"b6175f4562d72b18", x"08239904e8ff569c", x"0b954cacb732a7e8", x"9ddd308be7d3ca5e", x"b47f2b09c273f8c4");
            when 32317898 => data <= (x"a513c9072de0c98e", x"6beb9e73ba8dd46d", x"6241d81753d00ea5", x"786f8e54a6f621ad", x"e9dd685b03e7ef32", x"8615174c497a6cad", x"463604f3e8357703", x"91cc0d03421522a6");
            when 5472375 => data <= (x"dd6c95ea652dcf39", x"80891dce561c05e9", x"10c609953fdf27fe", x"c26caaaf646a7c81", x"fa88f9b1cc62732e", x"ed52be2dc6f4a700", x"008f14196d26447e", x"e807cb85cb51be80");
            when 27253347 => data <= (x"d2e110732b3bd660", x"ca52e50dfe73db8a", x"14b539e752417238", x"76bfbff3bf45324e", x"1e4478439bcf07bf", x"faddd238f5b9ac51", x"f5a43636c6c7b446", x"bf7385aa73c84ff5");
            when 9379812 => data <= (x"6a2f12ca8835d4ca", x"f0ba93eb4765c6fd", x"207e792ed7768d15", x"4ecd511394f43f56", x"e5ce6d80b4efb243", x"016f0ba25bc124b5", x"19929711b4cc1ca3", x"e6e089503ca271d5");
            when 28204884 => data <= (x"01b550b74c4dbe5e", x"4cd731dabcd9928d", x"782b6abc8b39cddf", x"387ec88566eb5adb", x"e2156b00512786f6", x"aef3de14091601e9", x"bc4bcbf50a13ddbb", x"96b915d8c41e3193");
            when 30792607 => data <= (x"be58c273ba3f0d28", x"8fb3ce97a2266ed7", x"af5493aeeaf21e95", x"6eb31cbc150e0e80", x"2657b6f5141c4c14", x"6699c76354cdd98e", x"07abfa88e1882a53", x"0a0e71faf42ba216");
            when 1530783 => data <= (x"96b395ed0afd4f10", x"bbcc201ed08e5138", x"47e1b637a7784368", x"2b64026ccd8ec4a8", x"01a1094fc70df7c0", x"720c9c8916dcf0c4", x"e67d10a83e1b007c", x"c72eee9cc806f916");
            when 17545728 => data <= (x"4068871658387a8e", x"6b2be45eebc3bb29", x"5207f788b0dcc47b", x"94617044541ae710", x"280c651ded56cf6b", x"1f85a7e4c31a70e1", x"01875f6d1cb005e0", x"7c00c7ad971d4fc4");
            when 15546068 => data <= (x"79d3679940d2acf5", x"744932e411e0e494", x"302243a831436a83", x"7aa7300f9677efe5", x"c367b29e1c026a8d", x"11033c7fd77d727e", x"6d101984e5c3e424", x"74f2e039f1644c46");
            when 20497508 => data <= (x"ca4322993f4ac66e", x"47707e6291a4278c", x"c23a65cd4feca7d7", x"2c376164a2d9d424", x"3470b1a218885355", x"2708757b9561dde2", x"d746d204a9812c37", x"08fead0c95afdcea");
            when 3101847 => data <= (x"d1d52a0a1dff4e39", x"164f090b2ae2cdb0", x"328ae3077b398fc1", x"f56916f10891f0e4", x"4bdf24eaa60dd2e8", x"b577c077c48832c3", x"6913039bb4df1d55", x"ddb4596326af53ac");
            when 14833478 => data <= (x"90e5189688538710", x"3eecd4a26f88b5ca", x"3b6b22cc46c82156", x"0e81343c7e72e596", x"f178ec550876cd7f", x"bcc78762ef896e00", x"ead859db9a05e129", x"f14b1a8e6f7160e6");
            when 24695771 => data <= (x"02857357aa0b7488", x"e51bbf8b53fce1b5", x"cc745df974c4a43c", x"7762a448995b698e", x"cc00feeb387bf64f", x"1ab8e3a735286f1f", x"1aec53f03eb2057e", x"d6b406e1da2102b5");
            when 22456716 => data <= (x"9fe6c45b0108d3e6", x"3efa0f7f7a6d7b55", x"3d031bfd6e2dcf07", x"ca89b5b6d3922c8e", x"b401fd9f9998c133", x"be8715bef6852bb3", x"4031a47e94cfd2e9", x"9c0f9766b7573730");
            when 21733619 => data <= (x"34b1ae68b4cf9b6d", x"b78e411b39afb69e", x"a2ee2572089a88f0", x"7666da9e0bb41101", x"0ed9c7e2c75dbf86", x"61e2e1419f0f82d1", x"3ec010e3c28c1786", x"2dc58f0831557c1a");
            when 3345309 => data <= (x"d0a2e9f96743b7c7", x"affe59eafd778bf5", x"2b3f7bf2a50a8129", x"ce0a33be735559b9", x"3a3b84bf2b227404", x"357d15c3aeb74d61", x"1ca0d0fbe4341b99", x"eb3ae509d346febd");
            when 27264631 => data <= (x"30ff573991790df3", x"971570ca39ed91a4", x"62d03e9d99474bfb", x"15c8134ae7d1f97c", x"1810a8318e8de1b4", x"7d99625e9adf82ac", x"f9c2d4c97875dbc6", x"c42ec49002b70436");
            when 19345944 => data <= (x"e5e3a342d61cf426", x"4ce6b506a9e17cb2", x"cc7eec4d03274023", x"c1d64bb06f624ff9", x"63b0f9fd256de53a", x"35c73d4e31ada962", x"9f30eb620a3f02fc", x"81fa8e5c7262def0");
            when 3775833 => data <= (x"860c214e96951a2c", x"30343f16a76bc25f", x"9908a559a976ee6f", x"71aab9f3f8603bd1", x"1086d6161c699729", x"98170d92a101c354", x"2f4932286a40a284", x"1baf5f5f666c90df");
            when 13397616 => data <= (x"109c5465f9d9691c", x"ec59849efa077dc0", x"4fffcfffca55bd12", x"a7fcf66dd7a14708", x"f178ce829cd8b433", x"671d8331f09ee61c", x"51e83a0809cea509", x"4cc3fd57c8e5bd7e");
            when 22649470 => data <= (x"c702193101a3c3d2", x"b838a69b57ead917", x"7736a32d953a2192", x"8a34dd7b5815ebf4", x"a4370442419541f8", x"790ea09731c0c22f", x"7879518e00695318", x"23025633aee862f1");
            when 2289694 => data <= (x"1ed42a7cd2c6b21a", x"72ad05425cf251a6", x"ff53fd8dabf6b58b", x"57ee652975551de8", x"859d7bf6f7b55c0f", x"403a31b57e532b50", x"0b1a687e49bbedb1", x"59d328855eb4400a");
            when 2262034 => data <= (x"d8f90a97e7e9227b", x"d8a2f76c6812fbff", x"4917b04ac7e81a4c", x"2e1fb77f276084ec", x"c87b2c52546dfba4", x"3fabe1fd9cc6a886", x"ae81669b057d5bee", x"84f4ba8e8d325a36");
            when 21947325 => data <= (x"4ac1509963f4098d", x"049d938e14b8038a", x"0750862c041535bb", x"96648fd1847afdef", x"d7f60a1f80f42989", x"7595387bef06c11f", x"9d3f82c8153423d3", x"f73c7f970c8a1011");
            when 29552100 => data <= (x"37294d67a4a1e516", x"a03b15d22da8f0c3", x"ee385bf2d6aa44e0", x"3480b1ade2ca5452", x"607d4402bbe2966a", x"2a3869032e3e6531", x"cfd38bf39334befa", x"e4b9cab22d16af19");
            when 25938793 => data <= (x"1b307a39235660eb", x"18a84be02e6b8ddc", x"a74e52a21e7a96d0", x"1997047decc9e84f", x"c83238fd81b29466", x"1fb91bbb5176b810", x"de674488f0a4224d", x"d8038171e033af8a");
            when 11869752 => data <= (x"e338a42ef0145080", x"80e8768ed381526c", x"e6104af48150dc1f", x"7c00b8c7d70db097", x"0286735097867c0b", x"b2f0f67aca4374c1", x"cb621065bb779602", x"9fa0be0e923f9b1e");
            when 21294305 => data <= (x"7c173bc6c4e63728", x"0840de1f53ac7fe4", x"f6643026a80d426d", x"608af6a04a1c054c", x"94f6742c9d79452c", x"5c2c3f0eaddb4c5c", x"1dd9a3e74f14d1f2", x"198981c5f10b0327");
            when 23561965 => data <= (x"a256b7bc21d76e2f", x"eb952983a721280a", x"9955fbe3a627b933", x"299ca5e5c85bdd23", x"0d33783b9bfcf5e7", x"7e071a9d7d4138ac", x"10bd2e5f77821ec8", x"59bc7e9860949f4b");
            when 23788073 => data <= (x"033cab98435c62e4", x"7e69e4647ec71cfc", x"8d5c4ab420df6bfd", x"e096125943c6b145", x"11995bcadc41abe3", x"0500348f866b91a7", x"40889a1de3f4ed90", x"33c33448518592e1");
            when 22728950 => data <= (x"fc0aabfc2ee4fa48", x"06f026f528cad557", x"fe1594781ef525a3", x"39b20f499eadbfee", x"07b101808ad90f9d", x"f8bd94697ae48a10", x"78cfa51a41219ef5", x"3c161dcba4752171");
            when 10351714 => data <= (x"0f0e5b47d9477c5d", x"26af7bf986b2810d", x"e9d5afb7750689e8", x"00089461bd29d813", x"3331e3ad14a01465", x"cb9534caf3d800c8", x"fe126c39f501d3a3", x"85d27a56ecf78fd1");
            when 5028446 => data <= (x"45e3cd493240a605", x"0db411ed6d050974", x"24e072ecd5a4f1d1", x"fcc9a2d169b49a24", x"577cd99a06e63f5e", x"0f3c253cf0921acc", x"441c2a0853dae1ee", x"e1d8bd031040493d");
            when 24000382 => data <= (x"0d8ae78d0247e599", x"108e9fb2cda34c98", x"bd9e3e3a38d47962", x"8d4b474188b20d38", x"7cb21bc9a55ecda8", x"85d4a08868975b83", x"a092aa4b52fe8906", x"4385fc217e352388");
            when 30157653 => data <= (x"c2d83d6b75de4949", x"cd0886bda197ed06", x"e8c48503ad07f9dc", x"1844733f188949b9", x"7e934bc15fa7e3a6", x"6c7f64a7be6ce00b", x"79da2a3e799a1f74", x"8858ed6ec4626231");
            when 21971891 => data <= (x"07c2ee640832c144", x"385d022d9e51ef08", x"5bce1b9dbb05a3b5", x"cc2cf3975452c853", x"0ed6adbef143a170", x"8b28d4790dfaae62", x"99aca7134e366af0", x"fe3d864495fe7059");
            when 5968797 => data <= (x"0e4fcc85abe7f843", x"2877e53765004d13", x"986aba8e0ff2c879", x"0adf5727e95b1190", x"2d81398437727933", x"cce98426d33f0b4c", x"d6cab1b8fb218aa8", x"1d52dd2100702c4c");
            when 25686627 => data <= (x"06c177bdb40fd2d7", x"b5f7dfc023ad7a0a", x"f50aa45653079b42", x"3763856b05d809db", x"ff974c4608ddcc93", x"dcf00f5c9daeeb18", x"12708a3fa725bd63", x"e16a5e8b84d06cef");
            when 30211389 => data <= (x"6706c6f0ce4e26cf", x"b368215f4778deb5", x"ea30cd6fff1394cd", x"55a97c5437624d1a", x"2a71e27a5544fb56", x"f0d224dc1d1600d1", x"3411d916c77a5554", x"fd8f6b851bef3f20");
            when 16477842 => data <= (x"b1f0d368193446f2", x"1ff91db3d14e6736", x"5c3a1997dfdd29ed", x"07f18b463d41710f", x"f260821a39eab180", x"85aa09b6571720bf", x"caa8b517bee8c219", x"a83631a26b2a7674");
            when 20014417 => data <= (x"c09e3ecf1a1b8ca5", x"4487ce6acf44ab7d", x"99bdb24cfa6981b1", x"4dba9c8c038ab397", x"04966a45790add60", x"29dd4145ed5698eb", x"929e76bb68de2aa1", x"e6a7328cb5fce0df");
            when 3104905 => data <= (x"d38cc45758463d44", x"45c60d4343ccdf5f", x"46dd8142992451e4", x"fbef82b6e903049a", x"8dbbae9f0030cd5f", x"f0b69588ddafec10", x"028a5297989ca25d", x"a22124e764761d03");
            when 23950933 => data <= (x"b3829af8e04a19b3", x"66d691c13f535f19", x"60b8f31ece203a9c", x"9516d75d806a6b44", x"4347b2cd8b4698c6", x"aae5e6b5957598ca", x"cd49e0e3f94b633a", x"94eac096e90e6f7d");
            when 1444815 => data <= (x"dea17d929efd1cf9", x"e7dcabc44b4fb4b5", x"1182d0605cff7fb5", x"cdd2debd0c45190c", x"906250dd4bed8666", x"6de4ebeab9f0c855", x"99f502cddf461703", x"94ad666fc278c2cc");
            when 6403465 => data <= (x"cb02bc08fd118786", x"220021c7fd528d1d", x"f20ad58aa88a48fe", x"3ba6218cb36cd479", x"96a1fc9ea694b24e", x"b4084c1fb1887304", x"3d1c10266edce476", x"51ac85befd6d73dc");
            when 15881658 => data <= (x"1c5e41219b41a0cd", x"d5efb3ffad90fd9a", x"9a154757d7596bd9", x"45b3e160c811b6f6", x"4b0fc32119e8e1f9", x"351bdbfa8bfe4547", x"8c107e1034270839", x"e49c394d7c56d3f2");
            when 1988657 => data <= (x"7835599a7b734c7f", x"c1d521192484bf40", x"a90a2cdf86e84522", x"251f8cb2ac429aa8", x"5a982b547c97df25", x"39a995c01e474637", x"3433011fd696de0f", x"9fdb4b2170d27f90");
            when 27804449 => data <= (x"b3096d3e2d0c79fd", x"e798d34cb8cbe8ef", x"69a57a249f7d8bcf", x"29017dd877eb3205", x"19e1873d05bdfc1e", x"6c6304bbc9fb8a42", x"00ab35b6069474d0", x"a9700a2d1e3cf038");
            when 9639850 => data <= (x"56a7bc3ddc6573a1", x"d7986fb9dd32b3f3", x"305bf181d15de416", x"3c07e263ed02b668", x"83e1487e745d1cca", x"1b3145831e9b0407", x"76c9a651764fae66", x"cb0dcb12353ce022");
            when 28165728 => data <= (x"6564dd133cf16b41", x"6dc11850eb753f22", x"8d14c6745198af00", x"b52dce48f02be34f", x"c9cb2d9deb631d82", x"60b4a65bb433a27e", x"4eeb3c35d069beb9", x"9db1de1efbe1239d");
            when 33112751 => data <= (x"d6726b16bb2c24b2", x"8edd80db3f7deff5", x"819de8d393808fe6", x"757485e2022c189e", x"28aea85d7de6a943", x"e3e019aa410c5f88", x"33b1ce4bd1ef7d98", x"9e4858844427466e");
            when 13623203 => data <= (x"195bbf7697d35ea8", x"f4167676b64bd7cf", x"bbd1fcef2cef53b9", x"449959c8dd54f0bd", x"300cfc34a71f3e37", x"e554c9139f6ae33d", x"e9a2edf838b70fae", x"ccfdb4ec9f6e50ee");
            when 9871540 => data <= (x"90a21189ffe130e8", x"186bae1124c83e2c", x"9c3f4441a0977ef3", x"3651b42a86b4ec30", x"d145b4e2c3b0679c", x"bad71c717f5a36a9", x"1653a8585fac4e5e", x"883d5d5f02b3249a");
            when 5107640 => data <= (x"ff2fff33644e5772", x"a627689b90759dec", x"1c6adef6c1589261", x"fa48ab3873ac7e2a", x"de9c3988d768ed91", x"1e3de33120b7b78a", x"79833e4123cc0cd4", x"ccfddd64b658e5b1");
            when 3832390 => data <= (x"3e1df542bbc5a40a", x"abfd360056d9be16", x"85d093d380a03fe7", x"082b34b197dbf0d5", x"2615a2e80621d44c", x"429b952b30e6720c", x"fc81079970217b1d", x"b41fac0d848673de");
            when 32428703 => data <= (x"4dd5d494831b7738", x"92b2459a2fe3b280", x"4b2e0e940facee5b", x"99dd747ee693108d", x"6527bde7d60bfe7a", x"a54270f26b377e52", x"a20dbf58453bb721", x"9f6336a1633693ed");
            when 14667287 => data <= (x"f7afe12f8a23dba6", x"81e9c3452d28d820", x"b092997f3180f0a5", x"68dc9aebd19091d4", x"ec59ebe53b584afa", x"d8009d88abe2ecfd", x"f1a19694c3e1e0cf", x"5206457bc6498a67");
            when 4821518 => data <= (x"83adbeeeca5aa0ee", x"3f14c34d54eaf91c", x"86327317d2d93857", x"43a7b453df26a85e", x"c60ede5388f12aec", x"2342c70a5904a512", x"354b77ec4eebd708", x"33703c9eaa017406");
            when 12652246 => data <= (x"d509ae2b45698822", x"1265266b89fbbe97", x"77d2c265b164255e", x"c6b37b631dd945d6", x"17e2b73c99768610", x"332d35543fc19170", x"dabd68096970ee30", x"6a39132f2886fd9b");
            when 26365332 => data <= (x"4bd289962bdcfb7a", x"384b839d4cc8b747", x"d6d8709237e9a9b1", x"0c66059ea8f2decb", x"ceb45374ec5fec83", x"1af756e814cc9d4a", x"d4303941987dba35", x"b65b458c54f94e5e");
            when 14855357 => data <= (x"f2c1157a0bc360ca", x"070b9827fc0f9b9c", x"c42ff5238542e944", x"ffe7f4687f21b94c", x"6cae7c093a902e02", x"f5bfcded87a63074", x"42514d15f03c92c5", x"ac43323923164ebe");
            when 18747801 => data <= (x"5b57a53fe5df75c4", x"53878ff175887de6", x"f6015f6356435fdb", x"f4d847b708722480", x"ee892b295284b9ba", x"97933db4c2dbc8ba", x"d380fe21bf649b6e", x"29c1a00faf25bf9f");
            when 7454448 => data <= (x"7f9a81d3848df11d", x"323dfafe1280e208", x"d241bec58604c0de", x"246eed2b1152be3e", x"6565c18c15167792", x"f5fcb85347be6ea6", x"8db0be78bea573da", x"e563dd531493e983");
            when 16999121 => data <= (x"514bf4c6b00d7c20", x"f85d4664401637c9", x"f948a5a52e361755", x"7a476d09aa7e2551", x"7446e6de30226abd", x"ac89c373648e4062", x"264a4f55119f8e7a", x"6c55541658032c92");
            when 752256 => data <= (x"c5f0b59073748ea9", x"7ec5f6bbf4b600a5", x"fa5e7d7c4506a50e", x"36c998beb26b6a54", x"7a7d9e5ba5f3b825", x"e2b13477290aa6e4", x"62d2e62cbe64cf91", x"9765f8cc8e7b0811");
            when 5141548 => data <= (x"6eed03f06352828c", x"4623903bc03652b2", x"5543729893a3e55b", x"1bb5da8ebf26bc9b", x"606abbd649265290", x"32d2d17d320b29fd", x"406ce690c5b5fc31", x"19a9a5b7ea79353d");
            when 12725669 => data <= (x"298f71554dcb83b6", x"070fdcb08c2b55cf", x"9ae9eea98b0618fe", x"3734cf478ba40800", x"388f8fedb69d4a79", x"bb6d3facc09e19fa", x"1aeb4e7d488db073", x"bd8fb4234ca7fa26");
            when 15938278 => data <= (x"3a4b7f20c1dbb7b1", x"607e0cbb7ab3296f", x"fd696c2719628aab", x"e4e3643060567065", x"56a2715a8a36f98f", x"cba14d6b2f0e6e0c", x"c0b715d3038e0ed1", x"93184ad0ec3737e0");
            when 21490583 => data <= (x"9fbf2d16846c7c17", x"4abd78a074f7eebd", x"5d653bdb758ae7b0", x"d334b9b0319ad933", x"9a9e83f1415632ec", x"5446698d7a29e308", x"f597ebc5b7d08b75", x"95e24a4cca1fa700");
            when 14047136 => data <= (x"4afe30f678f76610", x"1d6c2ca062b918b8", x"bff50d44d5184f65", x"9e3147cce30e31bb", x"10635c18e95b7243", x"b002d1be34a6ba95", x"d2e5907eb88ba459", x"80a39b16c0106650");
            when 6220082 => data <= (x"a96551243db6319f", x"b795421bf43f720e", x"e8c5fd796ac7eb47", x"5e8d97d988886438", x"ba40b4874ec88e3f", x"b1b7edc319240573", x"06d1c63203a9f2f2", x"32cb7f833b24b553");
            when 8764089 => data <= (x"c747bc4680acf00a", x"c65e9a9037a2a8b8", x"65bc8aca63e14fc6", x"6e8c47370a6e06d6", x"1489174df9843917", x"bf841444e2e50e3f", x"d6148ea42d8c7c04", x"4cff861c43272f4b");
            when 705796 => data <= (x"e3dc2f18022f5cb9", x"44441630d4c559de", x"a6486d3246b61fb2", x"ed8269138496e0b4", x"89d9435c7d551d75", x"2ea5bece7ac33e5c", x"79660afe73c635fe", x"a231673a5177510f");
            when 13467475 => data <= (x"367243ef79a33c47", x"d8ab7c1353af1e24", x"b969f016ae86925f", x"e683b0b930102f17", x"8e50e09cf40087b2", x"165b5b445f7fbba5", x"9caf023e7251ec35", x"276992e0feabefa6");
            when 9486694 => data <= (x"7966243c0cb64c3f", x"fcde1faf0f99a510", x"d31d320f657692ea", x"aac339041f2fd554", x"eba09e030f937c27", x"0f3b49587dd6c672", x"5d311d9d32413aa5", x"65fe6aaee33c9237");
            when 29629081 => data <= (x"a1650a8c8c0d6ba0", x"70254327829cac53", x"66f7edfaed1bb13c", x"db284e5bdff70997", x"961ce6d25bac5413", x"984859156e905684", x"0fabcdc8e238e940", x"14213c3dfe617e58");
            when 19779229 => data <= (x"725e784797136e47", x"f2b6d310cd91b79f", x"087593f543b8f656", x"e23f409422c24c92", x"1048e6e86e07ba59", x"5921845313254e4b", x"c86c5c42242190b8", x"04159d546d2c1304");
            when 20541093 => data <= (x"62d9316a3c38e8b6", x"9a5ef886bd52c98a", x"9d7aef4a5c827866", x"f1967586e3347690", x"0bf6ea2b8d564d04", x"6952f23296e44b7b", x"ace0f9fe968a7b20", x"e2fec11e11d0444e");
            when 29342996 => data <= (x"4aed7d31a10823c0", x"ad43019670defd48", x"36f3a663b436846e", x"210398c4209ca9fa", x"d94312a5ef2fced0", x"d0770abbd84afa21", x"c45f61a96e834a96", x"3887864f461d028c");
            when 22342769 => data <= (x"6dfcbbdc4945d6a7", x"a5941195ca968eae", x"4c30c37245430779", x"d39de9c720bda5bb", x"9c3958dfde10d8ee", x"e2bb03e9139b9c3c", x"deeabbfb9713816c", x"0243f7f41646e07d");
            when 18833041 => data <= (x"1ab8e360e7fd9dc0", x"4deac09a3a784182", x"5a81e5efc1f86049", x"295fa1e059e74513", x"6974d36452897642", x"63f18e658f16bf8d", x"56b353d11cbc8e16", x"3b5ccf2b606cee84");
            when 32070361 => data <= (x"13d8b2829f1f31ed", x"816e5158c11df5a2", x"4496ddc2d107d8ef", x"2d89defc5585b7db", x"d1516cbf56c63d02", x"3ca89820ca5ff9dd", x"6ce31f657878c12c", x"afb165b2c356c5ab");
            when 14283740 => data <= (x"0f4705607e721fa4", x"9e683d419f1edaa2", x"86f9ff06256610be", x"387f5115d270eb2c", x"05d11d8b83790133", x"0dded59355a0e933", x"5f82260e82bf5f20", x"648610ac0aed3bf6");
            when 13329080 => data <= (x"89dab3b915cce0b5", x"39ca90657a98c7aa", x"1917810b0f24c3ea", x"b8b58cf6dee0dd4d", x"55cee03b9df4e81c", x"bfd089cf30dbb7d2", x"7739bf2c2081584b", x"11f7963dabf2ceba");
            when 27221327 => data <= (x"5f5ac663c277c2bb", x"cf25d823d169c0be", x"3bdaa156d557b822", x"1eb0684c6ba6ba6e", x"e3f16e8363451fc6", x"4d86cb1c7e731405", x"48ca4f49bca16313", x"80964893d39b85cf");
            when 30614734 => data <= (x"2f704befa7806b3a", x"f811a2f956e12d0f", x"8ed7eacb5d8cef0d", x"cc70b07fa2028855", x"54591090848b633c", x"78c1e1225d803e72", x"c4251bd2ae0e2835", x"f64a62568899f30e");
            when 22055759 => data <= (x"424f63b704e9d3c7", x"8a192be17e3a27a0", x"02ae781c0348b545", x"1caa7b623ef22a4f", x"b8a365bb7bdc9e8e", x"f14c7bd488d11bec", x"03a4ff92ba983f6e", x"decc238277b16cb4");
            when 9814704 => data <= (x"587b7a9ad7759123", x"6f1bb4719b431a4f", x"39872651671bf317", x"27492dde7ca2f285", x"3246c3fbb04d4d85", x"76bea63c709e5778", x"564f30e191c96c15", x"3fcb94f555d8deaa");
            when 28822665 => data <= (x"29d44571e5d2e849", x"7a98e06c165255fd", x"70e73a73a8b9dc09", x"b1d1d50f870447dd", x"e4a1a15afc8074cc", x"442818545ef475d9", x"45a27ae10a51171a", x"a231cf702d759212");
            when 14701149 => data <= (x"a8bf9ae12ecd5eef", x"66ec7913ffd0ff1e", x"23c7f4877ce86ea7", x"590bceaffdf36436", x"3b21fefb47577c60", x"7e366d13943c1281", x"1369ab83c64ee69d", x"83e7c49779180b62");
            when 24517117 => data <= (x"6e80e5d2dbaaf123", x"25bd06e8968bc0b3", x"9a5935a1eb393b1c", x"e99b12e806f192c7", x"608a2618c92249da", x"072a5467c3cda88f", x"7a9e987398fcf88b", x"1965a23d9f8f17c9");
            when 28974606 => data <= (x"105cc456d9b23dbb", x"1f5a4268eec95732", x"18574c08cb8f2b2b", x"6f0d9f60fbd8ae7c", x"1020a209d96cff00", x"e96fe83d21105c46", x"1a380bc3158fcc1d", x"40a0c2ece7bfb7ec");
            when 29409893 => data <= (x"410d4754f428ba26", x"68915899f0fdfe35", x"2adabb5c586b437f", x"957d5d6c3f34ec73", x"22190b98410b7e2f", x"6e70c9284401f2d6", x"1eadf50d99580250", x"c3246242c048cd95");
            when 14667915 => data <= (x"fbc81ba96e632ef8", x"96135531c1c8febf", x"dd55b19dbbce148d", x"c29c0407f39d7259", x"35723de0d660cbee", x"32392c2e1db83993", x"66f7490f387811c1", x"bd9d45c2792611b1");
            when 8625470 => data <= (x"7267caff86680078", x"36c87131208cad57", x"fa8c9395ae64ec32", x"997c80ab0f5f0969", x"d665d28f1d19c132", x"c2df9982d6168bce", x"5cefd18c473b4183", x"73872b5160724dd2");
            when 24190904 => data <= (x"bbfd0957d4ced8e2", x"cf77c6a0b31cd3d9", x"b4ed180f6b797378", x"10044dada46d5612", x"a4a6bbc698c25cf5", x"8db58bd5dd1c3ef1", x"94911c5048ddec68", x"6cd9c764d1fda3de");
            when 28616605 => data <= (x"8d3aad46c31ae6a5", x"ef1422a5010c3e30", x"f60b489cec11f7b9", x"70e9999b0079febf", x"30dcb18e059e4263", x"fcba545167d07189", x"cc7c9453fd06c853", x"60da36a7b042a2b2");
            when 20258687 => data <= (x"3a0bcaf68b039576", x"8abac25edbed68b5", x"17107b88c3b5dfa8", x"3b1b904513eccc1b", x"0df80ec0a4f3c546", x"068e3891a0fc746f", x"f66308c4f446a3db", x"ead86441b508d003");
            when 23431921 => data <= (x"c9ec4b3fc7e8c494", x"71ff655d67d20e6d", x"eb92ba8ba9877b40", x"147b7efff6e4752e", x"946c3291fb47711c", x"44c444c59ff9aced", x"7f6831141c14ac21", x"6f4e870c803d9acc");
            when 13401658 => data <= (x"09626a0b40608939", x"f5057c8c767437ed", x"b6f3967524d3aacc", x"f98f29e02956c993", x"3efc1513d3845ebb", x"f0a453a6fd49c687", x"a35419560979df14", x"d5b8250c4df5f20d");
            when 12656704 => data <= (x"69963e48c5433e4c", x"6b42a22d60f9c71c", x"80cfc70355044435", x"1f09863407fe2d9f", x"1f5ab8b700d15e62", x"ab91874cf24bed76", x"78733d6f520ec1a2", x"83639d5c85f65654");
            when 28566264 => data <= (x"453cbf9633dd8c10", x"c027be69f260349a", x"caa79c0beeb49720", x"d1141c17a5b76286", x"eff3101a1d7b31b8", x"917068b15b10cd90", x"066bfd32f83c4c53", x"2bf0df7ebfa5f719");
            when 32434068 => data <= (x"04ac73ea75284b9a", x"5a3a3f80c16cfbe4", x"f5230fd4f2d876b9", x"516bd436adbb0094", x"606a1cf4b5332d8c", x"3e0c2c98a241415b", x"f1167dcaa1185686", x"bc052c6198da7873");
            when 17676889 => data <= (x"fdcaaca1b1f3e8b3", x"95f86eb1ce0c13c0", x"129d8f8dcac35935", x"14094aab3c3cb08b", x"99df0ddd5c02d8e6", x"9de14c6b9d82a4c5", x"a8c74ad4fbc822d6", x"3f1da15ffd6c8865");
            when 664557 => data <= (x"ecf28fa038731ac2", x"3e0bf9cf56f0c9f8", x"636af1dbb21a8729", x"cbf071e4a7070970", x"4c035d76fb43d6b2", x"283df785733f31fc", x"2ba8edb2c41c928a", x"b791f98a6780fbc9");
            when 29066907 => data <= (x"3265f1d300a6250d", x"5da9ed15caa005c5", x"c985bcc22ac25eae", x"9d7804b9e18266d7", x"7a441961cd222c2d", x"249887a3823182e4", x"862ccd27fe076b43", x"745fd9f9c79f67d8");
            when 16798089 => data <= (x"590b903d8a768ded", x"56a6ba5177764bd6", x"183ccfa2c9625f40", x"95dcc7b9697613ea", x"c86993c8bcaf301f", x"1fe59542f56b614d", x"5e4a82d11816fe5a", x"595e1ed21693bfb1");
            when 2748437 => data <= (x"2e65869bf7105a5d", x"63714cdfa6f80618", x"f9edbce9716d822b", x"ac5c60747e26311e", x"5c80064cc09908f1", x"2b7c782413e68150", x"0076d7becb4563a5", x"a462a11b408bb27d");
            when 23538629 => data <= (x"181f2160451642cf", x"30b32a7a625f5fb1", x"4172d887fcf3b3a6", x"39bb59fbd84da6fc", x"d076c41c10b6d704", x"53d36343f455de0e", x"bd0c0882b47838a9", x"f8fe7d86863ab615");
            when 32462037 => data <= (x"369773a3f32374d8", x"55343265d521b61e", x"b44a3481d70d7a28", x"36cfed2f405dadc4", x"87f7b083f93f7ed2", x"0b5f65b67a871f89", x"da6c9e49c7f2c6bd", x"4d01221f65bfb950");
            when 5922848 => data <= (x"f9009bf8dfedbd63", x"d5ff41fc5db36df5", x"a3eccb7219f410ff", x"7c542706b7b0f398", x"05d64768bd14eb4d", x"7d8503a8a488035e", x"4a4ee527f715a605", x"d0328a0a310d9448");
            when 17768448 => data <= (x"8f1ecb61a5273ca7", x"f09ab1530ef664e4", x"b83dd742713efa59", x"05015c392a4f8d72", x"010149555e61e9ee", x"836be54c67782a01", x"ac2283ca942da04c", x"9bafa88f445a5da3");
            when 11379565 => data <= (x"f20506b744f28d74", x"0c0ce0850f4130ca", x"390810ced28dfc56", x"421611ad08435597", x"9adaf466d2ec4bb5", x"86065ca97d1a1fe3", x"c96f9c046b0f103f", x"f982cbb0c36104e1");
            when 5831795 => data <= (x"90d9b2608b54adde", x"7d476e3af26b5a22", x"da017ca7c63b45c2", x"17824ef3fa522cf6", x"95826b372b611931", x"a80bc296a8f948b4", x"bc1508e64283f1c3", x"493015eb9d25d8e0");
            when 31206511 => data <= (x"c488293ecf3ef9ee", x"806e841a9b2cccb4", x"e49fe2656c13fcfb", x"9a7725fc4f98e48a", x"e8f45c1bcd08ccf1", x"9b15caf69ca4fedc", x"4d46dc41887a27c5", x"596a6acd00536396");
            when 30144860 => data <= (x"906b4e11b02b908c", x"401ed9a295e5f346", x"51c8f844af21722d", x"640a073d11967f2e", x"fe3c96bb065e572c", x"eaf59150ffc35a48", x"d3bda465d40aaed1", x"54919f058115d3f4");
            when 5902065 => data <= (x"2106ea1c134f8e7a", x"ef21797fc1aed0c9", x"5afb8881426ff861", x"b47bbb32f2a170df", x"122ccb8766d4944e", x"45000336d1dbb1d2", x"a125d2cf3745e96e", x"7e9e7b14f7839027");
            when 28562892 => data <= (x"a0767f751fb1b4a4", x"ca1c002f1c3ddf18", x"fe1307e67988a113", x"2d580c5f967ba632", x"ebd6598545b5060d", x"9bf9a5a1ce83c11f", x"e5170885f94d7e6e", x"8e8bbed1126ad6ee");
            when 17966948 => data <= (x"3a192f0cc2cb64fb", x"cd001c5e7e4d9983", x"9806da41c9141b4c", x"19198578331ff3e0", x"3ef17fd1d4ed17fd", x"b5a76baaaa5a5f3f", x"a56c7ff57e4d48cf", x"14ca795aca3deb0e");
            when 25053327 => data <= (x"16c9197e72032302", x"52f9f2b32de538a6", x"dccc7ea79ff61c58", x"96b0ff674cdef468", x"99aad39c88d879e5", x"b1772b785587d0fc", x"4395983bbddbb5b1", x"0bd2cd51ba915f87");
            when 30801569 => data <= (x"f33313d80cfea7d8", x"2ce0c821b75c3b35", x"258f2bea97972c73", x"299ffa360d1bf367", x"12a2e790a6d049fa", x"a8e1b3f219eff41c", x"159fc3cb1cf3b671", x"2796d23ff239603f");
            when 12144417 => data <= (x"a484b3fd023baed0", x"21ff653555f27f4f", x"221db7a21253b748", x"d150188710401def", x"aa6860a446950ce9", x"4fb4382659c3364b", x"38ebed7d9085cb8f", x"9141f05c34e4274a");
            when 28756620 => data <= (x"fd7bdae74d821359", x"7f8e7c7d2bacf80c", x"c8a956cc708e1680", x"2dd2ccedee4640f7", x"c8e337f12da63689", x"c136629f167a217c", x"abacec0b71efc9d6", x"98e298ce960a5773");
            when 20099276 => data <= (x"4fe88fbcfae6d3ce", x"25d0016f7426599e", x"272627bcf9cda0f0", x"691fb746fa1ac6d4", x"15288041734e605d", x"1eb491d79905cd30", x"540baae94184b63e", x"a4343472d66ea96f");
            when 15274231 => data <= (x"5718bc208e1d1239", x"8136696a462f768c", x"0bd538259299dfc6", x"63eadfe5c6f64994", x"e2cb0fe471b80f20", x"83745fe3415db1b3", x"b941066177e844ca", x"3753fcbca8a73ae5");
            when 30483181 => data <= (x"3d7d3c6bd11c426c", x"4d222fb5d26cff6b", x"9480a59df5e5a6b9", x"9b260a088a0618df", x"ee31e40a6d1dd89e", x"be5512e3e0cd72ee", x"efb26e55ff03e142", x"f0be2c18b7ae8c85");
            when 24306132 => data <= (x"42b38db45f1ceda2", x"089bcfcb9cb37763", x"d75b3b3196cf5bda", x"e392a503ebb66c7a", x"b668f4d95f7c2529", x"a3d46a24affca8ce", x"b027e399b2284f15", x"e77053fc439030f9");
            when 18634532 => data <= (x"2f94933dd778bfd2", x"38bf9142b9f967d0", x"053926b86bf457fa", x"3566f8faca86b547", x"7ae453b9b949cb75", x"00995827eb0f2d5c", x"71a6291bea903dd5", x"baa4175879421833");
            when 9129634 => data <= (x"25bb0acb8c91378d", x"a5655476d52e8ead", x"cd0b76eda237b777", x"cc2ba7799c913762", x"09c75f19799930d1", x"84b80ddbfa7f83a7", x"3444eac2163b5da4", x"d42310153d5d6991");
            when 30402743 => data <= (x"18bc996e01b9e03b", x"ba917383fc5ef289", x"750f9de382b4d865", x"9690198b9b00515c", x"a15c4c95a5718d53", x"40975621fa86aa0f", x"3adca0ab94bf79ef", x"7acf604de8f4bfb4");
            when 18696974 => data <= (x"d19a3e4328de9d68", x"8a8da06531424f71", x"ad075b631231e3ad", x"eefb49ad2c0deaa1", x"4c4a7877e12f0b59", x"ea93ab8c5f3ba2df", x"0884d08d0aa854ac", x"c4546923e7b600d8");
            when 18487354 => data <= (x"2f06dc62484130c4", x"65d8a9afe5b86495", x"ca940dc60e62e387", x"0b3cecd21eab04cf", x"2a1f0429c3ee7e36", x"607e0b40330c22fe", x"870302d1263ee781", x"59d51b7432b7452f");
            when 31354629 => data <= (x"4241a7c37ac012ec", x"119162edc957afc0", x"c8b207bd44066be2", x"6868c874e916a87e", x"749dee164f3db4a4", x"840d8cc64d3e7c31", x"df45957ed8d53891", x"9a884a0313883f18");
            when 21889279 => data <= (x"4c7ede6ef98ea823", x"2e221b3925b55029", x"788578598a208743", x"e0a685150cbc77f8", x"39b5b9d5e39d4f71", x"a166fae1eb6b258e", x"61c7e8f721cf26b2", x"dc063b32ada300b9");
            when 32938915 => data <= (x"97a27ede0c2bda28", x"81e039ebceef1267", x"750b5a52047c1081", x"f0860a5e9e3c0bda", x"20b5948e65dd44cf", x"357259cbff1f1f68", x"edb25ce501c50ac8", x"5bdd35f34d140f41");
            when 24557649 => data <= (x"5b6cf84bbd03bad9", x"ee6566f37cb2d6ac", x"033a1cffa216f4a9", x"355c42d61427ef51", x"95faf473e14208e1", x"5cc201f69a864b36", x"44daef547e7b36b4", x"f0985bbd5b204e5e");
            when 23948118 => data <= (x"440614eb894a5279", x"3a5c678be40f08c2", x"1d4fcc96271e32d6", x"7285b6c2a51c0f03", x"18bf01812aafdb40", x"66115a2c5312c016", x"4a92828f48b14acd", x"bec834706b28a040");
            when 23295526 => data <= (x"8141b02540537259", x"8b3900ef4b8dad76", x"2ddb114264a714fd", x"d27e4f43433f9a67", x"e8da4e4585ee1819", x"9e379e458c44431e", x"bb53a7e1e0c6b58d", x"d5b128236ed11393");
            when 28939021 => data <= (x"1d7deca442b3e070", x"b2422eaaf98f6390", x"d908e484b39eca08", x"4c8049ee8e150ef0", x"1704e27adc1a1054", x"ffcbd39fb888de08", x"ba9886811a820211", x"4b110beff7e9ff5f");
            when 10461352 => data <= (x"feafcbede69c6a70", x"6eb00edf942e69fc", x"e526fcd844538d6e", x"aea02b58902b5aea", x"5ae2d36d92c935ba", x"c9f6c3926cd13046", x"5c2c4443a9ed9edd", x"d815c170a699ebe9");
            when 12843302 => data <= (x"97b77f35e7a1b3fa", x"74ecce1a88a38cf6", x"01cada64a37f9b3d", x"b4d78b8070b38626", x"9598ef27686a3409", x"ff51a0ddf4a652f0", x"f19ffbad23e2dc8a", x"f09a384cda23a974");
            when 19016768 => data <= (x"8912661877b89e42", x"b1d46e6a59744242", x"5b056cfd24028e88", x"a76931377df33796", x"0e44c4516061cf1b", x"380694933b9822d1", x"c57f118946b59a4d", x"fa838ea8ef5083aa");
            when 30996818 => data <= (x"94b20bb22a95a27a", x"a448071fed35c5b5", x"ebbe4436eb1301a9", x"34bf08f0b6fa6c4e", x"316849e2e7d24c9f", x"0ed2a52b31f702a3", x"72bb733b6f2c2480", x"a4f3e2d2542466fa");
            when 29642788 => data <= (x"eca08b098efd4eff", x"acde6040c2932651", x"cb82521f67bc83d9", x"6d65c896f6947a65", x"6a650429922a99a7", x"995c83a3d32e75e9", x"9fb79fc1435c994c", x"419369760955ac0c");
            when 6258503 => data <= (x"a18d84fb595c0175", x"52b2e03afd411389", x"6804a4245eb02067", x"40fc839c15d2775f", x"20217e2153e89185", x"d30c9b97aadc40e8", x"5957cb5777f8f425", x"39b20fe855657907");
            when 20885279 => data <= (x"473b1859665e2358", x"63e83f21a054add3", x"23a7ab4c4721a649", x"543e8f61f1ab0888", x"55a5e80e8fcfd974", x"cb45f0d755c618cf", x"74ba729eafd975a9", x"2e7c5a7f9aabcc8d");
            when 2211361 => data <= (x"9b87265f51dbe2c0", x"2a950cfdbd2b8781", x"dcab6de0fa8146d1", x"18d01ee99a92ba43", x"42fb1a4bb3e0592a", x"d9b24030bf162558", x"226dd3e74a2b7e38", x"0e530965bbdbbdaf");
            when 20793619 => data <= (x"6eea9bc0eee73d0b", x"5d5726a636cba61a", x"b5c2795531a0972f", x"93a33631befa6da3", x"283fc941577637ba", x"c6727ed64af9b1e7", x"e382de243f906140", x"1a1e586bae9b600d");
            when 27491751 => data <= (x"3e5f7f2e1a6b4db7", x"6bd92e4ceffee840", x"2293ec1bd716acc1", x"be48fb3047a7ecdf", x"3cbbc710161af214", x"e6e673e32e4e5cab", x"f6106d84cbf47834", x"704706554a10960c");
            when 7771385 => data <= (x"af12a60033e214bd", x"8f6075b10d0e0d17", x"af3426e955030b78", x"81cb40c42ba0f1e1", x"f8988dabfacb40f1", x"47d6db7335955e18", x"ddd849715c6039f8", x"760b0974e0f25562");
            when 10083892 => data <= (x"f6fad2b77723ebd6", x"842b57a10235d16c", x"49a8d2b0b8b8ef82", x"1b612f7d0a834624", x"3d698c8eaee5129d", x"64b9cf61b72a0f3a", x"e4fc9603ffaff97d", x"fa9599d90b297eb1");
            when 25313668 => data <= (x"b61f235ad9551592", x"74154eb3a57f000c", x"0a38e2e2ac7b637f", x"a69a80ac7c9a13c6", x"76595d2d4d447f8b", x"847e89e4c9846fbf", x"4b3307c8e157c887", x"32f09623b8ae7752");
            when 3275920 => data <= (x"49aa9b3565b22aa8", x"88da284dd051a61a", x"6d7397c6ed5f16d7", x"94bd288a6a59e73d", x"98f750ffef9e4944", x"997db244295eba0f", x"4aa79093f8e3f127", x"aeabddbffbfd921e");
            when 17025713 => data <= (x"e0137d689a35df40", x"1ff58535eb61d878", x"9240fa65ac0cfa91", x"4b825d9f58197a19", x"a4caa04361681b3b", x"7691367384c91979", x"b41a433bcfd68769", x"3001e4b24ed33bcd");
            when 21922934 => data <= (x"347f3096fd5baee5", x"6088708495d29a71", x"98a2855ab7bffd28", x"14e4fe1e06f2d293", x"0f27efad7c86a9ef", x"8da84a3fcf328d09", x"7a5ac3ae61c5abdb", x"385e616ce8ae46a0");
            when 30403195 => data <= (x"7e249f910337ba9b", x"47804bb9c5a191e0", x"94acd81c22baf029", x"4c6285b8c546eff8", x"88d8ffbe12052776", x"b4c620cd05c6c522", x"0e0f2f0ff9309a0d", x"309c0a0b72a0dc70");
            when 31005253 => data <= (x"4c75214c77ecad35", x"c2447f5196869128", x"97dd87b47cb079d7", x"262490a26e017484", x"8e55a92e76f5f7e2", x"f31202f111766aa6", x"89b43a72c90b2a9b", x"3972f27af8bed7b5");
            when 4049819 => data <= (x"e2bad238eb4d293b", x"17ad93f1c8f55e09", x"8a7afdb9a4da6fae", x"c61b5b3a7333fa00", x"5990dc29835229c4", x"b7621452bddfffc1", x"ca1c447ac44f5bc9", x"a8419a2a8ac025c7");
            when 18256143 => data <= (x"625a3453740cc9c5", x"918b3ae99793fb7e", x"2652f095018cea86", x"866118c1bc6fd668", x"2a0e07a163fc2e65", x"b52d91aa30a748af", x"c18af97c0486a2f4", x"47ec1ec22b93e69d");
            when 8444228 => data <= (x"43859058d0442d28", x"cf0749b50cd7d5df", x"57507ea91435c9db", x"b61028ab18ae196b", x"2830278fedbdafa2", x"04a0f38de411c406", x"c1c45d9fe1509fd0", x"0fc8731e93784290");
            when 27308643 => data <= (x"868e3f6b2350a01e", x"1cc373ef0b316b68", x"0400399714338848", x"33039b002fe6deb6", x"00d86ea2064a1d64", x"7ebb542678640287", x"34713244e17860c6", x"e789b859c55c482d");
            when 16616948 => data <= (x"11c593548eaa76f8", x"02dd8a4269bbde91", x"1638bb0e659d4526", x"ce105b65df63813f", x"991ff7bf4a516b1c", x"3285e968245b70fd", x"341f8fb01318cd29", x"c46d53f2ad83a5d6");
            when 27668262 => data <= (x"2a773c6b5375739d", x"ac03de5f1d06a0d5", x"201a0bacaefc972d", x"58cae28bc450ff17", x"9d2f6c2f75048d9b", x"5bfa99b4537b2f95", x"28a678e670919acf", x"1793b80fc639d790");
            when 4483627 => data <= (x"e73b70b80774f500", x"e678355f9483f173", x"0677c076d91503ec", x"559b121b7d3d1f81", x"4275359394320a16", x"b0efe132305b9e16", x"0501b253b067eac6", x"0c5edc7f051d7618");
            when 9512219 => data <= (x"9ef33a78d6f0444e", x"befdb2d6ceebca3d", x"9361dffca2e5458f", x"45c223be0c005d94", x"36346263a3f6ee5c", x"62aea26894ed6d13", x"76fc7235f8ce7662", x"becb22f31e5b0d18");
            when 20401299 => data <= (x"94ba079567b8784f", x"a916b4828603e719", x"1a1c9c273ab68181", x"b6637c37e665b74b", x"5c7d75740aede4a6", x"9c80a580f615cf83", x"d3fbd9089e044e53", x"227b4785cf90902f");
            when 23723493 => data <= (x"03c16293c59d066a", x"9b195cfbc5469b5a", x"4178f3381ea4b700", x"3cfbb15edda939ef", x"bcd7c17cc2a74599", x"39b11db9d9f49819", x"d49d4e10030c067a", x"ddca0db652130b25");
            when 22345039 => data <= (x"37433bd65897712a", x"a4a4a63b84c82104", x"0c41bf82921f04d2", x"e7a1727ea1a9f098", x"707bd3ac44707309", x"7a33b1ac47241df9", x"b021858e99f7fe59", x"59b64221247e2ec2");
            when 22890961 => data <= (x"a0a96da45f694b41", x"e017023546b6ef6d", x"e8e744150184cd3e", x"20c7814f280a4f61", x"9f350ef55f3b3908", x"0e26d01acaa53399", x"9c843d00d615de39", x"091771b40358ae37");
            when 11635034 => data <= (x"c96745387887b74a", x"82f1fa8cbe62973e", x"a52df839de69cccc", x"166a0dbf854d5ded", x"d6578c87f92534fb", x"baa308d38be1ecd2", x"c1eafd621380c893", x"cc861ec9f778746d");
            when 9503222 => data <= (x"9120c8cb186575fb", x"518e68e484335529", x"c400306c648686ee", x"010333b5e6ae575e", x"9025d7d153e4d2a4", x"02dc7a9742556e11", x"d5915a1abb759440", x"b29822ea85912c5f");
            when 26481973 => data <= (x"94071307f8d9e62c", x"81515be6b6c95cf5", x"3b9250fc94a6feaa", x"3504d18c762fc1a9", x"3d0f88761c284cb0", x"9647ef4b07c2e3eb", x"b638ea164281c226", x"9cf643cbe924d4a6");
            when 12777006 => data <= (x"1c3ea88e4ca9ebe7", x"a41ad6e0dddf556e", x"7af417e1fd076246", x"a1f5f7bb638ea928", x"ee6d0c9df25e3299", x"6308ff8d6f2cd5b7", x"7b03c4303121732f", x"da02bcef0f7ade0c");
            when 16445100 => data <= (x"4066481e019a0714", x"81feb9c8754b789f", x"bde59305c94a1498", x"910d40d0eabdc395", x"5a4ae08921bbd36d", x"8332eefaee51f2e0", x"ecb0b4c98ef743dc", x"349da9d929e7f64c");
            when 19444025 => data <= (x"6031f0b752f17e9d", x"640827c3ed88d8b1", x"fed25f93a6ffac89", x"b7844203e401be38", x"01712490d18a8c00", x"6d94615abc90fd5f", x"dc5582a3b0113cdd", x"548425d11af9f2ef");
            when 14962443 => data <= (x"b7f744008dd291ab", x"7e698bf5502eee22", x"7bf427e41e0171e9", x"40b8f99fa1fe4092", x"7f0b7c19ce54468a", x"f4130fbbed7766bb", x"dd2a923dd69b9512", x"201e140d620d4934");
            when 3887370 => data <= (x"bdc3f28d026bd652", x"a722d6cce0465da0", x"373ff01f1bf2ab5a", x"8b42445366328e42", x"ecbb5f6c81109c0f", x"d5a605d85690c61a", x"cbbc656d6a1da5a1", x"092edc6ee5a22957");
            when 33554653 => data <= (x"1a85efa9bfde9f6b", x"56e9d8217a17b665", x"ca3d2ba9e2246f71", x"8fa829b0c7d227e9", x"5ac5a820a93ad5a4", x"06a0cf5d1ca6f9cc", x"7878b2be5ae4e0cf", x"52880ccec8c93b3b");
            when 3367271 => data <= (x"2901b02a87629046", x"40a2fdccbd2e00b3", x"f7c657eab69784e2", x"0daf45ce3165e9b0", x"b70d1db6afb9b43f", x"a4b6152b786933d2", x"8643e08216feafc6", x"2dd29771859c1832");
            when 14651676 => data <= (x"7cfff02a2b705b7e", x"f0fa9570cc0ebe01", x"68821b535cfefa6c", x"ffcd45ec3e1e60d6", x"986494254ebd4074", x"24fe865905ab113f", x"f238ac3948b5dd86", x"f6eb73ed70a739f5");
            when 900330 => data <= (x"3f15cbb2f7840f17", x"0155a75db59f71a5", x"3486966e902194ec", x"18cb042034624bde", x"44a232fb2a80a3e2", x"4bd07f7bd74d5eac", x"c25e01e6cb2d5e10", x"0f1ad89ef7c42efe");
            when 17597947 => data <= (x"6886a31cc254457d", x"9c02b28cf96066e2", x"1858a0133f526af6", x"b1dc9ea640ecc52e", x"5aff14bdb6226aa9", x"e4ed372b3fd56501", x"64f245c1507795f5", x"bd41aa1fd637ceed");
            when 18650940 => data <= (x"a4f0d2ad1e088c02", x"1fe651f1e7e0c735", x"e3e6fd5ce8b57af5", x"486c8171ec353cdf", x"8087467ce706828e", x"82f1670d3b2fca94", x"7a9487b89b10caa2", x"5ecb8a6a8fd8108a");
            when 7420716 => data <= (x"8113233bb4b911fd", x"5cdecd6702ae7575", x"d3ac389fe0d9a316", x"cb6d8a6b48dc61d5", x"97de879e0fdadd8f", x"fa704a33be7b4004", x"cb85bbdc95bf81f3", x"6e60f32a2bf0c418");
            when 31586292 => data <= (x"65e0b7b215d5f179", x"860db0af1ac12b66", x"9450b6dc7f00d9b3", x"391e0df1bc8b0e22", x"bb818875dcc9f18f", x"018c784e0bb3cfaa", x"f870bd035e025835", x"cb334a3d487dab3f");
            when 26379538 => data <= (x"550ccf3f059317bb", x"46e9e00e27c7c909", x"6fdbe8d456ff2a7a", x"6247374e0ad0ad6c", x"6bd89f5a55688d41", x"3c7d3649e6297125", x"5631b0ebf98db45d", x"abac63e3f2842b0c");
            when 16291061 => data <= (x"1c24ad37cd3577df", x"e30347502fdead47", x"e5581ee640cec18d", x"aa254e8c03846955", x"0cb733f91de9904c", x"9a7649be9f0a9875", x"3527538d8a0db22b", x"d1b54d55d80892b4");
            when 31628657 => data <= (x"07e27304dfa6a764", x"d0292be7994bc237", x"30a0e9da1a087110", x"b0404729b31a83e1", x"dc7948ef12a443c7", x"16281db191c81f66", x"de24e7ce2dd805d1", x"29bd39168c8ba526");
            when 33488035 => data <= (x"878ed1a912e97d1f", x"b4947f1f7c396332", x"c88ec33034853173", x"56cfd5cbc7c9063e", x"fa2439ea4d065f3c", x"1dd38d790bf7101b", x"dc199729032715c0", x"7840b09889a5c227");
            when 28899434 => data <= (x"cb1f9a1852d928bc", x"af3938bf73d5c943", x"3fe9c8f5a228d377", x"d3a90b9cf2a45f4e", x"9bc4265278940c9e", x"ff02538bdd729790", x"548fba12a263b186", x"fe9f6d469316bc7a");
            when 17035634 => data <= (x"ab71ebb1765caa38", x"c2a7f60267928fdd", x"aab75ffd391ea7d3", x"c0adb6d36c1b59d3", x"79245acb29faf311", x"4f198b97f07bb5af", x"aab8dcc3afd59286", x"428b78229b9dcaff");
            when 4379203 => data <= (x"d455b63bc63611d4", x"b4a81c7fff0dfa6f", x"25b2301f3de205ea", x"419e7b341347cc9f", x"bc90344eb47bb2f8", x"1d920c9caffec725", x"08c5895d67a0a44e", x"4eb50a847ee014d7");
            when 32133830 => data <= (x"de261c17e1ceddd1", x"a83f065f55dd7af3", x"c656590869d9ae91", x"6ad7cf879fdf3473", x"3cdff58ef12dbb2f", x"77ee45ea743e4bee", x"27fd3afee98e9201", x"6ce35b14de6caa19");
            when 12348450 => data <= (x"157bf9af3eb80c9d", x"579448a535d689c3", x"aad04ed357524cfd", x"ec83e7fdeb3864a0", x"f0aca2bed79e0d4e", x"fbcaad410d2a10a8", x"b764d46a4052aa59", x"d1773c6ed2f536b8");
            when 10548736 => data <= (x"8a9892fd96492ddf", x"f61b9549643bc1ea", x"cf9a2b1ff15a39e6", x"ad312d69dde23223", x"5261e39f230aff72", x"73ff33e366275ba0", x"190a18e5949eae78", x"50a6e946166b5ace");
            when 25509811 => data <= (x"56a0f84e66fadba3", x"b9ce6212f9c5184c", x"6f0584f81caaa01f", x"ddd5f9cb8f52a08d", x"25211e27c3efa837", x"0f769a01cf8e5012", x"955529bb514aa8b4", x"bb4442ef535a8725");
            when 19855206 => data <= (x"40d01b90730e7382", x"20b2db7d17f8fb89", x"a48059d99a696934", x"a5935c7fd6eacfc1", x"b86415d80c67fcfa", x"351373190ea61f58", x"70f2682197a1ac0b", x"231b4fe9216ef07d");
            when 33566628 => data <= (x"0be8a7fdea26d974", x"c6eb9e347f9fb72d", x"7e5657ee0cd96d63", x"3278faef319aa89b", x"286b29e6fbdb5fe6", x"5eeb5d36de20e2ad", x"ea62ecd4f095a1d2", x"c5c44f0a46ae9305");
            when 8811046 => data <= (x"5fc3ada5fa25a70c", x"bf2e0788995b8c89", x"da01814cda34d124", x"115d366e18ed8f47", x"344812ab5046e257", x"de13520250288fd4", x"114287688da87718", x"62a0546885125b2b");
            when 7682654 => data <= (x"4a18a3b0194d1076", x"b574666af7ce0ace", x"92dd8cc1960fa4b3", x"278dac9c725ba9f6", x"00138673426db833", x"0e19fb58683b3393", x"5b71fd6482990a85", x"f5b8911411798453");
            when 25431935 => data <= (x"b2f27fc848185223", x"759fe2d8d78c128f", x"e9dbf87c63ad8f4e", x"8d85dc4fd4b4c3f3", x"03965e9c894ba271", x"d15bf0bd3fa52326", x"43f4fd255dc5eec6", x"8c07d08c400c67f1");
            when 30896130 => data <= (x"eb99ca95c7e741a1", x"4010591809634a3c", x"3072f5c7187c93ff", x"a7476c7956654167", x"837c3f59d1dcd844", x"7c91c2990e6f0507", x"32307fd1f32e9d79", x"b701cc746a120d5d");
            when 22853428 => data <= (x"5b4c01806207d921", x"02c9ba1e51e8a434", x"6b92c671240f2582", x"9d902918cb70857f", x"acaec2c8c410ed54", x"91b044068817ab6f", x"986ad0523d703e51", x"19fd67bda16c37c0");
            when 15772396 => data <= (x"29bc6a753381b95b", x"e9fca5b5e89a8934", x"7c2d20e4144f5de7", x"fad42f5da6057a5c", x"d9ef4fc4aefdb974", x"7c8feba23408bd6e", x"6f6b66df37656bb4", x"dd742b1580f812db");
            when 8562135 => data <= (x"ccdd5a0b8a72f956", x"e8c99361470cbe3b", x"dc259e0f6d676cc7", x"0d21e4b99cc7fac3", x"0c9766c2eb840376", x"55854b9def6b1e06", x"82663c1fb75bbfba", x"d353d433d8a8638e");
            when 28273117 => data <= (x"1b98d5e94864efaf", x"7065e640a913c255", x"35bc846fefa901c5", x"27b6fd7b9460da38", x"30d76e078824a3ca", x"dcef0160e4a19697", x"7c012fb2ad83f1d0", x"5fe80fe9b9741126");
            when 11255898 => data <= (x"8037e87d0db55f67", x"575b378d95d6d54f", x"24a0b80ab8a1430a", x"0c340d32abc3f98a", x"0057758ff9ad6cdf", x"8d1b0cfb9a90ed2c", x"3b3483e240a8830f", x"2c1dd7a686869b21");
            when 2593793 => data <= (x"0a619aa947429a5d", x"d913ffdd42a38d27", x"785041076e5f7b0b", x"dd11fb2c5c13f211", x"b06482ae223399da", x"2411385bce97ed7e", x"9a9c315823b1ea16", x"9427e3e88b2e26c3");
            when 13367577 => data <= (x"6462c2ea21ebbaef", x"5bce77a26d854f18", x"7baf7fc161cc8e05", x"140e6f29e09d6e2d", x"1a303352a5ddadc6", x"f75aab28ca6d939a", x"bd7e2ba57aa62eb0", x"7486bdcdde8f5bd3");
            when 31222109 => data <= (x"70fe807dbfcdfda4", x"b4cf1aa7c990e9eb", x"03270752e76379d0", x"c0f3b547ca30407b", x"e07f6c4489485b6a", x"21eabf4905359ad8", x"7608010db22f058f", x"c9f790c652da2be7");
            when 22534511 => data <= (x"6e7c503dbf5db73e", x"8c0ae105766ed050", x"52efc500c8522abd", x"efd854a6b269a95d", x"65a7882f20090624", x"577faeb2c71b0a3e", x"fae4ab0108b9147c", x"297a4c6f79a54f86");
            when 27812089 => data <= (x"6185c26919a8b4a1", x"e6af926073bce732", x"505cbe18385e0bfc", x"0cd023383b857f5b", x"11bfc9d6dbf7dbae", x"76a2730d4f162e6c", x"ac362ad3f7f1be0b", x"ef4057b1e9dbba36");
            when 30045332 => data <= (x"4629753fcd5ab101", x"5262261a3959adcb", x"74bfe4c761906f6d", x"e1081c4128893fbb", x"88151234fff781e5", x"941e5d4f32a335fc", x"c32d1b7db81a9d47", x"61bf76b1e7f8fe0b");
            when 32666018 => data <= (x"6f608dfd624c00d8", x"d8f8b56b6ac7c900", x"7ec01bb96fcbf359", x"aee5f8a1a70914c7", x"becdb37ea80db621", x"bd0de373dc49eb5e", x"33689c95bd4860b2", x"117388a0f72d8aa2");
            when 15381193 => data <= (x"b81a778348cdd207", x"55fcedfdb63eeb97", x"07039c1cba381a1c", x"9482835238e90d3b", x"499d142d9560d9a3", x"8996e3189e9015c3", x"97eada49cc2d72ee", x"b218959bbc871c3a");
            when 14660225 => data <= (x"d35c684df1a012c7", x"c047780c26a53de1", x"228ecac1e8735bb9", x"4a24bad2d1fa08e5", x"a4ce6b4f2804b498", x"b7e0c4256ac65c5b", x"c4a1f694c1cc2fea", x"7447d8db0148d924");
            when 9867605 => data <= (x"a6f2672f9bf21a10", x"f52ee3f941160088", x"2d660556e60ae514", x"9712236fcf493d6e", x"f0ce0d60a78e6d2f", x"5b3fb16f9a052638", x"d76e264402bb080f", x"64959453ab75b641");
            when 11130069 => data <= (x"b8e88a2e81060bed", x"4dae129d95533d89", x"78e177a5adf2e985", x"207b91acf040b94f", x"dbae693dfaa38afb", x"f2c7b63f0ffc6cc6", x"f2368d97cc16254b", x"3d4d7ad3848b5a73");
            when 19502016 => data <= (x"217229229642e6de", x"b5c30e72bc1df846", x"f803f16bc2ec8ef6", x"c7226674f3e9dffc", x"241d0ece5ce8255a", x"449d5b4e18f9f421", x"b7b520b0488f32ab", x"955351a9bcc49baf");
            when 6444770 => data <= (x"2c18bc282f37b778", x"999ec5ff6e47c602", x"07bb7fabf8e9897d", x"c445fcd8412b7726", x"9b41b6695488b83b", x"2d060e551d8aa495", x"06ace43399f6f2d3", x"3535053b077336d0");
            when 18755807 => data <= (x"6931105367f66c22", x"27b7927794d055d8", x"acd617217fb09e11", x"0159863ef67ac117", x"e2834acb9baa0884", x"ae784bb950df6ae8", x"29170995b686dd7f", x"072cce52c2bbac91");
            when 14480926 => data <= (x"24b8a5aa715ef28d", x"225522ddf7568892", x"c20d6c2eb6856b36", x"6cd8d673a52707b7", x"61406d0652b13667", x"6bff2ce5c667e2e1", x"4ab8017593829a4f", x"73c726414642a9ef");
            when 9786843 => data <= (x"ac562be4cfa9e627", x"a0e3feb02a6f162f", x"0f16912b50d2ceed", x"3078b0be97074da4", x"5f8eb32e5c34e2b2", x"2560c3f83aa47787", x"a8c5b2c22367a52a", x"9ba9ccbcd15b507e");
            when 13848926 => data <= (x"30d19a5ba1ca5dfc", x"c2d9bfb5c431ef12", x"0d4aea37f36d0175", x"ed249ad83b837393", x"402ce6ecfd81d869", x"7d48afb2ea6dd61c", x"0c584db076bd4555", x"7d4889366b704157");
            when 7848646 => data <= (x"f10a6285f52cba10", x"5f284786920beaed", x"fdb650ff6467ba45", x"5cb668d3bdbdb3ee", x"c8ff0d0a36854a5f", x"df5059224333bf0c", x"9e4cba2eed06c727", x"9e020912b463e754");
            when 21712365 => data <= (x"ae15cb0413ad27ba", x"f612f182db60eb68", x"547c0acf973ccc3b", x"e08c3f7a26501ed3", x"b919c98db634de3c", x"fde24b5e6df70ff7", x"a354e0417e254098", x"69426d41928c7e41");
            when 28356949 => data <= (x"e288df5f1b092d21", x"cbbe266b1beb5eca", x"1484e300a0aa0776", x"554cf8e98e2016be", x"8aca6c060764ff03", x"0d4e653aaa227612", x"53ffd0dc5de132df", x"c026f807b3f84d4b");
            when 32811852 => data <= (x"bbbebc60ef437553", x"2c4df87f7185896b", x"7db9cf31fb035c1b", x"2313803d1b8c7a9d", x"7fae868928e155f3", x"06b8b87c3386f2e8", x"ef0ab046399c26ca", x"06994be50f64548e");
            when 6015909 => data <= (x"296905cfdeb140e5", x"029931bb3311b4c3", x"1971afc4b80eb473", x"c8d31a58919f96e4", x"3ef3e4fe588134f7", x"6b3bb34582a6225f", x"51d1635fc0f34a7e", x"727cb6d323c29a1e");
            when 30904630 => data <= (x"8dfef61e72b4f03d", x"10ae38c31552becd", x"aba8cc1a3619d66d", x"ec10d76bd2d3c243", x"67ff685990788fb1", x"ad26ab105480e5ed", x"0e4c375f1ba8d27d", x"9a305fd1dbb397bc");
            when 7051889 => data <= (x"6711e3d1a28640ff", x"8afcd77176301e03", x"cec372e4e1c7a56c", x"85763bb9b947e9dd", x"c577d9bc732b0472", x"71889df4476b93ad", x"e835cc52a85279e1", x"9d714d6cc9bd5605");
            when 20627079 => data <= (x"429902435713108c", x"4d0d27edcc7728d4", x"13a34794d80ba418", x"af15cccb4cee784c", x"b0c086277ba70a6d", x"8d7709376531520f", x"e0a2d27dcc1e1b31", x"436521e576cc1b1c");
            when 31626863 => data <= (x"ff022e9116d1a293", x"2a2eaf735d873916", x"4953447bbbe82594", x"874dad5af0b3537d", x"8935221abb27cfda", x"d40eca3415f28cdb", x"a0ba025f540bd9a9", x"d58cbd306682531f");
            when 13397610 => data <= (x"109ab3fd0f3a3744", x"1cd9d4ccd65917a7", x"182d668d39363e19", x"d54b75340ef9231a", x"19fe3deae0ab12a9", x"0513c512e8ac99f0", x"0d4892ae87a0bd65", x"975628d7d367b19b");
            when 15789012 => data <= (x"eb5a11e544deabd5", x"dd9318a97471b6ff", x"8e5e260a752171b6", x"cf9035c3942d3920", x"38bc3852807a6807", x"e806c31cfd2655b1", x"1e54f5f8e9c88380", x"415c07da0f6299e9");
            when 5443245 => data <= (x"985ea425fea3159d", x"6b6fac410824bebe", x"71af534341c01dc1", x"7410b85e0f2db375", x"ae4c6d0a0f48eff5", x"a845442663fa717d", x"78bf12751af37056", x"28bb885f3f7a1f71");
            when 21947185 => data <= (x"19e0b3ed8bb687fe", x"59a485a57436443e", x"a369cf7e33fc7556", x"96eeb4a91be92714", x"32a36f22d7ee110b", x"3f6b999a72f246f5", x"b937cc76e56cc29e", x"eaf433b8eed31e0d");
            when 3116910 => data <= (x"ddb99f2762ce1c50", x"9eaa54f2cc0237ce", x"0deb3ad87ad13b12", x"ce8ebba3f9b86ac0", x"3d308ea8a400c22e", x"dc76c72b9b03d052", x"683de1a01f6a69bd", x"ed45116d814c164c");
            when 19635146 => data <= (x"d900ea1b2a2f1a3b", x"efd61b0a83c8c59e", x"ae65a1479e45cfc6", x"43948acb50515f0d", x"60b40dc56322c2ea", x"4aa83b5695e0c7ae", x"8e6c2a01effb1a47", x"e6d2122db0267e29");
            when 21688573 => data <= (x"6cb5bc90c9acc9cd", x"e4e1d883eff3fcb3", x"70a9fef434e052f6", x"3d9c72f9862e5f44", x"6a16e62431477f5c", x"a0fe31430e9f49e8", x"52b499f880da8861", x"bfae6d9e1c32609b");
            when 18915156 => data <= (x"425fdeb4f51ed9e2", x"b948ddc0a7fba679", x"5aa0f3ac3bb688f3", x"d577650a5787dcf1", x"a884643457bb47d3", x"6c159f2f49201457", x"58d74881e9ac7710", x"1148ded27f625351");
            when 15784148 => data <= (x"b9d88a1fd69bff2d", x"8aee597081285d12", x"0d0d3315df482795", x"95719734cb6a1c32", x"7406ed88466343e0", x"567e73987a2cce1e", x"dd73124fd84f2057", x"93a1dc7653aa5870");
            when 16455392 => data <= (x"3933a31f7023d3c3", x"6d155d0be067b503", x"1fc3dd1b9c989e5b", x"06bf478fd425f1ec", x"a90d6d7b6bad526b", x"7740545d606afabe", x"1fb1cfe23e6ab51d", x"a05439d6c0343eda");
            when 10570871 => data <= (x"2e60bcff1567849f", x"5b2ba01b4aafee29", x"5a23d610b12f4a4e", x"2b2df661bafbdb44", x"a6095ecfedf08ccf", x"417b0771490a845e", x"e3e9e5be03e5016d", x"f7a80c5eced91c43");
            when 33691045 => data <= (x"271fffe0e324fad7", x"f60309e016318a61", x"057b618472d886ca", x"d78ca7bdd1ab7815", x"e09b09e4d10f1e1e", x"86e253ad60b329de", x"6ed95f76f2bb8fb2", x"19bc6a9b95e69c6e");
            when 22226806 => data <= (x"7a796084a290d90b", x"d00e873333815e8d", x"3dbb7420c338787c", x"a448b84c859edb8e", x"042aed97638aab6d", x"bb4d192f7eeed63a", x"badec88689082f50", x"2c505f51092d6913");
            when 27902284 => data <= (x"3982ed1e93230bc4", x"1ae8dcac39c74fef", x"d0c2495dde3cae99", x"72bcb128798da546", x"d9050cb2eb370709", x"738ed79ef50c9703", x"a474bf091751a6d9", x"fdb11e50cd3f11aa");
            when 13311116 => data <= (x"c5362f6f5029f54c", x"606f63bf5d9d3a83", x"fdb5821792c9c81a", x"6d0ff7a25bebcf1f", x"f10a1772913faf13", x"99a57dd8c30ad42e", x"6bc2679db71444cc", x"578704507a4a6dbb");
            when 14185736 => data <= (x"076abf7561f9c54c", x"e6b5fbcb0b28a301", x"74b49c4077aad340", x"84bba6e7fde9bd40", x"c2f4af7ac7929079", x"39f6e532b29ece2a", x"bdd35fdbf32f2b7d", x"43030b49d09c6e67");
            when 5864373 => data <= (x"fc678f1538042702", x"7676601b06d9e7c3", x"c7aab36db717764b", x"991f5af6a82c5046", x"6c1393f7f42ab7e4", x"40250212e5da44d6", x"530b89f82eb8c75e", x"1dd7edc471473e84");
            when 4636591 => data <= (x"9fb1ddf192f952a4", x"b0c7be9b801150ba", x"6c89d4b67e5885b1", x"d782175c359bedf6", x"dd3a0fef0caaa6c3", x"4eef754e08971ade", x"50cc5372341fbfbe", x"9b86f61f8251bbf4");
            when 26152580 => data <= (x"0e5a7022020c8302", x"fc10f0b2b42d6773", x"23243531fa09b8b9", x"d72c39b917eafbdb", x"45b2bf1166b45324", x"b66aba94b16fdaa2", x"64d106c7c8c1e517", x"da2dfd6ebbe00d2c");
            when 21861878 => data <= (x"de4588b77b35aafb", x"39af1eec4d3d830f", x"822ca403ef3d918e", x"2073f2952ebe9d0b", x"c357503af054dbb6", x"390174c82fad0179", x"bfedeb1cd9ab5d6c", x"00ef6fc0c5816a8d");
            when 12811129 => data <= (x"e23895ff959d789e", x"d5e03255d284c96f", x"394eddd9aba8ae85", x"6123a733a3172986", x"6d7f7a66d5869cda", x"7aeadd3cfc38c4a7", x"41b92c83c73b10e4", x"b2cdb1642be2469c");
            when 32283810 => data <= (x"7a17ea4171f9025a", x"a15465720772b201", x"fdc3183c7fdbf708", x"a0ce9876d47fc700", x"1fbc7425b8317816", x"c304a4ff33b367ea", x"b816c1383c849d3d", x"bd6b99e262b206a3");
            when 22501300 => data <= (x"028c68f8ccf3795f", x"5c844a2897599e95", x"45a88034c51f8228", x"37fb6e30812ad4b9", x"9b9f0c7d618aac2f", x"70cd622c0e63c82b", x"1b88364caa5fd365", x"9f96e1ac27e0b969");
            when 4456939 => data <= (x"532c08519ebd04d7", x"a0f39eb9c2a6af7b", x"0f4b502e6b16cd14", x"de910a64aa23b2d1", x"14b3717689008cd9", x"2220846ad7bb633f", x"cee2343ff5c59658", x"d1fce72dc8eb656d");
            when 26889814 => data <= (x"419e1cf216814561", x"4403cd0553ca5256", x"43b5cdbf575753b3", x"9cd717f3353809fb", x"440cf52e2eea77cd", x"51ebb6080659062e", x"8c816ef02f7db05c", x"a9cbf6f795c510b7");
            when 4161170 => data <= (x"aa705cd7416d732a", x"345bd0e9af7b2b00", x"ee8df79f5e825513", x"2cdb4fbaccd55328", x"abfec0767034746d", x"169c45665aa4a6ad", x"1d654bc60926a623", x"60b70c9b7b3b6042");
            when 19570695 => data <= (x"0f2f96021f181a8d", x"5b67b414b7e1e614", x"d09663271a7721fd", x"fa32f25bbb16290e", x"1736f0fd8d7f6cb2", x"b3ee9ed04efec7b5", x"87491c96c5a2985b", x"6ad2719749f13c36");
            when 19283298 => data <= (x"9d4481dcc282c1fc", x"76e9a72357d460ed", x"e86fdfffb69b951f", x"cc3f6194a34d7d2a", x"8c45415218bc5747", x"56d53b5cdd034650", x"964a1fc162dd838b", x"ebf3b476b3dba734");
            when 6816291 => data <= (x"170c150d00c62271", x"99e034397569abce", x"91bf8e72c6a943bd", x"6db66cfa06154873", x"705d7665d97c0054", x"9cf82854cdb56ce0", x"93a669472539609b", x"0de615f09ba33ef4");
            when 14795537 => data <= (x"199a8ff72e9e22e4", x"1e589782c855293d", x"50f372d47d13dfc6", x"89b4e14e1e75556e", x"284b0894e4f0cbaa", x"5037eb9fe2bd6b7a", x"3b92c903b8920da8", x"95182e1077b687c6");
            when 15647950 => data <= (x"3a02b218fc99c8a9", x"3a2ae1f1ddc28808", x"ed8deca36bfda1ec", x"7c850f7a7ab61645", x"4618db2affe6af14", x"5c72b1f0969ab968", x"4d4afb79252dcdac", x"b3180de4441f02e7");
            when 8588915 => data <= (x"f3eeb40d65a2ead2", x"0d7e03e1a32e4861", x"7b81b36600642882", x"3154354a6b07ec3b", x"0e39fcc21e770cda", x"bbbf02ad09ecf7e5", x"d69b6b5b6fb49e46", x"5a313015d9368962");
            when 30937113 => data <= (x"76342097532c36ae", x"a82c6b6ae378b810", x"4de0c1d028a312f0", x"4e32972c57f96bcc", x"fb217f39a6a3de23", x"d484d0c0de422e7c", x"f29c6ae27dbfbefd", x"014537ae4f60cdd8");
            when 8735423 => data <= (x"6b27e93188066869", x"3f044620c35efe95", x"79adbe70fa53f1cb", x"80f3be0c26de2d53", x"82b8b37cb4f802e8", x"0314f547e37d376f", x"9cb52dc2518b7d73", x"3d35feab125fbe3f");
            when 23609776 => data <= (x"2bf4c27608bf2fd9", x"bf12c2ff0955698b", x"8e0826f993df1191", x"8302cd088f5eb30c", x"69b432ddc8541567", x"8fafa129aa13087e", x"23e494d5bd015327", x"c92498abdb412179");
            when 8610931 => data <= (x"49177e8b6a2e503b", x"290f81bc11fdaf9b", x"8b618a677e2dfc42", x"63a1c4bb7cf2cf9f", x"8c6107f2b9a4304f", x"448bfcfa9e1fc539", x"58eff2721df07e29", x"167e4f017e3bea2f");
            when 12139353 => data <= (x"7de70b31972b1a88", x"8ef9575d7eedd4e1", x"8a36e8c0bf674360", x"ca07caae5f4bd0ba", x"d76c5f2fa82aae5c", x"99fe488cb369815b", x"ecea3515cb252816", x"397caa23258b629f");
            when 3754249 => data <= (x"4b4773d75eba865a", x"a7533305b731cdbb", x"a0696227f629119a", x"c247f8f97ad4af47", x"61519c47c05b659d", x"710593c83e7c9dc2", x"5ec007f975264ae0", x"75173a771116c8c9");
            when 5661715 => data <= (x"e05fb368f6ac25b9", x"0edcdd7dc096e1b2", x"9f5221e601f76389", x"e9f197c896de82c1", x"5a61a4019872083d", x"8692a514196031a1", x"c766744f7db1f378", x"22e7ba9e69c0a466");
            when 2922800 => data <= (x"7c2cd4aac1ebffcf", x"866047bb9e8ab7fc", x"6a73c245b903009b", x"ce96fb78a52fd887", x"5dc3c709f978c856", x"58fab1cf2823f47a", x"77fb12ccbab82a3d", x"35a335941490869a");
            when 15928458 => data <= (x"433b7a4794c3e07c", x"7351ba991089076b", x"44ba291cfb38f2cc", x"bbf3ba224168b923", x"e1afe0773ed0de1f", x"f3985bb6ec5ed74c", x"ea0a4a144aa3925d", x"c094fd74992dc561");
            when 26462350 => data <= (x"aec4621b8629ef1f", x"021becfdf2a95c9d", x"d017bb7f18da62dd", x"c88a390d19368d6d", x"7ff186f9d0ece220", x"995a8921e53e9b0e", x"dc5adf79bf8a48a6", x"156985b09e74c075");
            when 13992996 => data <= (x"a2f9986dd83e5636", x"96bbe897cfb6550f", x"474f9bee1cfd95f1", x"2e08f8d1a0cf7621", x"b9397280dda883a7", x"f7909bc67aefd1f9", x"8ae96b4c24e9ce4b", x"4d203abf492161c1");
            when 14259532 => data <= (x"bdb2f7e2f206389c", x"7854fd85df075d3d", x"66d9c1a1de37b8b0", x"becb2172c2131346", x"8b1aa350b88b1123", x"7d41bcfea671e847", x"8ccdb77cc66d202c", x"9cfe5b64f2213069");
            when 21247038 => data <= (x"7cf143fee7e80574", x"79510e896a941a7d", x"a17588b2e036fb59", x"c6a099b02a224ea9", x"ab93d017b0e4c9a4", x"1b066adc5b3972f7", x"ac6efb97e19874d8", x"c69bd820fee35c2b");
            when 13725640 => data <= (x"8899c5d2a96f0c17", x"3c66cbe8257ad2e8", x"b139e8df6ad6d994", x"b15725ebecfebf3d", x"dc5f1fdc29048995", x"e46d80930572767d", x"84c09ec11b0c0f9d", x"4b83f5189dcea612");
            when 569602 => data <= (x"1bde003e51589534", x"98c94cb9565eb1a7", x"a8001e46e60b1b95", x"9bf526c05dd32213", x"5a6b1e9a7ed25199", x"97dc28df9007dec6", x"bbe5208ab80e915f", x"6f92f968a806c156");
            when 23464234 => data <= (x"9501fa3c17936bde", x"f9e3ae4307bd1e6e", x"ccaa91dbcf170faf", x"0d2b6b23c27b396c", x"cd0dd3b3093a52b3", x"1214fcf3f3447019", x"17d2f458ce5407ec", x"19cb7d547bfefe64");
            when 16068911 => data <= (x"bc8187516504f38b", x"47682f4cea4b8ef6", x"1745414b01aed62c", x"23a7a37b62232c29", x"06f1f7a12cd40f3d", x"a5f15510e8933608", x"a39621e593b645e6", x"45985abb87930fb6");
            when 21968545 => data <= (x"79447e926279c596", x"57055ce51c81bdce", x"91f09571a9b55c59", x"8889f3bdd3f3f07e", x"34b1aefa1af661ec", x"a6c9aec1ce197875", x"752ae8e626e56667", x"fafe4bf0c5f53c72");
            when 13739678 => data <= (x"95de83c1be173eb4", x"2ee2bb259f9b679b", x"71d3e13c36c31635", x"a05b4a64db42015d", x"1a43c6096abbdb5d", x"54dc217ec299567c", x"5a89e71774212708", x"b399698fa3e57121");
            when 10870849 => data <= (x"c8184e304e55671a", x"9f8c9fc80e8309ee", x"3e5c9d8973cb9bfe", x"290880726a97729f", x"6be958f818559275", x"3ffc1df4982fe1c1", x"52e53e625451fdee", x"a325bd49ae66c1a9");
            when 30132228 => data <= (x"7ae221e7afc18c01", x"1dc96581cd540f37", x"d54c369a6b3e822e", x"65504ef7505289d3", x"22b9cdf82ca8fc46", x"4dc093dae3fab010", x"53d21c67ebd0b6ec", x"dbf7c2ad7ba3751c");
            when 18350627 => data <= (x"df90de4ec0daa7d2", x"6c30e9db349abd52", x"ac1bcce9136686a0", x"9b06b06db43ac73d", x"c8f95ddee77b9f9b", x"a1ef3f91011ffeaa", x"d14c086eff004d97", x"0aa66109de9f5bc8");
            when 10784845 => data <= (x"d9b6cdf6a860f002", x"78a8a119e7f8a3e3", x"5f7eba4c77835051", x"9e4cce224f1d6078", x"59cfe958bc700a3c", x"d97c9e5197af305d", x"066fe0caaed0a51e", x"499ea46285c17e1f");
            when 16873708 => data <= (x"eab98f35fb234da7", x"21fcd9562e4a86e6", x"bac332c6fd6a6f1f", x"756ed7927cc666d5", x"eed9e8d8a1ac56d8", x"27a741db91de7a55", x"dbf87967900de917", x"2f8315627c5a5655");
            when 13804263 => data <= (x"e155ec35e89df04e", x"069ca309c0ab9fea", x"4a4c06679d25bbf3", x"0866ab7c83f11623", x"d14184544f8949d7", x"890b6789a3613b51", x"991315a65cae7a88", x"47471f497b1c4799");
            when 15683607 => data <= (x"8de5f0fdc3befd30", x"2a45f080cd411f6c", x"4c574917766c8bd0", x"abbf08e7de58dc20", x"65f2d595449aa93f", x"a812a168b061f064", x"3207e39b8dc3c41b", x"367260a7a1f1d941");
            when 15785589 => data <= (x"a5a35f2b92eb8e17", x"90c77ab8f9ac819f", x"02b60fd2a245745a", x"5608f98fc0936ea6", x"5b40fde76e33437a", x"4462303866d0bdc6", x"5ccd1f50e399d861", x"2b4669f011cfc956");
            when 21073054 => data <= (x"aa658181523ebefe", x"5e3956e4c7199448", x"0b1e7841e7a818ed", x"a22b6d9e9ac15bcc", x"0bf27a2deeee1410", x"79d9e077a69e5cd3", x"b472355029bc8dad", x"c3784bd2d3d0c009");
            when 11092753 => data <= (x"3320a5b4842890bc", x"7e855b03afcd54c6", x"11e1e62a4c457f94", x"c4d97023a8cece41", x"dc3318f097c8bde2", x"daca20a940c0b454", x"7ebc37ff2a5af0fd", x"b7eb2f5b12ae39ec");
            when 15518977 => data <= (x"ecf075df55fcdcf1", x"c5fc42a39525afa0", x"c9c99fefc9271b3f", x"39adda88208e7173", x"d06adfe2a3f5e4f5", x"ef894661bfc1e166", x"26dbe003581e182a", x"39fb7dbbb5c981ad");
            when 15660830 => data <= (x"69b8f359a6a9fff5", x"0ab885cd3b4b1f2a", x"ab16c203ae71f296", x"c63b4f40a8bda2aa", x"ea940d2c8678cef0", x"2e79abdf6cc64451", x"8ae1b0fe217c4789", x"d03e7c12523c87b3");
            when 17117285 => data <= (x"d7538542d2691ae4", x"b511c64409a05704", x"db9a6fe36d0e8cad", x"72a2068c60571811", x"6d1462472015167b", x"a82b77ebe9460081", x"e654d6f2c2b7fe87", x"8ba79b58958b7dad");
            when 15445595 => data <= (x"df285181f3355e00", x"3cf60aac7ce3951a", x"0a1e610e715dd193", x"0371200785695beb", x"ca67f35225245852", x"384152b3d1de4bbb", x"65deca24682011f4", x"9dc353644dc46a27");
            when 22824959 => data <= (x"a35d9db620afc4c0", x"bc90a3bae4efec1c", x"079b3551fa82f4c6", x"5a0f44ec09e37b8a", x"589a2b6ba5305aa3", x"a3f689dc522313ce", x"a944a6e94811781c", x"fc864899b63179de");
            when 22306145 => data <= (x"ae4185c1884d90e1", x"e061ff013bd3fe81", x"160c54fb5ab0a8b6", x"7c0f31631498e1f5", x"39cfb5bf7e0baa21", x"5aff2546c1573978", x"83479a0e351c3468", x"cf4064a3da8b2e13");
            when 16187086 => data <= (x"551e002a88b1946a", x"d1f63cdf30e88778", x"1b97d1eec5d28f54", x"28b7daac9f9fda98", x"98363c1272b47f34", x"276a602f40dbcdf6", x"750296d1fba454aa", x"762d1c405cc7d4a0");
            when 13773924 => data <= (x"d8f989b86b433e92", x"fc73878bcd49bf06", x"4cec82ed213bd156", x"037ce8a64a5e1c1f", x"4daa4441196ead91", x"75d4c93a19716b5e", x"a7d89aa57f609021", x"10bf003862a0b459");
            when 18862582 => data <= (x"9adbfc35f21f7b60", x"c9b64fec40003cd1", x"f53825aa011aacc3", x"84ba3b323dfb4625", x"bf0eb51779256ae8", x"c94b572e8c5d4d10", x"98e954cf8cebc206", x"634a3d3e1dea91ec");
            when 17155786 => data <= (x"2da1e324d86a709e", x"6f0da2ee5fe8cd09", x"0c2540f9716ce9e9", x"64072307bd731058", x"829c0691d375499c", x"f27fdf9866bfa012", x"bccb12cd6b59bef4", x"14366b3c09d39e07");
            when 24744213 => data <= (x"cc74b5a610f7de68", x"a71a7333f5d71ca0", x"041c8db68153523d", x"93a3a2630742e32c", x"3e286f7cf236e3ad", x"64cc4786c00f4ebc", x"6f32b1087c529738", x"8fc101a3b6b15c2e");
            when 6036118 => data <= (x"8758b0b563ddf283", x"c0a777752704a858", x"61918a9050621b5f", x"00b5a563873749d2", x"5321de84dbe83e75", x"25d15613562811da", x"cc8ec45ac15432f6", x"ebd3ae4dc012e6cf");
            when 23333019 => data <= (x"51d1a6646a7853c0", x"bcf1f2aa88b19908", x"3e66a43ac95cd44a", x"9c6817c157bde54c", x"9f847451e284a84a", x"08055cbcaac928ae", x"0f6effff51871717", x"9985e4f8cc475067");
            when 16637513 => data <= (x"72287d670b1d8350", x"790d6469ab12e92b", x"50dab59cdc49b54a", x"710bf9d84346c1fc", x"52e008c337e15032", x"f0b6f8090a343933", x"8754aa6d14dbb866", x"3000bf91f910d618");
            when 22264969 => data <= (x"66f5d39fde08655c", x"0938b75b62df36b4", x"0f25260d342e377b", x"699ed348e46ec912", x"d7a1e9aa42b07eb7", x"9769229ed834e559", x"1ecd8d713717bca4", x"a7681aa1b027de9f");
            when 19719812 => data <= (x"60dfde1ea1de4aa2", x"6f3ee384c24fd09c", x"8f28c998790ea087", x"a7efa7afd17a08a7", x"2bb7de2e4ff5173b", x"ba7170f22baa22e6", x"0b042f569ec12049", x"780f1bbd9f68054a");
            when 25059093 => data <= (x"5d6e106365e4fa5f", x"b6720536f691bb3e", x"158ea7f160d3d748", x"70506ce5a775b395", x"ffd173a2a6e27d10", x"d31694cd51b9b5cc", x"ddf46d91dfea22cb", x"9c0a18954d96b2cf");
            when 5201859 => data <= (x"b44f245528b03fbf", x"c362debebbd07337", x"c9535521445cee7c", x"ddb6484f3009ecbe", x"656504afdf897d3a", x"34621ee89a50f1e7", x"378a77b62665b2d5", x"54d945cd46250514");
            when 25497122 => data <= (x"a9cb8287b66c72fb", x"a9c0fecd2dd038b9", x"fdf3f1ac05b1bd13", x"d2e3dfcf538a3e7f", x"d48d13b6895d29ab", x"0f357d0a8ca04e16", x"50f0878d326e4210", x"18ea21518d4600e4");
            when 2826164 => data <= (x"db91cf32efdee48e", x"0f30293a6a5b8076", x"54b4c69b32c29d52", x"99cf4a0b36ab1171", x"de6296481384af8f", x"82a155f2a8400fde", x"e63ed06f78c31b2b", x"993fa1b3d5c836b9");
            when 14945647 => data <= (x"88afd6d056973fe7", x"8bd74ff61a8580ba", x"9738a01bf6c71afe", x"3ad676d28aba61f2", x"899bb6859e914c9a", x"1fea07169d550dc8", x"d3d3ab30c0179d51", x"f238e9d7b8ff6f6a");
            when 24612842 => data <= (x"01ed7d3f2fb2a7c8", x"05cb91be4aa911c0", x"bc8989c230a0d49f", x"7b3d48f0adf820f8", x"0dfb8e8a306eae94", x"d97a589afe9b520d", x"e84ca3ccc31b2df7", x"c7e8fff05cbfd318");
            when 20179129 => data <= (x"aeefcc5ac94ecabe", x"8b0c6b937a9622c9", x"6a81691ec42ac57a", x"be2300a9ec4f2551", x"d1c5e12efac6e6e0", x"f18e9be2931cce62", x"73c4a5caadd7cec7", x"851bb4042916de3d");
            when 9453136 => data <= (x"b1bf8b84282490c4", x"667a5948c205a36f", x"1e053f08891a19c7", x"8b0b8a8d70b9e326", x"cc5ce244633359bb", x"2d481c62d7bf55da", x"71e47b6364a4833d", x"2f22a9ac10133a62");
            when 31512387 => data <= (x"beb137b8c5839f58", x"268f27c1211760b0", x"f5905c518850e8f2", x"b0433694c5c5752e", x"a8b50123bf38ef60", x"e306f92715ffba7a", x"8d5306f2bb81c0f7", x"9c7b9f0ea5b9c332");
            when 10016496 => data <= (x"8d49974bd742a68c", x"3ecafe8ecd168aa7", x"5ea76939dccdc4ab", x"08c734da5a775bf2", x"524c82402b9cf78a", x"afd22c93fdd58085", x"f7d72635e2fc8e7a", x"93682574d53bcdb3");
            when 6415834 => data <= (x"1946bebd0b8600c3", x"05c9a22ea7e25196", x"2183d6b49ade1276", x"fc2c70aefee96d74", x"330123156d8b0207", x"e476f7353be2cee6", x"10c5c2287c1602a0", x"fcaeff074076ee4f");
            when 1895526 => data <= (x"72234dfde87df48b", x"ff31b4dcda40be12", x"40e898e3308b58ea", x"39f1e225e843f805", x"87e33f6ea8ce5ec9", x"cfe5a212d770fdb2", x"86bacdf150b83cbf", x"bfdb604963c3e1cc");
            when 20192494 => data <= (x"a4f727e6966cf6a6", x"a9825f108b1075f4", x"5d6f9378aade3832", x"2cb23b837293efa5", x"df9b96b6170fdc91", x"f429915981586438", x"24b7b2c732131eec", x"9b013369b72e9c9d");
            when 25873035 => data <= (x"3cc35132ea0790ea", x"6a6d0c22e917d845", x"072afb53fc57086c", x"abfb87155fc98b5e", x"028423b54ff7baec", x"827f7bb7dd462cb5", x"a65dffa08d0111b0", x"df79858a6ad836a5");
            when 12391595 => data <= (x"dadb7be8826071f4", x"3ce10f8e0ab18857", x"4e0ade526dc43fd8", x"8f1902b73d3aa73f", x"3b422c22c9be6514", x"fdf939ae0405396f", x"779f62c3320f1b27", x"7c4130be7876ca2f");
            when 1959234 => data <= (x"8168f1cab67c4742", x"d1ef204a069f6df1", x"7a1452f98c6b2405", x"f2f759bf1a09ca2d", x"2f5f27ef609aa515", x"927d26ee9ebceaed", x"a507dcfb862a2847", x"b8ec8a6fd7d81795");
            when 6562184 => data <= (x"830f2d7f618369dc", x"618aacca7a1fe311", x"fdf3fe41dead3861", x"b01170dce0aac8e6", x"c3609938faafdb88", x"fd5b255a0dc0af92", x"5e2d93a0e98d7f26", x"92326a6faca5a241");
            when 20827168 => data <= (x"09b83c8a1baa6efb", x"8f220384bb68dd54", x"071f5a2cb0db7cc4", x"36e6b9103824fd22", x"be2914dc1f1abb94", x"64b486668fe0b970", x"ad1247f3ed234a01", x"d32e7188ee9fb853");
            when 5598937 => data <= (x"60c4e97f0086d80a", x"6d91fa505801fa32", x"f49b256229716ded", x"3c9786614320aedc", x"3989adcaa4d3d616", x"4d7caafeb1cc4abc", x"a6f8f3fa0f002c2f", x"2bbb2efb555a0919");
            when 6673301 => data <= (x"8a6c59b887a08f30", x"3f6f7c289b9e914c", x"13f9fcdba56666bf", x"270b386a60e094d3", x"94b3c5f4837f75d7", x"3003364401d07186", x"244a13bfc0de9c95", x"d25f1726a3f38e66");
            when 1901552 => data <= (x"d0fcf05b9621aa36", x"d5a1007375c08e07", x"0ce110401d940f36", x"e8e14134f801a70e", x"04efc465a6a4dfd8", x"312d20769f92ec9e", x"a7bf7552f19e9768", x"e6cfcf1913d09bde");
            when 16315876 => data <= (x"70c1564198804cd0", x"db6ab56aa8dd4fae", x"54a2775e72fb8aa7", x"e8ea6d9bf387b2c8", x"cd9b5785b016ad05", x"a50a1cc99db38c97", x"d97504d8c6d51b9c", x"f958d98982696a8c");
            when 24413190 => data <= (x"6ef18cbf8fae84d1", x"f21b80ec508fdfa8", x"8fcda6e217098f3d", x"1bf12b87bc0915e0", x"74c37f11c0db4b95", x"3e255faa769938df", x"e4223d1f64042375", x"17b735874c3294e5");
            when 18023408 => data <= (x"c0470585221c10b5", x"7d79e5d88e5074cc", x"26800ec9d7838002", x"71ad06bd514b72b6", x"e19e4e241fd75fa5", x"f206cde81893401d", x"c17b1b0da2d36130", x"3fd19b3ef477007d");
            when 28466906 => data <= (x"2ad879a2f9843b65", x"37ab1906b8f6a860", x"a2fad705e8b2fb01", x"47f5d65a4a749b8c", x"dd9f2d4492a43716", x"5dff0edebbeb0b41", x"a4c98dee3c466f0c", x"4eafbdf4d97dcbda");
            when 5142712 => data <= (x"81ebc497861619cd", x"2984f2f74b128aca", x"5918af850eae8fd3", x"01d3fe4250f31700", x"9a5724d36625505b", x"7461448ea9461807", x"b4033d2f80abc5c8", x"ac34e13f05ca2333");
            when 10928204 => data <= (x"bb2b141ad7f91398", x"00df4715935b9552", x"224b13d376dc56a6", x"d1f4617374f7e718", x"fd9227824d620377", x"f9150cac9132d9cb", x"079a2a5079ca84eb", x"805b5c2e003ef65c");
            when 18218409 => data <= (x"03f0e28bd19dbff1", x"cccb89329f15da90", x"2a0311c15cd2b240", x"8039270aae02d993", x"c1e683f16a6f518d", x"984fc27007e08987", x"d1f3311881d9e77b", x"619492d4f3015e85");
            when 18460051 => data <= (x"4c35370cea383647", x"244bc26e76617f43", x"b6efafd12d4a4124", x"0eed2b83d22f8103", x"56c9302018dd067c", x"7312e019034ff333", x"d7b8b2298520bbcc", x"8f97b55baf00e689");
            when 16880998 => data <= (x"ad9a4b6ccf269186", x"fbcd4b1ca304114d", x"b232d2ec8832233c", x"8a241993556c27e6", x"ee2eea22e3d6314c", x"bf5c97948d6f67c1", x"ae7b60c6872d09b4", x"1439606b0d0fab77");
            when 21714998 => data <= (x"c72be7219e066278", x"60511f0567b57ad9", x"1d3b817aac2bf1d1", x"bdf4dfaeca81c942", x"a943dc7a2cab5318", x"79584707f03383b0", x"d3a4d2dace48d763", x"06cbc0502914a0cf");
            when 32019544 => data <= (x"3c4ff19df470e434", x"dfad8f32eca37577", x"5c12c0f0bcc4dcab", x"629ace8e31fbccc5", x"3c940c3c68924cec", x"f783fc3a0432cca4", x"5dbb404e6d41f124", x"e866fadaea78c5f9");
            when 11063288 => data <= (x"0ff6ad4bedae89e7", x"f0120e0c7134586e", x"ac10035bf80f3b09", x"62ba478ae1034e1a", x"a74990c79a8fc077", x"8e6e82ce606061f3", x"fb499e78856736ee", x"20bb59cddc178946");
            when 30138068 => data <= (x"ce21d6760c923e5b", x"29403ce6fb08f6fd", x"ad13e112ec68964c", x"fbaf8a7da2db5716", x"80c443d24e294283", x"74cb83cfc9b99019", x"88c772e7ed231013", x"25e315cff7dc66c8");
            when 31953709 => data <= (x"65631e84ca0318a4", x"bf367b8b3301160f", x"9794a49dc5ed3b1b", x"c3d30f514a0111ea", x"7fabca31f4234f01", x"c07a86dc2d9b7597", x"33d0411b1fb4dedc", x"50a977d6dc43cabe");
            when 488228 => data <= (x"ad02da80f82fe89e", x"bb114ed248b382f1", x"f5f1012c61fee539", x"6f5a60113a953d27", x"0762b957931d9dbd", x"1b0dfc1d835ed79e", x"7d71f94fa62f71ab", x"ce0f2e194baa4076");
            when 3010718 => data <= (x"20c82a0106f2b13d", x"ffd5663da875bb85", x"47b45931d3d8dcbf", x"4e6482182c1b9005", x"c3b762e7857bd7bf", x"9850cc2a12c09db1", x"75489db84b9e185c", x"0e5c038d5f96f350");
            when 17021974 => data <= (x"f0e2740b0ce3268b", x"2f5d5a1b73c9ab26", x"1aaa5b03cf590f23", x"6b37622ec7eecb0f", x"6b31a2260ac761b6", x"2780d48204d30458", x"1cdf6a920f11c93b", x"6e6d7ffaa607e34a");
            when 1156539 => data <= (x"cee5b8f9383db2a5", x"b864c5d1a79e0e91", x"2311b115491e0bc4", x"d7d046ef409633b4", x"ea68a24cc722be9d", x"2dbc39ea4f658c01", x"fd5dfd259495bce8", x"e18ccb531a6f7cf9");
            when 28170762 => data <= (x"ad706deea58f15fe", x"796b3ecbdfd2fec6", x"9b85df8240dbea7b", x"30be0b0681c83a4e", x"66f9591785cbfc88", x"1943e40b04a564fb", x"912103b71da638fd", x"77726997a2348967");
            when 6211898 => data <= (x"2f6107a5012e08ba", x"c5cdfa9bbb0f84fc", x"2df9352e6d1877ed", x"cadacfa3499b17c6", x"8f21ba87055a2e5a", x"cd051e7bbd5eba99", x"c869ba4e9dea0447", x"30dfb0582e5c1c52");
            when 9165521 => data <= (x"27ed3b79f05821fd", x"9b4548c44d0eb3ab", x"0959e4a15dc367c9", x"98a2404a8c328068", x"75656d300320e20a", x"e225f4fef85cbe3a", x"239009199609845f", x"dc41595dba12e208");
            when 31437996 => data <= (x"eb1d029134d19017", x"b706663d4e7436c8", x"fb306d05e309d27d", x"c0ea128c0efbc8f5", x"ff4cec452d42925d", x"1b6fbdcf6669f7c0", x"df03a343ce8f9cd9", x"48513a920b2256e1");
            when 28054165 => data <= (x"7175b1433a79df8f", x"b32ad0447cd6b66a", x"0652947f974602a0", x"445e0eb439ab8484", x"c66f0019ea6d0f6f", x"091947b2a55523ab", x"e4390bb09595b527", x"b05ccc8775dbe205");
            when 27117059 => data <= (x"1764d8262dbe268d", x"cd5f5a1faac6464c", x"9bf72f5a69c0cae1", x"104874f56288e2ae", x"1ff3d90d6fde73ca", x"535009f6facae06b", x"e48bcc03f6c447c9", x"510a8cb5bc5a233f");
            when 14802183 => data <= (x"de49bbe09c156d92", x"7cfba56b4f539b0e", x"52da5ab6731b95fe", x"cdf5bf1cf27092b5", x"819766a9c7e94382", x"733cd89125f7ba9a", x"91d0c4418353e219", x"bc745161c4f49b62");
            when 8233346 => data <= (x"89bb24ad52ee8198", x"dae0319334fd82b8", x"1c507561ab982831", x"1c47f7d316bf5356", x"e1ede0644a9b81b8", x"d3ad2ccc4a6f0251", x"9bf3e8b0c29a3ef0", x"25ec41f2b77e2c54");
            when 18003374 => data <= (x"2ce518927bc224e7", x"19cedfccfe9b6361", x"cae90b8bfb14e318", x"64ce228c3cf3ed35", x"7e04fe530b671755", x"6e1a1f37633eb42a", x"78e4bd1ca6cd26b2", x"dfac440bc428b0e8");
            when 32998737 => data <= (x"cd4e3b0699cc3af4", x"6635a1a8a54b1a4b", x"7fdb00208a6088cd", x"971c57803d3ac6c1", x"a4bfbee7607bf6c0", x"8188318779bd88f6", x"384807fffd90b9dd", x"570327bb0aa9900d");
            when 14467993 => data <= (x"bb0845d37b2d1f5a", x"782ebf8f685c1f2e", x"394fabca2de4671f", x"0b2b78b9d5e51ffc", x"799f5129b5a3702e", x"781c439ec1916d65", x"29133c629126c69a", x"53a835f01ce3edc8");
            when 21995722 => data <= (x"4b1feb470ae07b1a", x"daf617e9bb9d6a64", x"4533f1c91e5aa316", x"2e505e17fb1ef9cb", x"67af5dd2b425d4ad", x"5b0250a287bc4521", x"bd172a9687591c59", x"6376b5b374fb7752");
            when 5495741 => data <= (x"97c5ec2d0e07b1ac", x"d3e66439cefd1bbb", x"8185a2eb4f3b757f", x"e9640a34b9035229", x"08207d46f08e457a", x"bd81eb310769be2a", x"2da2c2c89179ab5a", x"7c0b6da3ea6392ce");
            when 16458851 => data <= (x"35b1406eb59be906", x"922b1c6492901824", x"16ab9540b6165441", x"0940f9c7a2e87c5f", x"122639365872fd11", x"60f35c48e7fc8131", x"69a017e44a615ef3", x"fd53e3fd1a195abc");
            when 22154772 => data <= (x"6c2fe0bb77af9b49", x"842af734af691f7b", x"002f7bf1f3a32a28", x"6c87bb39ce697a31", x"a0557d6469452f3a", x"4e0a9c873c0b5a3c", x"dda82f15791b8c96", x"474f062bef9134f2");
            when 30066556 => data <= (x"90bc2cddbd3c5c5d", x"9bbcabdef48e931b", x"912a983718e55c59", x"425c3d39e99ab798", x"5fddc28cde37d48a", x"62e65796f8e1af6c", x"f5667679965f7d82", x"fb7406d833ac5260");
            when 9348627 => data <= (x"89f034a852a75a8c", x"b6281bf87540a023", x"3446b5dca56e53cb", x"5e4436028a6270bf", x"aa077752f6375095", x"8a685eaaefb5c4f4", x"59b2317ce776bc44", x"8b07ca7eb0a15f4b");
            when 5139002 => data <= (x"36354866c039b999", x"f39866b78cbab814", x"7572f7e6bef9a50c", x"ec1f4107d6dc33f4", x"4cb266c494e1e2da", x"21f50e0adb2b348b", x"15aeb1d87a585d3f", x"7feaac0127711fc2");
            when 3965493 => data <= (x"8679e84552e6717f", x"0a0083260a4d9310", x"c7bb7d0702346eb9", x"2bbf8bbf1eeb4928", x"29b137e4f0d88db3", x"56d34718cf7ebd64", x"97d0106e5da0be23", x"5e544b0da5580a17");
            when 8957604 => data <= (x"4dece97b10f310ab", x"f3a00ba81c049717", x"500b2abdf9929ada", x"e00bb8086e0d96d2", x"7144d0e3a3fe28b7", x"f1deca27b0e34021", x"6b71c9eacf98f5e7", x"e0d040e6e8dd8e4c");
            when 11900980 => data <= (x"36ed843db151d199", x"2e018c7dad8e214d", x"a33aff2eef8a88c5", x"b781edb4138cdd82", x"715ac44493cd9d63", x"1213c39a265e2cf0", x"516a4e711a966281", x"1d8dc7916c432e72");
            when 3246584 => data <= (x"01681669ce026f48", x"d688db17b1ce684c", x"41b09a487c54c3ea", x"2651c3f0bbc29681", x"614cb98ec8ddcf19", x"6433a8bf167f0deb", x"303a49088edd0a96", x"b17c938915ba7ac4");
            when 14310410 => data <= (x"e7279a06a83f549a", x"d9c9c1744390e04f", x"840e364c457468c2", x"31238a52808b010d", x"0de14f3eb762ee40", x"fa2e45a340dbca38", x"f43e2df16fc40d28", x"e63e5b5fbfc5f945");
            when 9658042 => data <= (x"8f088654cbce67c0", x"292243711741bf98", x"59fe55f783d575f4", x"3e71c67f0eeac0f2", x"6b24fff62bfd9b89", x"f47cdde9a5a74a8b", x"df8d858c8493e05a", x"aa779ce796384fba");
            when 23939998 => data <= (x"a485c92413af65a5", x"85b41eeb20d5f167", x"f0cdb16263bdfeb0", x"f8fe7fef25e6ac7e", x"b4e4973de76b3e71", x"df1d06d23d424dbb", x"a9d98a4667d40e59", x"daa328c0b3fc24c4");
            when 18946352 => data <= (x"bdc7bd395f1b5a0c", x"083054e5cc8f1ed3", x"d4426eac8a8dcdcc", x"22e15894ecaefd45", x"573035ae8f66bf1b", x"5e6867f37822d66e", x"1bd578db2a290daa", x"00859ece9da019d5");
            when 9424535 => data <= (x"574e0a4333154084", x"5509a29df54c33f7", x"83f225c64d972da4", x"b752bf0391085903", x"a9766a99aad78664", x"37cfc248136fb060", x"25289d6a9fc06b47", x"0bc9bf65ccb36c42");
            when 1209587 => data <= (x"0e5c7f8ee9498989", x"b43a7123c7707d8e", x"c42aff457e754cdf", x"1571c6550a5e0992", x"cc1f7d718359c2ef", x"4d810977a1f59d83", x"486968fc764e205a", x"78c5a31f5414fb8f");
            when 33604850 => data <= (x"55195504f13265d7", x"01fc3ea19ab2de12", x"a05af57cd0ff1304", x"9541ff6c96cd8214", x"cb7e21f98255c1cd", x"e97a29e5082fcf9a", x"ab272fad7e714643", x"e32df21b393cbffb");
            when 25176947 => data <= (x"4d2e01707cfcbfb0", x"21e9c05c408dec89", x"87d40ee9e108d577", x"29b5cd0bf21c2ca1", x"71e685dd2c917f83", x"a892d214df999063", x"93c4400e44e4437a", x"d24a8063ed0cddd3");
            when 14691599 => data <= (x"6f31a12c8ce7a3e5", x"b7048d93310e1d18", x"413899a9fe4922bc", x"c1e25a8c4bd70234", x"c65df20895a27cef", x"3979aacdd1856ecd", x"b767c5e2c95f8ca8", x"7192141ba8b865cc");
            when 18309574 => data <= (x"db63664a7216d734", x"29efdb79cfbbe1e2", x"ecfbe27e88fa3d47", x"34750ff77245ac89", x"1792d42745798cb8", x"3186953d907819a4", x"7099f377aa9d4295", x"02c2d4944ca3da75");
            when 25744611 => data <= (x"918e24edbca72ccf", x"1a3f2a4bc543f599", x"3229d3b726fdc3a2", x"3193ff357219eb64", x"7596d14f6eb5c6b5", x"f38c9ebf3a383e72", x"1458ec6cb3a1f88e", x"0e3094059fcc1fba");
            when 2792198 => data <= (x"d253254ef4f008d9", x"bed6e38af1a2cfbf", x"106adba271d57d13", x"a6c469e3455b87d9", x"fb97269a0620f375", x"9d58c39cff1c259e", x"7974820228252d26", x"f3922ee8814b04fe");
            when 28427787 => data <= (x"3e62990faaa56caa", x"c1dbfaf29e04b90f", x"6069d583c73187c4", x"57bfc775e70f088a", x"150901d5f1f8c4a5", x"6ed9c41d9621bbaf", x"dd153a0ed2ec44f6", x"db4c676db06316b2");
            when 12889041 => data <= (x"4b65dbd9f3f80a11", x"c8bb11102c4a0ca8", x"7845ff9861b72049", x"5c08d4667d242648", x"ef4ed920391d6d42", x"0dac6e74cd317f97", x"59155ad2b693335c", x"d23229c6aebaa2c9");
            when 17566683 => data <= (x"42f748d8f121738f", x"60f2f64bdfa4c20c", x"68f8f486430d49f6", x"271ad9d0cbe0c04c", x"64da94dc4e3a5660", x"e03d44f0a1067390", x"7afd30b0d61b8eef", x"7c34ed97132a5cd9");
            when 23406661 => data <= (x"709a80e203e39311", x"f679cb41867be386", x"348324a7a2f7c5c6", x"904258ff00bd9467", x"ee6572a180859539", x"2b525170211d2f23", x"402aba2d6a39bc72", x"c3995d70f8c3761b");
            when 25694517 => data <= (x"98bf425f5146045c", x"d4a66ac24d257c7d", x"b5889aa257a864d6", x"cb121e7e36104f76", x"98495f2684cc4fa6", x"6b0fea50f5ef06c7", x"a29d49b89cd43015", x"e8edfeee4fb3a22d");
            when 24740590 => data <= (x"26a880df2c4b90b4", x"48952ba0aa7552be", x"eecb3f76278b5bdb", x"699bbb904cd25db5", x"51cfa3eede9133c3", x"8b501aa18a73a613", x"d2ad8d2aca5d6a26", x"7d544710aded1042");
            when 28708804 => data <= (x"9cbab27ccffe04cb", x"79aeba1276151131", x"f1d521b29be63f0d", x"4c8f9f68f59cc239", x"77e696949c2b0132", x"502a1be444906409", x"97b1d9a417bb0a6a", x"04ca6381210456c6");
            when 26632751 => data <= (x"89ff69542f904461", x"aa07e50d48c6a44b", x"05140ab97c9da76e", x"12c8a1415fb34a86", x"136cf9bcd1a07c10", x"016fe3c56c34cd92", x"d026c889facd3ea6", x"8d7ecfd8aa69d2fb");
            when 12253071 => data <= (x"2425eee77c645859", x"ea2e77c634533c84", x"e20d46a3577f65c6", x"1e0638f30524f4fe", x"56dda069f3662758", x"cbee7b780f1b5134", x"dd0cd05cb3ff6130", x"9568a6278d523767");
            when 25231587 => data <= (x"63ee20cb1f1c4cbf", x"25b7e909ad2656fb", x"4e58ae430ad3f3c6", x"3a18f5cc9901510a", x"0301fc19dc588162", x"e8d172e416dc20c7", x"ef14d14fb584d1ea", x"ef931c087381e1ab");
            when 7191221 => data <= (x"5c40c8d176389bde", x"e69809a114f29724", x"6db51f26e27ec762", x"003884a81fa710c2", x"7bf10c12c0d1dc4a", x"83a7b00ca53a7f45", x"2de192bed4c48a4d", x"8deb5d47e854aea4");
            when 31253932 => data <= (x"6988ad32344aa93d", x"7e6dc50e54d4ace9", x"360842d4ea61360e", x"d7d9e907c99d8942", x"27d0aa2654b124a8", x"6c56a05b06249603", x"2cdb3a3ed5cd0d11", x"95901f5f0f526b7b");
            when 31815433 => data <= (x"1c7c629fb0a2db93", x"18ed1fab00bc8160", x"abebd613904e2f0b", x"5b3fbdc24388b99d", x"58c1e01ae8a9069e", x"d41075afff8d7842", x"7f33d0ce3525f27b", x"d663a1c54364932b");
            when 22861694 => data <= (x"211263080befd465", x"1dc7d3f8a9cf2a29", x"e1c5cfcb19ea26b3", x"454c6efe5db8907e", x"a5f7ff9defa74fb1", x"a894c94eefdb3e6e", x"b5a3c79db58972e5", x"636b7a21fd1f1587");
            when 13627294 => data <= (x"4b0a0d223ee53387", x"f82fcebf064297e6", x"b330bd2ef9f74cf4", x"83d1249c5241a538", x"3a5d95bb8f68d1bb", x"bbe96ff839510ae0", x"0c1e38f0c27abe7c", x"33639d270fb8fbf1");
            when 14407910 => data <= (x"9fabde8e52d52469", x"ac5c456bfa5f48fd", x"b98dd02d81e4522c", x"0257cd9bd9733bdf", x"4daaf609a2c2c3c7", x"0888213a24720ac1", x"1a1f4c7a72254d43", x"c62900c43f481d68");
            when 30400287 => data <= (x"1ee5bcac5b8c3316", x"478c212ca3010709", x"78cfa756ad7e1323", x"4ec04624b6fa3ef3", x"87bf14bce3ca0b45", x"a53deb7f072413f3", x"f6725187376d18ae", x"c34a9e13c25d8a8a");
            when 22649637 => data <= (x"8c06119df92a8b21", x"ea03595f994ae8bd", x"488000c849e45649", x"2ab51a929bd37e1c", x"c43cb0d050665c73", x"69e19e0100e24b0b", x"085e2d6e3e73d8cb", x"8593f52bc7393d50");
            when 25307872 => data <= (x"8e3dea963812996d", x"499aa4abffb267e6", x"0b73901cbbb03f7d", x"dd77fa526fce841a", x"820424a2047fed53", x"6bd077fbc60d622e", x"ba7d490646567c65", x"fa81e1866c36d6d8");
            when 24657727 => data <= (x"4ebe13e657f11af2", x"79b0d11f808dea65", x"cc8c2983a746da9f", x"aa5cad9a176b8242", x"7cd4a8744332194d", x"47f4d2e328a80f0f", x"e41a9b699771a642", x"3da32c51b11b1a63");
            when 3455746 => data <= (x"29277c9f773ffdc8", x"1f6710652d4f0685", x"647bd346c12bf348", x"57a76c5ee0d344ec", x"9fdd6d6ba0694535", x"52321b3d1adf90eb", x"70cdbc30ebe640b5", x"3b3dda4886d0fe75");
            when 26793996 => data <= (x"e49dc1571cf8036d", x"7581477049fc55ae", x"63e095eb9ec2139e", x"0582145be8c4be9e", x"cecdc9bfd6636b7c", x"7bc3295b5f3b4713", x"a2582a7e8741b7ca", x"0df14354c9db2cd9");
            when 10700296 => data <= (x"09fb65911f1ed953", x"3172fcc5d65562a0", x"07cd1d7b2f956259", x"c13c8862360e07ec", x"f637ed38a11b7159", x"83c92ab36ada1a9d", x"aec05028639f7d8d", x"063dcedea52b63da");
            when 25897773 => data <= (x"a22cc6c609bb6b4d", x"812acbbeec8bdc7b", x"028f771e4eaa4364", x"932e1239b7f4f567", x"55206d2f2d106ac1", x"5d9fcde3fe32722d", x"23e2044fe71345a4", x"d41a5fdb4cbe95a1");
            when 10158043 => data <= (x"2a81aba05bf98ee7", x"b20683cbcda36504", x"67741d3e032d6e89", x"1321a470347439d0", x"6b0a1600b692f756", x"a6ec7a5efeb7a124", x"16bd62d8a0648833", x"6d61df9ead27ce9a");
            when 16600514 => data <= (x"4186b4ee4431de41", x"c9e2d5969d2e6c12", x"e77e15f4e1161457", x"0ed154ff6a451647", x"7fdacb94c72091ac", x"73703a35d22a08d3", x"cbdd341ed8a6a5d4", x"ed23262fca32a295");
            when 14766492 => data <= (x"fbe0dd8d878a6515", x"887a04cf765ccbc9", x"2c6786a726e55811", x"849df77d98505e17", x"b98c3a490820f6be", x"971b0d645204c371", x"2693c0f4862b8384", x"9078d6e59e9802e6");
            when 11968279 => data <= (x"8b2e8ad8d36928b3", x"baf1bfecd9e2d444", x"ddd14cdbbdc0796f", x"bc4165064b55c68d", x"c74d9ab62c8a1d1f", x"f2bbe788fb0b7804", x"d11e2bd603bb45ce", x"ad5768ac895899e4");
            when 8910867 => data <= (x"c19b89f3e9d87a34", x"62eddbad24ec5275", x"57e0942fc0fa104d", x"191324d7d4777aa8", x"f5bdb2d6371247d0", x"1020c12715958803", x"295f3ef0829e563c", x"4d558b7138fa70fa");
            when 25460556 => data <= (x"fcc1fed3577f9e18", x"3ebdf58113806a6e", x"3cadc84df82c94c3", x"511f9708b916f7b0", x"1463b6d23965144a", x"98808b368b48e1f6", x"a6cb7061168209db", x"d3b3ec9e004ed483");
            when 16021028 => data <= (x"a32631dabc012e01", x"f3e385eb3c544749", x"95aef05725da6feb", x"b5a31f07d2498f47", x"7b4f835584354b26", x"5e0006c330dff2f8", x"88ee4ab687d82744", x"6b4126d5a54c43f0");
            when 20626796 => data <= (x"7344e55eab239f29", x"a4e36a3697f71d58", x"eed611280b6cbe92", x"665be71e82862f41", x"8dae32eae2a38c79", x"8393b2f9f156e412", x"29ac8656729e831a", x"e80e543fada494d3");
            when 19596089 => data <= (x"36ab78abf08e48c5", x"5acc09d8a579856e", x"4db1a98502cd6ebc", x"849efe76554c9f21", x"6bc3cc4d42ba660a", x"e943933ceb846140", x"a08ddb3e434e9db7", x"7583073c205c417a");
            when 26930941 => data <= (x"94c8bf7ae1a7b1e2", x"28c5604cf63b8f68", x"0fbd6bbcd05cb780", x"e14bd843a5c53c76", x"b3b5d7b586b45d2f", x"8adfd151567db711", x"b489a5a598f04a6b", x"3375002933cb2a4d");
            when 15110947 => data <= (x"14d28979d519b9a8", x"06f919877f19438b", x"1dfd48ac4a0d96d0", x"7a6d3c772f241474", x"3426101184a3e585", x"3a6af3f5dce7edc2", x"3c09f5b76d3a7fb9", x"f1aef17fd4294b7b");
            when 3292246 => data <= (x"30d0225cfb16e78e", x"9a5d695a56183ebc", x"b6c2d923f9f4c9a1", x"2fda9d08081cf9ef", x"b8cee5d55953a944", x"3f574ace4b9d1258", x"3400c0b2814ff314", x"24e847141c7401c9");
            when 1864625 => data <= (x"2f121777359331a7", x"0034f6011a367b7b", x"37f8b3f8b09715ee", x"a9d52b0ecfb1cb3e", x"8bb55414b0305d21", x"71ff4d73c3670a0c", x"52583d9f5bd049f3", x"fd642d0517f6e8a8");
            when 12168465 => data <= (x"0da248633d5e85a3", x"997c750133695dba", x"335c6ae18644d951", x"02ff0c7f2d5d7037", x"ea727ee48d83413e", x"8ee0840913bc119f", x"e0ac86f951e1ae1a", x"7ec3578265abf335");
            when 23554382 => data <= (x"b26e31a2a608b184", x"79383899f40f42ec", x"4cf19d17fb780bce", x"5d376cee1cd50f5c", x"73978edf8f962fab", x"08573b1a017568c3", x"c3cfff417058456d", x"e067379ea23da7e5");
            when 22517904 => data <= (x"ce10784147ce06c3", x"8e4e665d6f394be2", x"03a54b9db5d4e2ca", x"b0a35d2175aece55", x"ac7ee51d1b8d92a0", x"d40775b40c35cac3", x"038258bcf5003f1c", x"ba0b0f3aa920f96f");
            when 23929377 => data <= (x"0187755c625890c9", x"41c159f6bdecac5d", x"7d41af21d91ca002", x"9f3e58889ff200ca", x"bacac9a3bbe397cb", x"41cc81d36ee209c1", x"3ebac5f17e2f0bc3", x"6fa7804897b68e89");
            when 7478079 => data <= (x"3f58139256e7c78b", x"6909c23be11ca9e4", x"f5dbafba4d0fc10f", x"1ffeedd85aae372d", x"3826051b0373c029", x"aa6591623818981d", x"a44b10006cabe04e", x"11d5b7b29e93ccd6");
            when 19666514 => data <= (x"d154ce56de6fc8c0", x"a121500a35c44ae7", x"eaa1f0ce717dbed9", x"19d16207e72c5107", x"a64f43d5d2a1519f", x"d200d91ddec98309", x"ab118925dedbd7a2", x"543de896aed327e0");
            when 26379779 => data <= (x"b000dbddd7e10472", x"9b892fe2d00f8a4a", x"efbc3e41695bd292", x"1931f78f55794580", x"290546ba2275402b", x"537cffa336da01f5", x"cef0984b976973e2", x"6bbe52bfc2af00b8");
            when 8715955 => data <= (x"771a72103ea0c6d9", x"c38156db923cedd0", x"5db627f9175a1ab1", x"468464526a9f06df", x"cd6f130b6b51a61f", x"82e522b96b436767", x"e54f688e6f831956", x"cf8932aff719e3bf");
            when 19477073 => data <= (x"b100d992beda5dcf", x"b7dd96a1fd25803e", x"c84d018b05743fbe", x"28e596fc758e1fe9", x"a775b5dff2a689e3", x"cd0d513c12eb44c6", x"37acf2b5c9c1efa2", x"59fe3abd18fadb12");
            when 25942713 => data <= (x"b005b35c1d21d1a1", x"015101aefa87d07a", x"bad5c45c656d9e0b", x"9a945ff361d36b9c", x"9ce7f58707208ace", x"25f8466db0ec5bb9", x"ca068d40a82333f7", x"7df95c137e5a6d48");
            when 13611254 => data <= (x"b949dc8d6c53441e", x"65ea719d70ede1fc", x"cf79492c09dd0624", x"8cfa99d4a5f432fe", x"a28d885e37101706", x"591128d53b28766c", x"dba78fd955a8b322", x"52e735acd630cf83");
            when 6700705 => data <= (x"0342b4553b71fc5b", x"e1dbab7d92d3dfd6", x"c96a7f75a61b6621", x"de684e5407abba99", x"4513b208b45c5401", x"393c8f1ee056f891", x"fef4734ee0c36195", x"1f4720c75ec944f1");
            when 1302695 => data <= (x"65a9154eea745229", x"e36d55235183316b", x"693c68feacdd309e", x"301968f70ee2a403", x"129d57ba3225f1f4", x"4d3e5e210411ef72", x"84fd99916b4e894d", x"8db0c25c0a3a1424");
            when 31855031 => data <= (x"48284c9c9588d2d2", x"2a7bec2ccde8d765", x"8523a335653e0b81", x"172a13f1ffda0149", x"957a44c0e5c46537", x"78359c41d95c8c06", x"1149a8a8995e1fe0", x"4340c2fcefe16150");
            when 15331305 => data <= (x"deb885471f5ba7fe", x"a47e3976258b6b20", x"23bbbc86b37632e0", x"3291008d640949b5", x"1e285816858cf5a2", x"ffa7700f6b98f0ee", x"bb602a1ab0837c13", x"0e3361de5b0f870f");
            when 4793942 => data <= (x"d603d45ea75383b4", x"f3023c2753e35066", x"8ac184352adea853", x"0d3e0958bb7720de", x"79ceef4bb3c6a2b6", x"ab4e137d43ec8bee", x"2009570ff5b70cb4", x"0ba15cc8901a50d4");
            when 3790209 => data <= (x"c8572a906921a586", x"8c3cd53f94788dc1", x"f7284f6586729ea0", x"c5b62af8f5f0ec96", x"baedfe316a81e950", x"e9709ba59aea6c99", x"5b0e8238fd21e9e3", x"a453511686dab86b");
            when 5998706 => data <= (x"9e290a096e6b4ab5", x"e971790abeb66848", x"c7603da90bb6191c", x"325b603be6fb8340", x"d6298f13a834bdc7", x"1604b75381e4c231", x"0f99424eeaab5eca", x"df9699dcb0adcf98");
            when 30207808 => data <= (x"6be866881e884a60", x"480613efb51aa247", x"38f9d4d851432feb", x"8cd4fc3f3dd3e8ad", x"a0dccabe15b83764", x"15626cffacbb2573", x"09c245483a7d4e5a", x"2b9c198b22b3b7e6");
            when 14221835 => data <= (x"25c6be6aa4a83680", x"637359b39688b7c4", x"052d2d4f17f16955", x"090b11e63d3d8223", x"80667a2372fc4eb1", x"bf59953ec36da2e7", x"5186d3d1b68766d7", x"35e4a2298f14de5d");
            when 23559398 => data <= (x"216c4dbbdf8f1972", x"7cf5e1821df02b47", x"6940463e153b32f8", x"54d23f5de21a84a3", x"9beea4b1e82f451d", x"6bff88b37ef707c7", x"369c2ac92eafb321", x"c851abf21f426265");
            when 2927426 => data <= (x"3a42f5015aa259b2", x"7af2b79b1c3898de", x"c9a3a127df57e622", x"abea133705a47d68", x"b93ccdcd67c936d9", x"40f60234b99fac49", x"50ee4b5efca9bbbd", x"8a2f9c458791d641");
            when 12667120 => data <= (x"b188c434ec2e3153", x"50c958decb715ea7", x"490ccc6fe4512c66", x"30dea5922d431af3", x"0f9ba45378a58836", x"b27f975ac06701e1", x"e59b6f12b0727450", x"e7f8043ed7e40d5e");
            when 28781999 => data <= (x"0fcd933f871df96b", x"ee11141854bf7acd", x"be8ba360f8e7bda9", x"f238be5cad671486", x"9821df67eed6d56e", x"5bbdec01d97539c4", x"e94b6c71db849fec", x"7faf934d49e0b6d2");
            when 6651136 => data <= (x"29f2cc9dc1cf72eb", x"f46c9a4c57691aad", x"613a6569d7f5086e", x"075d1c4b02b5352a", x"bfc2e19380404d30", x"405e05c59e84547a", x"798c7a9345488fd7", x"caed83ce8b9b5a77");
            when 7872661 => data <= (x"7a12b5e1dd2300f6", x"f0c5851a37b2ecff", x"294dc36552733bb9", x"a007ced904521512", x"c66c3a324b47e625", x"144dbb848e6ec3fe", x"acadf36ba38016d5", x"75bb29b627fe018c");
            when 18145631 => data <= (x"81877aaef4b2f579", x"7e5a73d04a8db3d7", x"3c7316548bcfead9", x"e3194872a5efc1e3", x"cd99c7cae483b3df", x"c853a2405f9898bb", x"2c535a1b8264e33f", x"6748a198c7dfc826");
            when 11943329 => data <= (x"2551f8c9e3274e21", x"79356f64640afad0", x"463c6f7755fd20d4", x"24ec55846cfdc030", x"b411b375bed1a327", x"13c4d00cdc4aa9a9", x"9ff27c99ebe1cf66", x"6898bb867271c41d");
            when 24836082 => data <= (x"67e01ced947f70cd", x"b66aded60eeb828b", x"cbf745426cd27919", x"356f7076e0bcae4c", x"4beddd6b817817fa", x"a24d30a37b037897", x"8d9e8b2d56416edd", x"ab6486e04ac0c384");
            when 23012451 => data <= (x"a5c4e37172af7aa0", x"ad12fc7334b4e678", x"4ad4ad9c1ea0373a", x"008142d97b1465b1", x"b47961404032fab5", x"f6eae077c7d10561", x"95bf18e7de36ea41", x"2b3a72a3708340fd");
            when 30907129 => data <= (x"e52ccfffdeb6bffb", x"606f1956cc506b22", x"edf0b118f9581341", x"e5b1777c6caa4992", x"d16901c540e78620", x"dcea51da17314d94", x"1320639f130cd800", x"827a1073b52f0335");
            when 14895878 => data <= (x"9efa19120a83d10a", x"e012af582d13ba79", x"6fb08b8fe784c52e", x"5c14c85b998b9ff5", x"9f183b999cea33f8", x"dbe24c5dd8e681b8", x"b79ef220da2a7708", x"eb3e0e29acd9fd5a");
            when 27570149 => data <= (x"0c0e9f6931918695", x"bc7db9cef91b086c", x"b1c27bb29bf76687", x"5eb0dee1869e154b", x"a438f0a928dc1c1e", x"37dba6378d0f38d2", x"f1e07608895d3f77", x"44632e527aa9c3a9");
            when 8859131 => data <= (x"b9674cbc34777694", x"7a988940f793ecdd", x"4e556a39ca9be7e1", x"35b9c466b2c53a33", x"f9971c3e5d227e5a", x"c0d2b8f894d5e61a", x"09190c1de7f97339", x"b61870fd63618c02");
            when 6816383 => data <= (x"4d602a13bb634252", x"dd5a58584f08ab35", x"2da4be6a4da53e27", x"6e71a42274a96541", x"14ce7485c22b96cd", x"95b0474666b51167", x"8e2eb9a1f028daba", x"662b922ea360f355");
            when 8350596 => data <= (x"832e3a4061595c5b", x"312bde66db93cf51", x"4103e122870dd242", x"dd1dc3eed346fbf2", x"d4ee007aeb8957a9", x"a87a5cea1dfdb0bc", x"60f1aeb534bb9cf5", x"eb5cf93998b1772d");
            when 8002759 => data <= (x"0d69550048e81c04", x"ef4cd3189973e797", x"13f78fec9b362cc8", x"d3437691d43f8621", x"798f5e152ef548e8", x"d6df8d56954b2e47", x"d4754cf6fe93f379", x"f946b868387d346d");
            when 31345019 => data <= (x"057e0da981ec758e", x"8c363d72a9946ebb", x"6b08215695e9aa4d", x"f24b06cc9e19b4d6", x"70f99b0286ed0d56", x"0f3084afe3037620", x"676416afdb0e54ad", x"6aff40c59f5ed1fb");
            when 24344238 => data <= (x"282d4aed21d0fd6d", x"0dd4d2d4d52667fb", x"ea6f209c81a47bc5", x"298aa327b7ac83e4", x"ab9219176e0407d9", x"802cbfba42a1b196", x"7fb56264a6573a70", x"255d20bc9e98ce8d");
            when 20455664 => data <= (x"0eb2ca8b972ff8eb", x"d7b1eae6255a3b7a", x"d3e74db5b63503dc", x"fb054063476eed94", x"3a93fea755cf86e0", x"eebf4f2bc10f6b2b", x"58511c63ef52bed5", x"5429132036194465");
            when 27026193 => data <= (x"9629df904dd67204", x"a8b045f0565164ad", x"a757afbe431cec4f", x"93d69eb2ea6b3f14", x"b599ed1dd34d5d0e", x"4844de3b930cd8d0", x"2438347d5cd949eb", x"efbcca74cd147338");
            when 29965878 => data <= (x"1830182cb3b3d4dc", x"a373225a38739b79", x"0b2671037af9dc1c", x"fec63aab7c7d9792", x"c2518e96a4621915", x"23b45124a91143ed", x"1b935a2ba94ad887", x"828daaf029d2a1d9");
            when 22655147 => data <= (x"975e78ecae57e7c6", x"45981f6cae4127ed", x"36bb1b056596edf3", x"1a1ff1144ae03b43", x"20c0507534c63e60", x"df123d166bcda1aa", x"c5ff0372467f37ac", x"baa97a8159fecb0a");
            when 4723502 => data <= (x"4d73a40c654f43a8", x"c0be453626766008", x"197f553ac35e8fcc", x"58fe55e5e1f58bb9", x"e0aac73638e6a44d", x"1bdbbe4eb07ab7bd", x"49bc9e59be87a55c", x"20203ff7b96770f7");
            when 20169046 => data <= (x"eac4b907f2ab1442", x"ad5379aea2c321bf", x"fed0a55b7c67ec91", x"a0f25b68b5d0273b", x"783237817a0f7565", x"06217be819ba1e6c", x"2e28a72251e33924", x"3f1bef7168a75945");
            when 31704067 => data <= (x"9d33de5c08be49f7", x"f7c89e3c5c93a1f8", x"c8a021eb7db59db1", x"b2cb05ba2b0be927", x"27615dd2f12f1a63", x"f7eb43559ef28210", x"f10131df94027d30", x"34d676265de31e67");
            when 7590837 => data <= (x"becf7408e859ee49", x"a48b13f47617d13c", x"cb0fce8a01f5a4f9", x"cc25e45c25be4b7a", x"028d5460e10a5134", x"f54708ac93842d81", x"76ec58b59e30c932", x"57b62c6b44e8a512");
            when 3820474 => data <= (x"7c547bb10ce4ae23", x"5d2512f071e9bf84", x"7c789d4327574de7", x"e75515db21fa0819", x"c3dcdfdcbc9d9b4f", x"ca6f3301b29931f7", x"10b93c37626ed584", x"c7182dc3dbb04cf1");
            when 21028951 => data <= (x"054f5c814b83058a", x"9c4385f10c4447a6", x"4de7f456cabb29f4", x"2cc551d41d906c40", x"8ae13be17ebfe876", x"ffce0e1bca443e30", x"8a1110469250ce79", x"4df682a54950ed6f");
            when 3509627 => data <= (x"ef1b1db74f4249ad", x"5e18325c8ed865cd", x"13ab3e6baf7cb4eb", x"c10ed8c37429fd42", x"0736030fdaf7d3b7", x"64a55ed76e3d6b3c", x"779d239e87b0f28c", x"493f53f6fd7fa8df");
            when 6007133 => data <= (x"56eb2c7cf10efed6", x"8797add822eeeb0f", x"f1c5394378c3f800", x"1bd922a8e4428a20", x"9cb99088057d1f95", x"8848f766a3d93fab", x"d8dfb714404d56d4", x"b3faf539f9176380");
            when 33701420 => data <= (x"a470c9f95e202170", x"45cb7a08d3991dfb", x"fa69c4c0753e1f2b", x"2f3e78f98ba40bb6", x"847f0eb1dd6b56a4", x"a5ad26ff800bb8a0", x"6b06288eaca45427", x"78b5c0c510589d55");
            when 19174237 => data <= (x"58bc6df021c9203b", x"2ce61d869e582c23", x"bad505fa9e9c0742", x"4b9bdee3bbd9f17d", x"96a91739b5ccf133", x"f8426d8a62039e7e", x"76e86c2264da662c", x"0777eb3512726943");
            when 11814141 => data <= (x"f97bd2a2e516a045", x"f95c61a77f111c58", x"88f603b5f08b8236", x"4f327d4233652bb5", x"4258f6965aaa1412", x"42bfb0883eeac587", x"f219bee62ceb93cd", x"197f22ef1bd14e33");
            when 3823736 => data <= (x"d020fa77c27729f5", x"37d8b2ebc87a5a8f", x"5b30e8cae8e2fcde", x"51337cd6c3de8962", x"edfab199e7a10eee", x"5c9a8f9708d349e2", x"3a113e3780747c41", x"5c11515db2f07f4f");
            when 976035 => data <= (x"b298f33fab2f1112", x"da35c2d4d8d337ff", x"6cd190aa742bab20", x"f4d9b6da95e6c99a", x"a79cfb9a1a30dcd3", x"8448be4a70d0a30c", x"d5dd761427561339", x"e597d90272e1323f");
            when 10443658 => data <= (x"7b4d160bae66a458", x"7d9af8f0c3139ea0", x"523431f5f0c56e77", x"5d53c223441c26d6", x"58bed96e213f0c4e", x"5adba7e6c68cf4a7", x"49e29f25fc435961", x"eae9483039dd647b");
            when 18265303 => data <= (x"790771b9786991ca", x"815c516963b767d8", x"1d0cc55fbec6345c", x"2f09a3f30002c505", x"bb38b5eeb85f738c", x"912b2bab800d90c3", x"27d3979bf7d4c6a3", x"4b32b9f1e34a050f");
            when 4315389 => data <= (x"820b1a10a449b872", x"946b6242dc96d65d", x"2dff136e97dd82c8", x"11e4d5bac3b2163f", x"89f6a3283d196aed", x"545462f97b890998", x"36fc3d0ebac9f24f", x"87920794253d4dee");
            when 20232009 => data <= (x"5e1a67935b4ca4b6", x"807ed5be112c15b6", x"43cab1781976e10a", x"9ba699d2c7460d0b", x"8dda134796b3c3aa", x"dbbe6a9a14841600", x"ec051965b51447d2", x"56e2ff38471b19e6");
            when 6292133 => data <= (x"5a30171e9aa92fe3", x"3d338cb535e1ee8f", x"7eb02288fbe88c99", x"d1f156f9a8845ffd", x"9af5b4a8c05e006f", x"eebc66eb600da4b2", x"279c3513bfa51b19", x"683425b6b4b58662");
            when 4768520 => data <= (x"7ea2e2d980883cb1", x"3b5a2515aa9c88ce", x"c586200e28502b14", x"1e8752c8af01805d", x"bea9204effca11b8", x"665b5a681c98b88c", x"9fb277f0239835bd", x"e3321fc6cc2eb049");
            when 27723442 => data <= (x"297c5af98bf4ce6d", x"a8e2188449b17673", x"254f39aee991e29e", x"f90b2524b91feaa1", x"7342f7843440268b", x"dc3c01033281073b", x"be203c004f7014b2", x"54f8499c0c8c534f");
            when 7268635 => data <= (x"5ad246620918584d", x"779b6583f2c365f3", x"78b3b0d90bdd754b", x"78371d5533b9b54f", x"5cf0629202fae323", x"ce7b1cda88a6c0a8", x"604cd76461f92733", x"141718ac220b82ab");
            when 19587281 => data <= (x"7b022e47894c6ceb", x"a156f71b8b35d856", x"9c0596cbb998f11e", x"31033c27335ae57c", x"5bb94b4e214546e9", x"b0b0a720b0fe446d", x"6c66218bed4c7fa9", x"eb96a483d806e867");
            when 11556142 => data <= (x"690c45f4496d0cd6", x"bf562e2b4b72d681", x"f72197a11cfde174", x"bc7431d258bef8b6", x"fbfc567faf3174d7", x"60a2834117ba9ddc", x"4dc2375c27fb43c1", x"b9db2971af9a38e1");
            when 25935426 => data <= (x"0d788b01139efaaf", x"586d25e6d91bb0d4", x"d647ef3732a2c881", x"55c8e43980fa7ae9", x"e243ab5d75e6c6d2", x"ab8d6a0854a2c0bf", x"fa37eeb262f8b6af", x"86096f4d8164a18f");
            when 21173386 => data <= (x"da41823c15ad5eeb", x"a9e8de4a1b51da55", x"9183f9a70d2ffab9", x"e0d3dd242c757490", x"d0173a8a3cea5c07", x"2685dc1f3ad3845c", x"561853c7b798fb01", x"cf49845b01016b15");
            when 6445758 => data <= (x"6a91dd70c24e2428", x"debf2bb18691a3d7", x"d321f1e4bdb05777", x"bafa6c92cbc22b4d", x"da8d47895dddc843", x"ab0d2ae339b442f8", x"1dbed3d1129cb232", x"ed85c006a4b68bb2");
            when 3962679 => data <= (x"92b30561c5e58b78", x"99a6d3675c6dc624", x"236f813eec0855fe", x"00081317a91b47e8", x"297f6c084b2e82e4", x"8811094f8f1c81ff", x"4ba5cfd67aa75988", x"92a20716d413f57c");
            when 33049608 => data <= (x"42bb57f37f1eac02", x"c0406935e0aee7d3", x"761f9bc277ee17bb", x"bd901ad41ccd817a", x"999ef186283c70b0", x"96a44d002677908f", x"e33f8969d9a48da5", x"4d01342b8d9022f7");
            when 21723161 => data <= (x"b1da96a1eeb03c44", x"a2dc17aac42fe721", x"a0dd0571b87eec8d", x"5ce7997c4cbbfd9d", x"fb7c2e32703c60e1", x"f42d88b199ab0db8", x"86ffd795f9d4f7f5", x"639c8d11676ae96e");
            when 26862972 => data <= (x"7c4194b6167cbfbc", x"2292b7b52ccce701", x"aba890b3993a4e9a", x"35e591de4d87960f", x"24278d96fd9fa677", x"4019662bf538d400", x"fac32b1aa28e884b", x"17c0b86412c3561e");
            when 26424414 => data <= (x"a6a96986168ea090", x"abe7c86b67d2fa1a", x"324e8bf1ba6b42eb", x"add9e51502c2f57e", x"934756ba7c5ce672", x"535431e1d604066c", x"bf839e14f04bcfa2", x"dff2c7a0533d0def");
            when 24561097 => data <= (x"0c5b4c3d81f33cf4", x"96ee6b681c62ebcb", x"c6a21f2d10ea31a0", x"91d3db506d22b33f", x"a4980b00b02766ba", x"3ac808269f7ff14e", x"13e5e69fc10a59d3", x"80068cc1474721c1");
            when 2821311 => data <= (x"ea3a81520ab1fb1f", x"3b4c4430171ec250", x"26b8b4c5010667fb", x"9640a9615977a172", x"4e5bfb2390cfaf13", x"7fde7aa40bef61f3", x"42e183bb933cf2f9", x"18b2b5d182860c9d");
            when 6559751 => data <= (x"cb7208cd0b382e7d", x"3d6f7cc75a189e92", x"aab8f8ec22c386ae", x"ff6d6e15fe92795d", x"98b80d02dd546bea", x"a0c0a69ac85957e1", x"aed6f1309dd30f7f", x"01f73dbc68aaa4a3");
            when 25842139 => data <= (x"53aaa32b5ea82f48", x"0702a12f0626827d", x"2aaa8c8810cce91c", x"0195b17e9e057d3f", x"f054e672ea56dc22", x"583c4626bf3fe6e4", x"3809f85b048ca921", x"c2da12b05e2fdfc0");
            when 18695570 => data <= (x"d8cec7a608fa75dd", x"c7bedf3a6cf26eb6", x"a3e9a367748367de", x"f15bb0db1bcdb445", x"5faa57b94eaaecea", x"00e78435cb0edaed", x"855309757f147fc4", x"fbb63520920d09d3");
            when 24099915 => data <= (x"8ffbc629806a0f41", x"06b57469a892aaa9", x"bb9a44f0981f015e", x"d1d7bf2e8e77bbcc", x"cabe3af5db9d1688", x"0aa94e8c9fd34854", x"434dddbad9fb9a24", x"22b314a5243b96a6");
            when 2993166 => data <= (x"2cee24d6573501c9", x"99628638d0689a75", x"6cf7e7e29cb6750c", x"67b848ea92b3b39e", x"e8459978858f8482", x"0b591a53e742018d", x"70a896d6baef2f6b", x"b94d8c42d9753f49");
            when 27145557 => data <= (x"cf560222e5703c89", x"1f2e4695e01d6965", x"2066e54a51e71e0b", x"e8d26f24f4f9bb03", x"558435a29d7adba8", x"07d923c7e1408445", x"965e5c041ddfec0d", x"faa599ae1ca3c660");
            when 5257415 => data <= (x"1a17bdb54a60dc1d", x"e86f3da352e19501", x"afc00c0e3bb0473c", x"417dfeb8e3cf60d0", x"3e65f6252042e507", x"a99e3a436f34815c", x"fd44aced3a3d741d", x"ba2141807f03b32b");
            when 3232144 => data <= (x"4a2f4fe0733d773c", x"a4a6bf0d418862fe", x"311fa48a0db0b5d5", x"8f673597fec83aad", x"7f20308337cfa1e9", x"af1eccd7de59b281", x"51cec1d0809a5f1d", x"22e8d23f3a310b74");
            when 4782364 => data <= (x"f530948a7bfcde71", x"c5f3d6ff67a4e702", x"6f4d73fc6e9429e9", x"20b337ade5e40362", x"b23ea128d850cc09", x"e54b1608105641e9", x"54bd67cfe1ee7a0f", x"5646a997356350f8");
            when 1560103 => data <= (x"f31a3cb78caf8aa0", x"1196493a97de0380", x"c56eb98837086b77", x"a048ed3326c4c999", x"8f4c203c85ec55f5", x"d31f6b68331d440e", x"a54e38fce4d3635b", x"f376aab1b9d0c96b");
            when 22228305 => data <= (x"9532ff2d4d73aece", x"a726d730bbee6015", x"27542b754fe7399d", x"22b318518767deb3", x"97a402a935a5ae4b", x"8bd3164bdbfe69aa", x"bf825f96c4ae9e0a", x"5e743a61385e63cc");
            when 7999093 => data <= (x"849156aec67d3bf1", x"711fca4094ddf209", x"72d0ab11ec686311", x"21de0f5e1deb2d49", x"e11b9937cd1fa1d8", x"321a582d6826b06d", x"668ebfd0938721c8", x"d7bd6f32bcc23ce3");
            when 11880775 => data <= (x"32999a5e76795671", x"a0fd70ebf2e13b38", x"0d3fafb8106926a7", x"acebfbf3cc33ccc0", x"c032d70b6efd816e", x"43978818803c3fb2", x"714ce6e4f26ecb45", x"7c44bf54f811c332");
            when 30377781 => data <= (x"e73505959e839f77", x"671c25cfc6959c7d", x"a1e65fb7c8c94b95", x"fae29992dc904ab6", x"650dc30ccbb61d5b", x"f8fee255a1a89ad1", x"d38a8a2ea5ff10bb", x"54f78fc721bd867b");
            when 33364926 => data <= (x"b5e6657a948838ed", x"efdd9b84ade65f72", x"c107742e3b1dc18b", x"adb9fbf99e8632ea", x"08802ea30909b393", x"b88a3672e8d77c81", x"5a26e117142b0a83", x"c3df3b88e7f1f9fb");
            when 27337129 => data <= (x"d9ca1c6c9bfd49e6", x"1181fb443ea2aafe", x"f9ea606f1457839b", x"eff98ea8bc21708e", x"03585326b13aa2af", x"548569f637257c0a", x"21de8e9d0230363a", x"8843ba8010e6b547");
            when 28618179 => data <= (x"3ec796a535474268", x"c52599133e542b10", x"73f95ec74eef3a61", x"988a2e3a505fd6e6", x"29c68cceab26306e", x"2aa9d9929c6fae4e", x"46492d439a8da4cb", x"0c419e15be6d99d2");
            when 31032435 => data <= (x"6bca793dd7c4bd04", x"61e52cd70bc77754", x"3a7e7bf926f9b1a7", x"52c55f59cff286ea", x"b8b8e45928279868", x"1963963df0cc3ab3", x"3f9bb8720ad426b7", x"54679b9a985d6554");
            when 11002996 => data <= (x"43243f16fde8381e", x"4d6126a5d02aac5d", x"2e94c200128c2d98", x"df4326a108b53113", x"5950f9729074f524", x"764c98ff4876160e", x"a728b7cbfcea8a03", x"37e52f6539300960");
            when 21123002 => data <= (x"0ac170c6e9a9e005", x"efad4ae13e62a763", x"e12251866e4f7f12", x"baae0bf85572e19d", x"f7c4ae80bda7f8f0", x"4da897ae4b760eec", x"feb2a35f5405ea5e", x"b25e1b6f942e837c");
            when 20942369 => data <= (x"17d317ab43a8f613", x"96c20ea89d81ab6d", x"b25616a435ccdeb6", x"18399003d6321b10", x"f7da194d1833b400", x"573226ddb532666b", x"10788a64a4c9851a", x"9e1cee8d75be9578");
            when 26024811 => data <= (x"217776f83aaccf62", x"1c724117c5c3f50d", x"938add20ec8c099b", x"277e3bf49e40a401", x"4d0aeaca67e3db1f", x"933ed72b0c5bff33", x"4d21918ab934cd00", x"dc0513f70e06ebba");
            when 15204307 => data <= (x"b4bc7da71e689713", x"52566b9ef7644d39", x"023128cb4045dc5d", x"be834da490090334", x"d11e9a72cd2bb5ad", x"ea87a1d0e85e3103", x"6f46eb8d2a26f98e", x"5fc6d8c098f88ee4");
            when 15582713 => data <= (x"5a8f4c0f24793c29", x"3b6531f8e5b9be0f", x"65c826cca6ee7568", x"629c25f1c53e4167", x"9ad675de3b9c7914", x"c8e2b18af8a0ea8d", x"089258aa2a8d5b10", x"ee157a25f561cc94");
            when 17178650 => data <= (x"1c7b26ce632dbb49", x"9edd82a2e7c022b8", x"e48f2e78fb7efd52", x"b90129558278c340", x"aa0770eaece3903d", x"9f63bb325b068923", x"2a99c1388495e151", x"32dbc86cae401b40");
            when 5388806 => data <= (x"6a9a6b0a3443aac4", x"7c0fecdd6dc98290", x"94103ef4ff948979", x"584081b992775eca", x"12ca393f6df06ccf", x"76371cf261f25f52", x"d653bceb510db3bd", x"ecfa7580afbd06b4");
            when 7106532 => data <= (x"6f72389874b34183", x"bfeb2acb5109668a", x"cff75ca0c78f294a", x"48e8dad026bbbccb", x"879d0b3e631442d3", x"32b0f39c67bf6e91", x"7a2936b9be9621a8", x"58ecba934fbbe2d1");
            when 21698908 => data <= (x"eaa239d1d296262b", x"9ee91742c28c489a", x"ce21cda8eb245e88", x"d691a3e8df57881e", x"0842c9f5a0196cc7", x"18bcb76259bdf73e", x"35fd9a218ede28de", x"14db0ffea6ac15f4");
            when 6063779 => data <= (x"40990e34a6e81832", x"435b01a80f1066b9", x"25582b0ee2c02274", x"8ba759e15ceadb70", x"68363907832838cc", x"bb429f527112b174", x"8daf8dc9f596c626", x"d9e4c5314abacb09");
            when 8778234 => data <= (x"fe1ec96e4d5d5880", x"6c991dcd68aa3b8d", x"77b5f6fb60030f7c", x"34dfef6225cab8f9", x"9b35bf163840b3ba", x"df670980ce4dc6c3", x"c8fcf1c5a4ad2425", x"5ed00982a395fb02");
            when 10813890 => data <= (x"1eafa1c14bfc96eb", x"fdb0d451ea04b280", x"48416c3fd184c434", x"1fafffbedd5c60c2", x"3ed2f261b97898e9", x"13e724af9b219339", x"0ebcc6da0ad9db30", x"57678b7288f567f6");
            when 1123674 => data <= (x"797079a7441723e3", x"34cb4745a834abcd", x"7ebf31d6562f1f32", x"bd12d271cd3f635c", x"33b2a6f32307f6e1", x"f670f6d051dc1eab", x"b51eef2160b6c22e", x"1091e675e78b1e4e");
            when 8018474 => data <= (x"6f91bbaaf687d82d", x"13ff7d136d068f20", x"9c989814985c885e", x"0aa549e70fb1a17f", x"0c421b42768d2af1", x"5856a0a7a4a9c305", x"cce398bfc7230dc4", x"d195f87a4f762aac");
            when 31718035 => data <= (x"d556e2292fb4f27c", x"e49d6ef6ae6aa6fe", x"76ebb38c8e1252c0", x"4efb6b72ca68937e", x"b13ca9b736d106a7", x"72073a39c6f358bc", x"58c9b751466c1980", x"d97388dad83811d3");
            when 1569661 => data <= (x"6fc865b42e0e0713", x"2fa48723c87503eb", x"24265be987e8c1c4", x"0cf8f3cd39d62317", x"b87920d1dc78b75a", x"5f7965daec1e0b5a", x"1de211fa2a43c441", x"765c93a14ab192f1");
            when 14226436 => data <= (x"dc92a01125e6e87b", x"830ba38efdccf3cf", x"84fe4b0f627d557f", x"dc50cec8c5f7d704", x"344d164c4d80e45a", x"44ba7df2519f49c9", x"f4eb4276ca7632cf", x"032655c1128a80b2");
            when 25063046 => data <= (x"434593eecf432e27", x"bd47e162a9dc11ba", x"0035946408fafdbd", x"ce23e48c0243f077", x"188dede3885bebb7", x"0b1050ccc61c9594", x"d2e9dd938ff6364b", x"8ede2d7f210bb2db");
            when 1344870 => data <= (x"1f024ef70d86902a", x"8f7a7bb96c87c09d", x"6d1619393c88fd80", x"4bf66cabfa3c6706", x"9a31817f2010862c", x"8b8bccac52f6ba67", x"58a3c99c887200a6", x"47a9da3917aada7e");
            when 10445380 => data <= (x"a4e30677b2068a2f", x"bd1c03e6f1b9f288", x"e522a9cb1674b237", x"0aecea6e5254bc69", x"f08841e6c9ec589b", x"76dc8da84744d79e", x"b7323fd81c954c71", x"a24d31b580f243c8");
            when 23632532 => data <= (x"8e832457c531c12b", x"769e8f34b85e8d1a", x"e01115aa4bc443d7", x"dc26c17e9ff9102f", x"3c8c5a83b5557d23", x"a1c96dc835676b87", x"4cc82bc2032ee4e3", x"ccadb31524bc558d");
            when 33511200 => data <= (x"c56281f12c2f9136", x"787328837f92e35f", x"e13cda5663e7962f", x"adcd6d00d1afd1fb", x"b5052523602cd5d3", x"6f74d091c3b8faad", x"1be7881619638aac", x"7684caf262724ad6");
            when 19682672 => data <= (x"0b8706810a62658d", x"84e05a8b1167e22d", x"0fb3df80a5f8c759", x"c398d6ff439b0005", x"3bcdf7f9b01bf105", x"3cd0fe64194e8a04", x"a23e791f4d7f8fc8", x"61152bdb93fcb893");
            when 10817017 => data <= (x"3a3c8337b644ff3d", x"bd2687964e00a546", x"da11889c4a9d502c", x"348cc5130914d163", x"2a772a220939626f", x"ca037e6c5017bc49", x"d62367a251cacd60", x"6d05f0206695af0f");
            when 30767408 => data <= (x"4cafaf34573fa98a", x"2f691998f47ac179", x"d609aa8d68a574b6", x"144817d92e9104bc", x"89f3a8184a9c476d", x"ce076236ff762ae3", x"8b80f615f9ef0b62", x"1e6dfe7c4fb04884");
            when 28722234 => data <= (x"9b410b1d30a5f26a", x"76ce228acbb6fe36", x"91b2aca5b8ae6dfe", x"10f95879a3b23ead", x"ad44a69f8c05353c", x"0b815f8fdab854d4", x"ac19c954d923ca77", x"9d33720cf9150ae2");
            when 1572620 => data <= (x"481c87912cf4268e", x"e79d4f70bdfed39f", x"4c543aeffbdc1091", x"db1707775a7c943e", x"d296f3a2f00e0339", x"5699ec353125a42a", x"85a8c1552d2862f1", x"d1485826f685acb7");
            when 13077924 => data <= (x"afe82a0a8adbc350", x"0b4909c1ccbd3f1d", x"b50f499eeb67fe44", x"f95992723a051fa8", x"4457c64e4ce7f0fb", x"d403378efaf2ac88", x"13233c2c924eeaf7", x"d16e25cd02e87447");
            when 11181090 => data <= (x"386d899fbc518ab2", x"53d73f3872b543b9", x"551b7e5e9258c0f1", x"a858d354c223cef6", x"d4118a3a5a858199", x"20673ef291793e9a", x"f535c3594c3859eb", x"bd5caef686d73795");
            when 33727815 => data <= (x"b06d829b50dbfb34", x"88d5c2724d1adfb9", x"282b7c352a6773c7", x"365aecbc8bc21d4f", x"06f69016ccb6294b", x"7a5894ea5a57049b", x"336c5ec65300a3ae", x"d5fbef1fef6c15fb");
            when 32053200 => data <= (x"0f358ead00ed2899", x"46730f734ec25c1b", x"3721bbc4c2d18a5a", x"c8bdf6b3b2ab8f4f", x"ceaddf9bd2c1cd6a", x"80c3258a3aa34f95", x"65afe7a58bd88bb2", x"d0c8649bc18a5cd6");
            when 9092891 => data <= (x"81aff971550e36f9", x"410484447f924639", x"2b14884676d25849", x"140fe658e5555d10", x"381737971d3d3b7c", x"36629d5fa952dd95", x"44e93cff1d90bc93", x"735dc2aa367be64b");
            when 8886272 => data <= (x"494b00e22ceb64d7", x"9bc85604dc520dff", x"c649adb231d6d3eb", x"dbb838892843a4a0", x"170e5c66c4bfad53", x"d51011b7a51bb17b", x"4168e49031473c32", x"16593b897b552a98");
            when 24949265 => data <= (x"96e71f2cd7282746", x"6e45af6b0c61d7ea", x"406718d222cb2069", x"8ec44d921f10654f", x"ba717c02c5f6e291", x"227f67c3d4ebd0ab", x"b5219ed784a10df0", x"c3f99ac48bd604fd");
            when 3621801 => data <= (x"8dde1faa0127890b", x"8c96a47ddfe719c5", x"0f94205723507260", x"8f6ea6811c1cf548", x"a011cd20beabd532", x"db4fa1dea98be028", x"322fb7243979a85f", x"14b3d5c18368e412");
            when 19966192 => data <= (x"1ac9066d49d3b099", x"020428300f19d963", x"9c6894a0a5f47a12", x"87b3316994f7f9e8", x"66290b01b10faa2b", x"effed227c14d0987", x"efe77acbbc5f177d", x"3125bb966dee7c40");
            when 9820164 => data <= (x"a605c10c167889d3", x"4997006f0a9d3dc7", x"00ba2b99867146a9", x"83b6b76e84583d4c", x"13a16d1d951823ca", x"03cb573a64877a3d", x"5f8fd1f2406f6ba6", x"95da051a6d62a9c2");
            when 19377473 => data <= (x"7afa09e9390cd60f", x"46be60d3b259687e", x"b16435a73f14e811", x"04a64ab2afbef082", x"133193d601108970", x"eb237ffb7f68f80a", x"8c12bed71ff1c37d", x"b2164cdb5a031f3c");
            when 1560284 => data <= (x"5245cd56103e6da7", x"5fe20cf76f5b9aaf", x"2ecf798a09a42fe9", x"c74233cebeecf0c1", x"94340917e4e45ede", x"21328d89f7a78f8d", x"5f24c1dd0e372aa1", x"006a4553e5980585");
            when 8508027 => data <= (x"180f0da57e05ed79", x"8f99fcd81263e9c4", x"dfa892103c542668", x"31ab21b93fa21a31", x"0b0d0a10ba148e89", x"775e3674f7e9352b", x"bad3bb1da73600b6", x"d55043851a494beb");
            when 12700533 => data <= (x"5348049523a2351e", x"b0c725f169f2a990", x"b762c380cf2af839", x"67e161ad2b5f5573", x"583406e0cd49b5ac", x"fa0341b15aea1ed0", x"5e52d05a0ab93587", x"e7b2b7a801b06397");
            when 5809884 => data <= (x"72360082c8b685d5", x"276660430e141c42", x"258e2cf61428f505", x"4d8d566526b56d41", x"cf64159d35c72784", x"dcd8e57ff9a65c04", x"0e782dde1330c471", x"8ff7cecaee443892");
            when 19942627 => data <= (x"559c0fb39cdf67e2", x"aff0e71d39c8350a", x"7ec676d0aa61fbd5", x"9c73ad0e601c665b", x"d3c907211b30a243", x"ed9b6735160e26a2", x"3c57d0c98db158bc", x"f2208b96b9a93bf7");
            when 3112236 => data <= (x"4c1e51461a5549a3", x"b4a60dbe6de04c49", x"15300fc26bd20333", x"131a78898ad217b2", x"87cdccb0eeb8af70", x"8f5f47c33c27a575", x"f30b2b28fc7fe301", x"996c8b1a70f8c288");
            when 25365922 => data <= (x"35d7dbd160f60c84", x"5facb0959dfec86a", x"574badb1784445fb", x"07a0c24922e4d430", x"2409ded30eabfa24", x"4813499fb5b3052d", x"5b3993f045be7bc4", x"e61f45b52580ea35");
            when 13084631 => data <= (x"724030e805acaec7", x"3adc0520610a6ddb", x"8b757342200abe4d", x"a57f1029d05713d8", x"cfc0519dd60ce411", x"b302024a42cbe65b", x"19b5a0e7698e8341", x"f880a5b1f478eac8");
            when 8212370 => data <= (x"65daf8bb46b9da8a", x"08e19f5cf235418c", x"2b4a6de078d0e4ef", x"31fd2321192d7571", x"5a539c96c3380f67", x"471e7dee55e1d000", x"f3e0039cfeb22dab", x"c73e4f575c10f9ee");
            when 28196118 => data <= (x"a2c64ff76bfa6271", x"3c58b5e20d168212", x"2b9208a8a6c74763", x"9e81706f8b307490", x"cda618d5587a68d6", x"e4557ee0a27b8f7e", x"2f7bc058df96312b", x"9e0a17c30b997e42");
            when 4735111 => data <= (x"ec9efe5971ba0132", x"38f2529c3b64f344", x"4c3a2a08babbd576", x"0dd53412951e08a6", x"b27135812cd97613", x"79f5b874485ffa13", x"14f02210c1923170", x"706750f482fbf6cd");
            when 29997748 => data <= (x"d6cc3f0dab175b44", x"aae6684556a572dd", x"df450c1e5eeb3ee9", x"5db0128893f5fb1e", x"788d0f54ac039804", x"60a42f1765a2259a", x"f3b084a7b7874a84", x"054a089ce411dea2");
            when 22873917 => data <= (x"afc4762c14d09175", x"7abeaaccb4c6ec3e", x"4e2e7c81759e79f1", x"b962d3d6161afafa", x"87c0fb3a69f31a26", x"1348959c8061f3fe", x"43e30d7c11b381f8", x"77aad91420c933b2");
            when 23675657 => data <= (x"bf613d5a7e746242", x"af8b2b3097c93336", x"3a4a9c397ec1b451", x"db253e8221cf7298", x"e54bbb20efa74613", x"63f622db1550ab58", x"da65a11c1ef28d8d", x"468d0c80ecfa1ffa");
            when 16816692 => data <= (x"d9366e9034f82606", x"a26a6125374ef7f0", x"f8de466f6fc81f27", x"1037beb1e5521806", x"8eba43931db26892", x"568277e9af24c636", x"a07af92dc61e527c", x"b1e7e13e690ab3f8");
            when 24252161 => data <= (x"5e406bd2471d2622", x"27c221d40ac5c472", x"f5bc30e5720de539", x"a99d0c3741b8909d", x"94879a73db8ee5c8", x"09857d9b4403bc40", x"aabd02b7b956b0a0", x"06522590bf633761");
            when 5591028 => data <= (x"bcdafa21cc59d18a", x"a9871d2685b86170", x"57f273afaf149857", x"d6c2d829bc7ced19", x"68e73e41fa7002a5", x"187f5a0ab5372584", x"fe8c62982707dcb2", x"27ce3eff5736852a");
            when 4016222 => data <= (x"b7aded0706930959", x"d2e88f308c87b63b", x"6427577eeaf51d51", x"e46ff458d5206a0c", x"d8675168249cd68d", x"1e400a7b992a2cdb", x"6fe1ef086be0952c", x"cfbc704335b049ca");
            when 4703042 => data <= (x"49f06cd4d1a05355", x"9341c857d71c3992", x"c017cafc97546137", x"252b883d9e1b506a", x"68d1f1de8d4fa1e3", x"c4cc7d476b0dee08", x"0259ee9c5ee9b300", x"c311784eb7b82d0f");
            when 33329131 => data <= (x"ce27be9cc3a102a9", x"66d862f49bc7856e", x"b7b2ddfc28b031a1", x"f189a51d81dc764b", x"6be1be0cd1254330", x"dc0d1054f96caa05", x"cf9a8d164a9379fe", x"245a9c25e73fc38e");
            when 10559094 => data <= (x"01768f1f16877811", x"baf9c0936105b0db", x"4356720810f912d5", x"e7fea86e883c1ee2", x"737d1dd2ac8caa8e", x"1a634eb0cd096e9a", x"d412732604105d08", x"9625a20833ee5fad");
            when 20381050 => data <= (x"7753a1ff19066c7e", x"dcb222566bfcc2c0", x"143c12ea8b52aed0", x"39d453fbd9fab25f", x"38768fffeec4a05e", x"19f270cc0091f063", x"54f51ad6a73a28ff", x"9ee393d08fff1d8a");
            when 6874247 => data <= (x"99381c9a65e41110", x"61a06315f34efcc0", x"651eb26e08cf6214", x"a92bfaf3e98cdc33", x"57e478cac67ff3b0", x"d5469bf980f58050", x"4c57e7832971b7cf", x"a36daf02669c0791");
            when 15668390 => data <= (x"deacc0435bb39a34", x"4f9aeea9c46b490f", x"36b7a43ca393e392", x"5abe015438854069", x"9271ed8e5c0e61a4", x"503404044f94397d", x"008a7d1a5808bbfc", x"860b6548f149f702");
            when 16107536 => data <= (x"25f10016b76a5d28", x"2f675a9e67dbaeac", x"97acecf4ba55ca1b", x"192e46fd4522e751", x"497dd4651c34d5d6", x"a10ba4a817f4616b", x"240358f7370bebb5", x"9280759f2015a535");
            when 33173791 => data <= (x"d0cd92f699fe32ef", x"f5d93c172c774c24", x"fdae8c8e639a6d11", x"390c9be2bd6e8266", x"cfcfd4972e411f39", x"ed4b190d960de861", x"143b8292e86ded77", x"0baf85a741e76088");
            when 18679295 => data <= (x"85903669899fa9dd", x"2b50df73ea54e019", x"202eb5f41487ba06", x"e7236fb8765ed8a0", x"59b96c5913f26dc2", x"3fc478d510263f98", x"68f91d0fab6862a8", x"67c89dd622ffce02");
            when 19837595 => data <= (x"7e5d2671487862ae", x"1b1fc4f583435825", x"ab0a38c949d31a0b", x"a95cb5ab42867ed6", x"eb31cfc08ad6ed25", x"de499881d0396375", x"b8dd4d2acaf7fa45", x"c07e4219626d64a5");
            when 25597990 => data <= (x"01d6909dbbd05fe2", x"7ed96a55680f5764", x"737144a43cf3c6f5", x"8869ee997fd7c916", x"10783cf21a47bdab", x"9fa26a03c71e0ecc", x"c1655fa155dbc594", x"51c8b6d1c351b412");
            when 765705 => data <= (x"6470e83beb834e2d", x"f84351bb0314c3df", x"fae191e7a5af0a88", x"a24e89b6b4f756be", x"c3094acc85cf32a0", x"1864d39f5dee91ff", x"c58b9ec2432b7ab8", x"071b0178f0321d30");
            when 22581830 => data <= (x"5c4d814149b7d099", x"c2a5c2264bc350c0", x"2d12b0cdbfdef720", x"7592663b0d3e7836", x"0d8b9f2e2a9a665d", x"d04d905df65c190b", x"8c761a682dc8d5ec", x"524296a799a6de50");
            when 21468085 => data <= (x"3f11d749ef9acbe2", x"1d834bf986c6fd08", x"4f524fd269760a04", x"8450626778f2376e", x"8abec72010e4958b", x"623155acf128afff", x"22ae740984a29351", x"aef1383007ff8b93");
            when 33865287 => data <= (x"52acfa9330325f84", x"c500d8c682486055", x"01323f4326cca016", x"951e4dbe2a992550", x"7c318804e1822470", x"f92296a56d93f31c", x"4c8826e3aa14066a", x"f32798a10d4eca59");
            when 32407188 => data <= (x"631be4b1f423f336", x"9a8b194eb93bda77", x"649a99b990379e46", x"9566b1a53a80468a", x"8e382c55c87e8a0e", x"16c0bf7a47844e32", x"7b1e3368a4fb40e8", x"f3667ea5b1778ea9");
            when 25495010 => data <= (x"9bce222b20b6b440", x"bc767e931e009877", x"3e61722196e5792e", x"13f7817fa333e9da", x"f77cbbacd7faa87f", x"ffbdeeafe038e14c", x"d6ee68ca1ca733df", x"57d8b4f46ec02b28");
            when 6264019 => data <= (x"14e3fc6fd5572405", x"4b43c30653973bc0", x"c87ec6d7a2eb9149", x"5be4d240ab8883d7", x"775dfbc3e2848b71", x"84bf1f9a9935aeb1", x"91b5a8f99bcb88ca", x"1d67e255b5778066");
            when 20283311 => data <= (x"b3da00a4bb98b145", x"6ba3480c1512ce6e", x"69fa9884b4e15fe5", x"0107c20b0ae7bff5", x"5e683be16b3da2a7", x"db0f995f599bcbe1", x"44c0ff49e5e5e0a9", x"0280532209417bfd");
            when 6091966 => data <= (x"071112560f58ecec", x"26cc5a84874898c3", x"d68ab43d807cf1a6", x"47f3be3029eb4060", x"0462653f3d781232", x"1b77bd59c039013c", x"4b805ced9d0f5585", x"a0b10a0584af8ec3");
            when 28595206 => data <= (x"630914a27cc27c19", x"1324ba4481998db4", x"20f74ca102afe3c2", x"9d4f010e51f5c70e", x"f50153f17c17a080", x"6c472419f03eb464", x"e7a65023c697e66c", x"e699e77aef5b1460");
            when 23687961 => data <= (x"e93f1fd0c9e042da", x"c7aef67c11361744", x"31b5b7833b6dcba3", x"365751afae276db8", x"8205e4e8317b214e", x"ead94791663024b9", x"ac964d639311783f", x"f01838ceca4b2efa");
            when 29604028 => data <= (x"baa12362839d140e", x"0d16cb31c077f907", x"d96e2e49ca7e4b71", x"80b500827c024225", x"ba49757de4e42b4b", x"fe83480d5d81b5ad", x"f1f52091c25b995a", x"28418f3553f23233");
            when 12885810 => data <= (x"a91007cce0620d2f", x"2aa1ac7752774ceb", x"8278593557c58554", x"44e666acef52795a", x"279d09a83248a37e", x"343b65272a05938b", x"2cc4458728330beb", x"a4dc5ccaaf83e9d9");
            when 23107261 => data <= (x"8636cc95be225cc0", x"15212a1222559a8b", x"c2a1c2d31f0657f7", x"78d442b98b01079a", x"284278cabc176e84", x"9b7c7c654b1cb83c", x"6f8ec95175ad857e", x"86de3d0f7990e704");
            when 12870976 => data <= (x"5fad81fc855a37d1", x"4a84c6ab8b7affa6", x"22004dea246c2abb", x"5c33f4406f9eac2a", x"41aec3b4c0f11907", x"bb5d6d1ff0196e3b", x"b0e7c641133ec67e", x"f8af2d7dcd110cc5");
            when 26945202 => data <= (x"5ba52cd6e7919b72", x"f22ab0554f36792f", x"14de6c4e613f58e9", x"1fd86bbb77bce7fa", x"7c0c3910a5eb8a27", x"6be94701ce2f6226", x"ec9bde0d2e1feb62", x"8947d98402ef2bfb");
            when 14013849 => data <= (x"010dfd9c1f696788", x"6c221b703654e562", x"99d3e6fe127e10e8", x"4c2f15fc42ebf1a3", x"bccbc0c3b9dd220b", x"7d2f5753201e161b", x"c41916b6f9fbc262", x"620d5a7e08a7c12d");
            when 2598320 => data <= (x"aa288ebe9c8be151", x"d30947fab46d1e41", x"0bbed92ffa4837c5", x"26e8cfd68ad71bb1", x"f0ff9f7b91cdea2f", x"cb90e4f315cb0a48", x"19509a1db745a57a", x"bca8b9d67e259097");
            when 20807524 => data <= (x"dac6b43e9d70417a", x"6da289b8a6116a68", x"b9578cf90e2e3682", x"a02493b4cf1c5b75", x"067bd15154312cdd", x"22e250ede181c065", x"74221bc708082dc2", x"66f478c751583d4f");
            when 16151925 => data <= (x"e79533bc8b92421c", x"44b8f7017443ac4a", x"5c03d0afcf1dc158", x"d2024a647fd383d5", x"672427f99dea567f", x"dc39a6390fe0795a", x"153e417d38f1d58d", x"f1617845d3454f39");
            when 33576173 => data <= (x"432a7bce1e680274", x"9167fb648a164e2c", x"e4f9a9963d91ba87", x"79c6abbf587d18b6", x"5c0e84e4915bd14f", x"03dca8afa473ff70", x"c06a1f9fc23547be", x"42116a0d3205abef");
            when 3243800 => data <= (x"37304521836c7da6", x"167389d99c49351c", x"39fe14b267de0e1f", x"bc66689768f14c2b", x"88818b60c055b121", x"9f723d3ee2a7bf87", x"40438df6cf576952", x"6217ed6cd987c3d6");
            when 24218441 => data <= (x"833d3ac20d6afd43", x"faefc8e319d6cd36", x"41abfda7dc198bc9", x"f921bcae6e1518e2", x"44aead14ed60a2d9", x"7fd3008f94e90f85", x"6429624568afd53b", x"95abef50eb2ca292");
            when 11844984 => data <= (x"b9f5cc659bb224c5", x"ca764dc0f88b03b8", x"2697d8abb5d11db1", x"c1fa15fc7e29c9db", x"39e1d5becfbfd84b", x"65cf3671f51ac64d", x"87e8c6273f9b684d", x"af9bdc2b3bccb80b");
            when 26060517 => data <= (x"f5420b944b3fa0df", x"82af2adc236efb12", x"9e85143bfd9b63ec", x"da97354b220314e3", x"5400763309787a09", x"8a867cd77757d122", x"3bf20e74975b6c5b", x"7351ef0d59f07595");
            when 18729905 => data <= (x"8c9811fc9fd4ac99", x"eb7f167ecb772eaa", x"b0f1047003fbef74", x"ece74e19ada6f9c6", x"33513b0b52f66642", x"5661373bdaf8d871", x"b216822b3657ff81", x"9aa797919330b0d6");
            when 3930209 => data <= (x"7342c5f97bf04e0a", x"526925a7f26ede86", x"df14d1a2f5917371", x"504396848e19cbd1", x"8cfe9bb2f8622ab3", x"4e2c15b7562be9aa", x"44c927a12d0204c6", x"f9bee7edbc88c1a7");
            when 19678915 => data <= (x"accdf1fb234a1738", x"54ee8c0d3e9444df", x"fe61aaf678ebdd7c", x"6f30b16739a7e8d0", x"8b379bbfa286557e", x"56476a770823426b", x"7e02895105d614dd", x"130aa22c010f0f05");
            when 20712945 => data <= (x"f04bab98536c60c2", x"ca4c8cccc75e5ac7", x"dc4b9c57fd31c25f", x"f96e2a3225ce84e5", x"0e86d72dd22b8d5e", x"63628d67f2815527", x"287c18735ac38e1c", x"39b699a753cb40a2");
            when 18789966 => data <= (x"9b283a0ad3f599f3", x"954fb6165e427674", x"e2be38ce7ad175ee", x"f41ed27ada3f21fa", x"a0db89052c139f5e", x"c308e3775924de24", x"19b0d49c7494cda4", x"ef85e8028c17cab7");
            when 20377207 => data <= (x"8f61e76db806b342", x"0f5d20228fd2082d", x"747b07b68559de38", x"abbc373059a30236", x"720d79d9da50bf71", x"c08fbd62009ef74f", x"534b9589dc365e3b", x"21e556aca3a17f7e");
            when 25330359 => data <= (x"e5fcb96160dabc69", x"628500feefd649c7", x"4695b26293a7707d", x"216819037d1bdb2a", x"db80db99b7f7ce68", x"9f01cb002153ba85", x"1f3ca6526ea5d196", x"357ffdb40e78f0a8");
            when 7128361 => data <= (x"e95a8a61b060e7a3", x"221d1ffc7036a481", x"30905fae90f6a706", x"c2dda15d3cc7d6b7", x"f7c1e12c7737e800", x"84d6666078de7378", x"9331a73fecb0007f", x"9399f08d83890996");
            when 31943587 => data <= (x"d47730cfbcfdf260", x"c370cf527318eab8", x"0514264c0ddbac4a", x"b7b32e645ebfbb04", x"49e443cbe1eed3e2", x"de606a431491fe3b", x"ffd8fb9d53535941", x"2bcd7d9579cae3ab");
            when 3787143 => data <= (x"d7f941873291879c", x"38057d6a49c2eb4e", x"6ef2f83afd1d32bb", x"cef1e35fe67a745a", x"bf2eadca8b9c5513", x"ecb8f90aa5c223c0", x"a00b11821b6a19a5", x"39ccf8205f8770ea");
            when 1085295 => data <= (x"3af0bba6e03e7a03", x"b3dc52e9a447acf9", x"183145a213a5fb85", x"1ad9705ae980035f", x"b2bbccde015e7faf", x"2b2ac1087a688e33", x"8f29ba826c3ec87d", x"204fc3d81eaddf8e");
            when 9286154 => data <= (x"013d258f4e436adf", x"8608dccec955cc84", x"4b7f70d8b3cd5757", x"50b60e2c9aa22d7d", x"69b9b259f7df5beb", x"76ad141380b26806", x"73abc5cb974f9186", x"519a1e3eaa3d6b72");
            when 23364859 => data <= (x"2775ea63ccb67c25", x"bbed0b92f9d34f3f", x"405776d908d7a432", x"077c715a7b3ef46c", x"5c49524629d52636", x"a9a967556e81b88a", x"f7c09c751f67710f", x"b928a46f5d5b6b8a");
            when 20287658 => data <= (x"1591b63110ed184e", x"eb71e312715bd48d", x"e146fc7276f57829", x"37e3d4707c8c222a", x"ebfbdf1ec3ca4e7b", x"c6a7b5dab75bbdf8", x"0ea5ef748c346e07", x"aa592bd786e0781d");
            when 20481823 => data <= (x"f578281667f3ee6c", x"675ead2ae1baee8a", x"7bf9e016ba72f0ba", x"9ebcd94d2557efc7", x"dbf168cd2a8c7217", x"071e662a5f6def7f", x"7960320e9f4836fa", x"9be80e5f4dfe2e4c");
            when 3063420 => data <= (x"4fb44385934ef9f0", x"9904ab04370f9813", x"ab19e8a22a2a767a", x"9da7b047eded6721", x"3ede7b6542d14862", x"767198a107360e25", x"67b7f77bf384d8ca", x"fec136dbd90c3177");
            when 30768621 => data <= (x"4c520e515cf66c55", x"a9211afb544297aa", x"bf58ebd56b7dbbab", x"7938335aeb6d58b9", x"80bb7f56390738d4", x"cf557133443e1c5f", x"deffd129ac3c202e", x"f9d0535d60aa38f9");
            when 26232864 => data <= (x"37ad63fd00dd7bbc", x"a4561cf4e2287cc5", x"1651d9c2dc7fb377", x"88f9850a0a429451", x"f97e4642c7b92df2", x"8e125f451388b0d9", x"68f6ba423b755418", x"536e1b06cfcedfab");
            when 13817603 => data <= (x"e6c38bb84284f488", x"8e4440a5ee680364", x"b261ca93a9bc6b12", x"bd85104b29043762", x"ff5b5c42ba86fc11", x"db2a4a883f9fb211", x"a727d063ded16d72", x"852b643e38eff94b");
            when 4503908 => data <= (x"2eb3af07483ba82c", x"68f2d6cc352d5b9f", x"a6a90957a6f6743d", x"c4fa274f62e7e44d", x"4d1fcc7d2c9ff5ff", x"8fd05ad94ca6c42c", x"3b3c8666d17de46b", x"63eed4e9a4eb6582");
            when 13751681 => data <= (x"8bc67bda2883c738", x"d0218187d4135396", x"780ee3d434617442", x"aac3f122459d9bd9", x"1cd671aeddcecdda", x"d390c99c73aa5085", x"859dec70c58e401b", x"da65e6f99dbc2766");
            when 15903420 => data <= (x"06cabad7f53c9537", x"df54e2a83bd505d3", x"1a6078814e188f20", x"ae34f4f8c7ecdbb1", x"29cc7f039c9bc4cc", x"acff3105c71c522a", x"76fd2513b2f1ad42", x"3fd98f797b979bf2");
            when 2993154 => data <= (x"711e5fcdd8959d54", x"cadbeece0a1f9dc1", x"94fbd8822109020e", x"b400cb97d731bf9c", x"a1764c9b5578702b", x"d89cd2b615d552ee", x"407fb9dfc8d8fecb", x"f364389cd3c0cc76");
            when 9149475 => data <= (x"d3d4a49fca36b979", x"87f8d1b4e9e367a9", x"13fe48bfa131c14a", x"2d39ac87e25df82c", x"49dd080bf6a382b3", x"15e1faf10359e147", x"0ad2a7565fd1f51e", x"555a04066c3f9a38");
            when 32346792 => data <= (x"707c8ee8ce7299d2", x"7e4550582cbc1f90", x"100942ddfb12d80f", x"141b52ce88ee0576", x"b2f06d9207732b00", x"87e57d7d08473e19", x"45750766a2cfa436", x"dfb0036dc9dfe134");
            when 24275215 => data <= (x"0ae3b73c1b4754ae", x"1b1349d3c73f16e9", x"2725d32a032cfc86", x"37868f8865074526", x"62d6c2bbb1a6e7b0", x"ab8fcb54982cb6d7", x"800347d0c2a3907d", x"ef6c70626dab093c");
            when 4430761 => data <= (x"9d21ca2f2925d849", x"c19697512a0a6b3b", x"5d247d59ce545cea", x"6612f3d2a1c77bdd", x"0e64dc43772cdccd", x"210e6acc38c6c4cd", x"32fc2cf49ad759af", x"fb21e14b145a478a");
            when 11762732 => data <= (x"140e7245e12b3c99", x"34e41de4cd1d8da6", x"0e9594b3d6f42569", x"52b955e1874fc646", x"c9a456780417ad40", x"df22620fc8a26ca3", x"47d1267579d8a714", x"921b51b5bab3c33c");
            when 18984800 => data <= (x"ff8a7e0019a4842d", x"d43daaa82955af77", x"ca2668e5e6aac948", x"e0dae94c919acdcf", x"f11359b0c1f6eb38", x"d3927e24aac254d1", x"e2aaadc9da211983", x"0685e65283fdebb1");
            when 21282792 => data <= (x"fb73fc7b8dbd6611", x"ffe0b66d320a89c4", x"37c6e76bf9359b33", x"ee6e3f4ebb21be24", x"50587e4e090f7d2a", x"d09cd75cbf4e216b", x"012224e91845a2ce", x"a6ec7091ce88e7d4");
            when 16617056 => data <= (x"00f2ad0f58d87f71", x"1e9584cdd53dc0fb", x"d2415f4b10102693", x"1ed1d00967313456", x"27b6dd0cf8f402ad", x"d6da978cb8fa3364", x"2e852e02bde95bb3", x"c2706856ad6ff0df");
            when 15612877 => data <= (x"7708f919d963426f", x"2acb8403304b08ca", x"b412c6b38b1f6df7", x"3c14abbe7661e445", x"9f74c8ca822e8bdf", x"e53b8f0d3443b912", x"c1c049e713af50cc", x"0d0be277842515e7");
            when 8383848 => data <= (x"583c71c43f0ce61e", x"ca715517966369ca", x"29f30a18628edfe6", x"e1056556a97563bf", x"480e564d50975d9d", x"6c9b2da9f15fd732", x"e691e896cd20e40b", x"e57f6f1a8d916a33");
            when 12355187 => data <= (x"e8c05ddb2992e48a", x"5b99f12bd235f15b", x"8f9896b0f9d9180d", x"5f00597b486bc9e3", x"73210b6d8489d640", x"ba96b34d49c16ac7", x"49b51db001ac7e4c", x"3c848367a0a92600");
            when 33377282 => data <= (x"9a97ae3c5ec0ee76", x"47d84710ea5bcfa9", x"022831d5af950459", x"66f2d48ad21ff7e4", x"336a45ed0d558f94", x"c98812be7c328fce", x"4cee726cb9124a86", x"58ce06d5228e2aed");
            when 3131265 => data <= (x"37d617f811ed6a17", x"c74a9f8165f104ec", x"3758fdd749bc1f52", x"b2ff900a841909cc", x"b86d64f8487d766a", x"b8870ea426c6babe", x"ef4ca878f3a74646", x"21de6c089e03861d");
            when 10106375 => data <= (x"80568d4158e16178", x"37ae68b0cc960106", x"87b42ebe2881e878", x"ff4a8ba27c946f83", x"2717b301207a762c", x"39b27a2bb314e4ef", x"4d937d636b8ece8e", x"4168c2666d928bd1");
            when 1148787 => data <= (x"3d6dd59b3ba5ece0", x"bf9ef7b5f68bf0ec", x"6a37139e3a27bad3", x"6e6a1544be290aca", x"2a81ca6c4578be85", x"5bbe14c10a0daf9e", x"603d842f3c37b6ba", x"5459f9588c448ef8");
            when 31106638 => data <= (x"76321b632a7f3091", x"4d23cf460e1c93b2", x"207dd4e240a5da07", x"e37f76173bd227c5", x"def38c3919b60b5b", x"4caeddf3795a3de7", x"2e66510e8355cf97", x"e1e8f1e4133941f9");
            when 27125390 => data <= (x"43b4181ce7f86ae7", x"f59d0c4142b4ee12", x"1c1913d0b69fb899", x"8e1c457a99f23dd1", x"6c77a282708a5a05", x"7d695e7121e9c5da", x"e7668e3f28129466", x"a6e7ea4a8677a393");
            when 28851768 => data <= (x"5a6e2130cf076f81", x"416de5b33f6429ec", x"a46fb5cfa3fdca42", x"3982931784af8926", x"70afb9868344975a", x"00121f49fb0e3e27", x"0337d390273c3e49", x"3fe52d71be907b34");
            when 19069225 => data <= (x"010cbcd3d267fd61", x"95858890e02fc79f", x"48ed0a665d5ba317", x"78d280e5a829b3ed", x"ca2d652fbf0f7b98", x"1b9f4ae12f2be619", x"2fdea8ef5c099bc7", x"d533848160ea51f9");
            when 23545822 => data <= (x"847089ae5d493961", x"be0b9d93075206a7", x"91d807296e4a637f", x"1ac7acc9afadec20", x"6aaa8be7c16e445e", x"2423120dcb75bd46", x"8b3fc64d010668c6", x"669b492be293ad11");
            when 15704419 => data <= (x"0221597e49f94922", x"81e84778849fee49", x"44244a55b1a56738", x"8b5adcaa8b22505e", x"0f8ec329949fc624", x"12823905fe80507c", x"a337c6f6a7636881", x"85a9bb8c3952c8cd");
            when 13532335 => data <= (x"9803ad8607706ce2", x"bb6fc1bd991b245c", x"749c182992a3f866", x"04db5d5952b823ea", x"6dac2d1471a016a1", x"1b7e9857e71aba67", x"29e36a10c40c6dbd", x"b6547ccf54f13542");
            when 6090259 => data <= (x"58d3541aa52db0a0", x"82a24d92c7e972d0", x"063c2796c8d513a5", x"5daa63ba1b7bb17b", x"fccb792b1652f685", x"94914feaf6ac0702", x"589d688ec25554bc", x"476e81822cee3286");
            when 21966062 => data <= (x"980278997b77fdf0", x"8972c3632b3dd95f", x"58770cc7976ac11f", x"ea5b4110b5c426f2", x"7dfbbb02ad6ab54d", x"565b3aa762f25d08", x"59c0bd4ae7411073", x"b1186702ad5fe53a");
            when 26030143 => data <= (x"98d064bf5d29f503", x"67914c88f4a87381", x"077bccbdca93b929", x"667adbe078a2a049", x"63ae6bcf4b6c6da6", x"8713944b3f753362", x"6526175d204acf8e", x"a9d6eefd25e0a03e");
            when 22070791 => data <= (x"6050913a8f1da6ff", x"208470e1fd1e4440", x"df35609dc1b1fabc", x"2a11b14f58115ac6", x"40b3bd4615175075", x"6c10c9a624d3eb97", x"9bc68c6ffd6debc3", x"b43dfe143c548a64");
            when 15062450 => data <= (x"e238b9affca726ba", x"374aac7ce718c2ab", x"441bbcf569960c1e", x"98bd48d36ee3a9c4", x"0749d589de429baa", x"d2dcddb95aa45353", x"bd9c5db958e80086", x"72a4294606ea5cf1");
            when 23689312 => data <= (x"f6168927d67d7cee", x"93c076d48dd97c69", x"4ab80696b54461c8", x"7760e9de72f16071", x"8c605b4024cadcb9", x"5d3fa7f9f02015ce", x"0813f6b5ec69fdbc", x"47dbe17d116234f0");
            when 7056474 => data <= (x"af713483f4d1f7cb", x"eadbb99b12ce8142", x"83a739b9519114c3", x"a7d604cbb74c7696", x"d6407523034cd1c7", x"c83a5d1ff1a53cb0", x"e5881970bf1fc9bc", x"2b79a1f0a7867c06");
            when 3357277 => data <= (x"f296f4b0b1d4b422", x"5c278feb82942753", x"37f6fa1ac114d9f8", x"d75ff9e1309b1c58", x"8bd5beee29363427", x"1c1bfcdb96024a7c", x"512d3af8f62ebcc0", x"dc8b37148b130a27");
            when 27433332 => data <= (x"3e0c058e0eebdd8c", x"ec868bea106eacc3", x"01cfd184d8f85f2f", x"dfa50fe6f13472d7", x"4f9408bc6da8a044", x"0967d4ab3a3f31c7", x"0e6e98fbbb706c72", x"0261bd9df7257d70");
            when 12552745 => data <= (x"9255023484d1388a", x"0953189b7d828082", x"d0dd0186f0eb2423", x"dedd41c342d56b0a", x"1b391b405058e3d0", x"8ee43952a32452b8", x"6cc2ec9b36c8fce2", x"4827188033872193");
            when 1871684 => data <= (x"9bf053695a7d450b", x"590de331752b5a26", x"2740d8da9cdd1d85", x"cafc8cd9faa826a1", x"f9611cb155cfc4ce", x"63f2d1953b15a1cc", x"4d8dbf79f06ab9b8", x"16399644daa86d75");
            when 30601442 => data <= (x"df6a079dfa049914", x"8a2b9eb7060b7f46", x"3f786cdda2639aed", x"59109389670f705e", x"41b0e266dafd4418", x"8af66e25b6353926", x"3364508df1efd3f6", x"4bce8942843d2ef9");
            when 2021944 => data <= (x"eca18796792c698a", x"1fad10167db1f75e", x"9fc651f9784f02be", x"18984b885d70da8f", x"fd6bd335bf569777", x"fa86efc625cf949d", x"6824f3776783ba09", x"510ffbfaad82a601");
            when 5321171 => data <= (x"531c903398504f45", x"f0444b2d797cbb7a", x"b5d5e12bda744080", x"0f024a376033126c", x"5896297dd5fec8ca", x"606ed52eff95a8dc", x"1291982dc3b6fffd", x"7e92a6253dcc07ec");
            when 7045043 => data <= (x"cc62f3b21c59dac5", x"6ef39427da13bd22", x"18820d9f1cdad9ed", x"bad5505b5eef934a", x"8147fa1985c96f6d", x"27326efb449dedb0", x"61e6b0e9e419d3e2", x"c5126cc9b5848b92");
            when 26370589 => data <= (x"ad8d341f6fea554b", x"0dcdafd1f3fb360b", x"430812bc8ffdf170", x"a24724acdb221819", x"8daa7b6a02a9ba89", x"56b3a1aa230e88cf", x"1387cfa3b479aefa", x"69514a5c788494a2");
            when 11398819 => data <= (x"c39a2bc7ab9fa171", x"c205496cfd0128ed", x"e0f77129cab36980", x"300d23440106afcf", x"873f6d41d61da40c", x"c1bee1d9ec129fab", x"24bc8a31df41a53e", x"911a79fca7502430");
            when 8547786 => data <= (x"0e9fe8d7410484c4", x"8627d387e7753923", x"8ae1144ee414c854", x"8cae1c64e4a901fb", x"f95f76c63c0c8d09", x"030c7b1135520784", x"3dfcd7da67e4a70e", x"b89909113efff28c");
            when 5165091 => data <= (x"b0b015852518f9d4", x"692e385f3e0c38e2", x"3e264106c516ffc7", x"9d6216a18f0049ae", x"13e6867a1581374c", x"bddffb429c67f228", x"2f33671addc279e2", x"d66dccd1d65cebee");
            when 27090308 => data <= (x"c12f3b0eb2679fc7", x"4453f295b8da2e18", x"5e88759eae4923ef", x"1e34d72c383456de", x"4d6876b888504f1d", x"db575c3f793f2b9d", x"632602e6b11d352b", x"b0c97f9e6acf8b47");
            when 6087768 => data <= (x"84c1e13cf7d060b6", x"d0cc1a36f48f69b9", x"9b4106686491d9d1", x"3ea24e114d81fc6e", x"d834128cafa10541", x"c76b6f992462e823", x"42f9635c8b4b4ea4", x"c48470144c474d53");
            when 2848017 => data <= (x"773ca3d3d1c58257", x"8ef77259bd25eb3a", x"c986af2687c15a38", x"c556493867f8c27e", x"6ac366793aa3bc58", x"982d2a0c73ddeff2", x"3e01aa8f9c078008", x"c117500943df5135");
            when 6309356 => data <= (x"ed3cc8e2fe7a3b7d", x"216043ff7423e5f0", x"321328d05a8964e1", x"a080f7f1ffbf8c34", x"ae4b19935ca5d4e4", x"9ef735b3289c5604", x"bb6bcdda3e9b89ae", x"8c235e1af975f3a0");
            when 3175886 => data <= (x"8e5d772b764bab67", x"103b55c9e909bb53", x"21249f73489e14f8", x"db7a316bf84c2900", x"636ddb7832cfe13e", x"5a173bdf265da9e7", x"164a7d5303c9d619", x"5c95ef10e508a060");
            when 20952075 => data <= (x"b3e5fde80c0d3b90", x"48c4d76f04bc8e35", x"4d663d677f6a09b4", x"818d23edb0b25e1a", x"d3d8ff5515a051b7", x"2c15e12dca3a7abd", x"c2f34aa012e581e6", x"2adfe078e2052f03");
            when 31050879 => data <= (x"4c4b89fdcb6819f6", x"300b12178fe8b57e", x"97e6e2f8f45ce32e", x"9ee944dac76b1c7d", x"23df9cf84ab4a0c4", x"02d904278d80dca2", x"ea7e6fd4b9b32be7", x"cfbb12e440b42358");
            when 33255021 => data <= (x"2603e26dcc930517", x"87d28a5777eb166f", x"b0a052457f8811f6", x"e277687766ab7b0d", x"e07995b097aa8149", x"ab738494f54ef5e1", x"892c001a70a689e9", x"fa7f7f8afac5d38d");
            when 6264111 => data <= (x"d23f2871899ffed6", x"9fd6bbd3e91242d3", x"7553006e98a1a759", x"accdf8759460aee6", x"19f25e14f0c1d0e7", x"6e44695a4e8518db", x"44fdf8841b38c928", x"9fe63c97ae14ab89");
            when 6880027 => data <= (x"1059a62a64dc0d0a", x"04a8782cbf61fb92", x"b78664320974b09b", x"c8f217af94a81d53", x"f91f431061c20955", x"67c1c1e9f58ae1a1", x"46f06cdf7ecc0c6d", x"3965ac5e7b3283f5");
            when 19420328 => data <= (x"b593eaea7e75d7da", x"b316c14c59835e9b", x"23ce822d86772a47", x"03742576428d8ca1", x"793588f2b87eeb50", x"a71e2fa140f68baf", x"4130f0deda2d9f4e", x"8926fe74b3e01144");
            when 3506994 => data <= (x"379849ccc4fb4264", x"fcf723c027ec4dac", x"712066ba89dbb359", x"6778b1d8e22e55e2", x"7d4c404f8e4f93df", x"adc70908df44acfd", x"8377b04510bee26a", x"a221d90a95ea595d");
            when 11108614 => data <= (x"0f216d2f7acde7e0", x"9384d33ec6fad41b", x"3d3960d092aabd3c", x"d0c8d76cac5f9b00", x"46761f25198d3ab4", x"f65063e7d14b28c9", x"bcebba560f5dab09", x"cff682582149dcb3");
            when 29138048 => data <= (x"b29fa69f34c65050", x"e5bd4de1759638ef", x"b88d624453ba1b26", x"5ef989559488c90c", x"7fc9c5c67ac2848a", x"09e42351642311e3", x"d38e00d634c523a2", x"5e0cffc5649071a7");
            when 21149206 => data <= (x"8022a59357849a98", x"71ed97b0b0d3b099", x"f6b35b3cd4b226f3", x"722edfc2e2349bb9", x"2f1dd88929fa5ef7", x"028a435c1704648d", x"7d05fc21976721cb", x"881406ce835ada1a");
            when 8717329 => data <= (x"430a01099201ade1", x"694594010990d1ce", x"b46b28130ca34b59", x"3772562e3030e37f", x"1b61adcb838241a7", x"4d50cf9d4c89b77b", x"e1e98c6e40dc4f3e", x"59885dde6bd73c47");
            when 30371742 => data <= (x"ada8932028fc5732", x"53261fc8d066dbda", x"3b9ed233941d872a", x"96389e19b58ec562", x"8d7056f256a017dc", x"f5703bef23365bb0", x"33940c36913d18ea", x"085f520b157dcdec");
            when 32802405 => data <= (x"4739ac88d994b6e9", x"f7f2ac6254eda7e5", x"9a5acc209fa7e6c6", x"e1d2d66b5516e29e", x"f2416c22159c7053", x"b3df02b7cee7ee08", x"193c82b2fc67c614", x"2fa8ade4d75a2c99");
            when 28393675 => data <= (x"348eb74c9e39caf4", x"d8967b51422f9d72", x"06757dabd76618b1", x"eac47e5d4a8d8bd6", x"e0cf1f84bce5d010", x"f889cfa2033cd054", x"cf4cc8b4603766b0", x"c2c5edf6e37523bf");
            when 16064351 => data <= (x"dc158d83a76f43a1", x"b0606d617c833578", x"4f2eb26440f9e20f", x"3f3e7e4be0f05f98", x"dff5c5880ba6edac", x"82768f4c6c77bd9d", x"25e85c31cfce4ee8", x"546f265dbf1eea13");
            when 26333132 => data <= (x"6408257974da20e7", x"e260fb352862f5e2", x"d7d84829a1b40ff9", x"378637c4898f1fcc", x"442dd2e7a3bdb7ee", x"dd9b3a948518ca44", x"be2f3b59db60604a", x"0568d1ce8118d0be");
            when 14303173 => data <= (x"932cf90a5174032a", x"d9c6fadcc56dd372", x"75cf343c95ee2fd8", x"26aa8389fd5dbbbe", x"66bc99e69af937af", x"ebcdfac392ffde30", x"a38d3bccf78f740f", x"6e325280efd504c4");
            when 20124513 => data <= (x"e26bae7698393bc4", x"da1adbc11eddd616", x"c59ba9b0b07716ee", x"b9d4bbbd722cd36b", x"c2a5c985543798dd", x"01e0091bf5d7857c", x"14474be3f0a37b74", x"bcd424b21dace0c1");
            when 7598238 => data <= (x"66b6f9677ea65f06", x"b0ea847db7138e13", x"21e39071b28d3641", x"e464cdc7e1e6996a", x"0d554edac3796427", x"f323de712482d587", x"37792dfb2a440041", x"1a8f5ea1bb098713");
            when 8990558 => data <= (x"5e62e8e02814a61f", x"0a18401efc7e5395", x"c130e33eb70e9489", x"ebd72d35336b25ff", x"f0cdbf95862ef338", x"5a46f717ae46d3fc", x"dc2aa31e971328c3", x"458aead1a866a7ff");
            when 27122539 => data <= (x"4acdafbe3147ec4c", x"57df876ab304201b", x"125d2ca8aca81d4c", x"94618d47911c0c79", x"821c7dacbc571a3a", x"8fd26ba957e4c5f5", x"43f2f7197d2c8411", x"67d15da367abc318");
            when 25889557 => data <= (x"53916425c5f4aff7", x"32f606024c4a87ff", x"428679993f4920db", x"898688fc2df58c7d", x"e6150adff301be1a", x"ffbf5b0754d15269", x"66e5018a2aaae43b", x"ec74c6519e9b5871");
            when 32424676 => data <= (x"42cabf92e87caeb9", x"bda06ff67f73ef69", x"721d9ad44f3f1c09", x"9f9b257e2cb91ace", x"f12d068f692d05ce", x"89d52aa7618fe141", x"ca5cf84a8ee4bc64", x"40248c19ee772eba");
            when 29737589 => data <= (x"244200b7cb6c18aa", x"069a472f477c1691", x"f26ccdb785a945ae", x"a7870466e46ad42b", x"e68c7a54146ebbcc", x"00bba2a59f16a358", x"65e75dfe568d16ab", x"cf8fc5f8a0c7b0da");
            when 27497218 => data <= (x"ce5a0fec86cb76f1", x"c0dc9a8d41307377", x"7ec719bb45bc99c3", x"6d34862f512a4a5a", x"23a8fb7de058ee5a", x"f9269788aebb5efd", x"cc31a7d6193bdd8c", x"47bea7236f8dd8f2");
            when 13050423 => data <= (x"8eef38e9bb61b65c", x"68bd64e9ac925da5", x"eee5837885575f7b", x"bd35180971d95144", x"e118fdbf84383d4a", x"8058245de8eb9b23", x"aa87e8d34a733c55", x"02fff05010a7dd86");
            when 1308109 => data <= (x"ce4a39f28dc54cdc", x"d61b72e5a71301ec", x"dba8ec6b9eceee64", x"771b5b5dfbc35164", x"e73978bddfa9bdcf", x"fc4d409c5eb88963", x"f03778a3428cbfd8", x"30514097257b04fa");
            when 10765273 => data <= (x"579f3cb906c7cda8", x"6ddce345ccab1f97", x"01eb792ff9314562", x"4ad18e0be28662d3", x"13f96149e5a52727", x"f63806c26b491f30", x"ef1a19b4337efb8d", x"6daa6e1d4000930e");
            when 12315309 => data <= (x"5740e0b2b87b7e49", x"153a41df04316a85", x"b3d56023297db45d", x"89d15833c42743e6", x"d94fe464c52a5f8f", x"3dd8520591bab063", x"5e0a015c302a5236", x"47ee2b3bf3fd7362");
            when 3988289 => data <= (x"39dfe1602c2e373c", x"8cc4aa0fa3ab6d0c", x"e41275f0ee9d3111", x"1f354cd63f59c5aa", x"7f728116d1bdf3d5", x"f39aa2e9d7df7b75", x"26e1264c3d2c5079", x"7fc6426b4e899e3c");
            when 12858520 => data <= (x"309582be87f0f700", x"cc2614243bd034a2", x"f9dc80fafe733f16", x"3590d950a3892f99", x"857dab4acf091426", x"4d0f8ea296178eaa", x"59c64f21e0ce0b27", x"7ace88a61873e8c5");
            when 25961019 => data <= (x"5119be7be5cb3195", x"e88144e776cdd115", x"587859af38295364", x"f16f547d711a365a", x"de7ff4244f4f35a6", x"57409c4263b51523", x"134c7e86ebfd5c6e", x"415bc4dc36840f4b");
            when 4847018 => data <= (x"8524a1eb4c93622f", x"085bf77dc591ce4c", x"52d2e680b35a3733", x"4860dc153baeaaa8", x"d32bde43e2b2284d", x"3d1454c379b48399", x"5d6a2d65eb9044c3", x"04f4ca8df89156b0");
            when 33366800 => data <= (x"eacba99e2b81a0cd", x"bbe497ff82b5bc76", x"044c1854ab621daf", x"612c5247f12cf2a8", x"2ca9480971e2ea4a", x"4228fff5fba2abfa", x"474d638636338445", x"fa715a2906646ecb");
            when 14501844 => data <= (x"c3c695be4cfdcfc6", x"fa5b0cc2df5df3ad", x"40b1c571109c4ee6", x"94f557d183771f4f", x"030550dda389e380", x"a690ee471ef321c2", x"b7db1c71ab36d6e3", x"a1027b6f303f410a");
            when 27758092 => data <= (x"d16761096f86ec0c", x"2a65350b78946b2d", x"9d43400097ff1b36", x"c0f1aceeb38d4dc0", x"460ecfeaef66e1e1", x"a59b51f819a2f1b6", x"71071526287e0e8a", x"738ad5e8b8a8eceb");
            when 11233873 => data <= (x"6f6ed2a1ed813fe8", x"6a64b0d139012755", x"7760af3e3f8986fc", x"cc956ecb27759f95", x"4527aad031878b08", x"980f616564a69b19", x"29a9fc1d9a6f07bc", x"ba84c463910f5256");
            when 28740808 => data <= (x"f85993e6cd52426e", x"30b3fa984b854242", x"f2a8f3acfab99d32", x"e7867443a7d87cd0", x"1330bf5a5b229745", x"65cbcbab4c470dca", x"6804650559d84e51", x"3f58dbf8927f5bdb");
            when 28553820 => data <= (x"2d70b65e222294b2", x"22bea27e0bbb5ac1", x"8ecd02ab946f4d9e", x"ea7c4e61565f6ed5", x"570856798914ee7e", x"45a30de1d3d55de2", x"a3260ac022b58002", x"b63c2a5f69e859fa");
            when 5111985 => data <= (x"f44f66ac5be10957", x"f78eb607d2a8f3b0", x"65cac5be9713b9ee", x"016e9398eb052489", x"d175ecbba7730ade", x"3197f5c535b24994", x"7cd08c9f90c863b0", x"f25647781334bae4");
            when 33918795 => data <= (x"2bf6a8dc15f33add", x"67191859457cfd9c", x"1942929f87cd8b7d", x"08eeef901031f503", x"f99776a5038004cf", x"4ef5d8c446be74cc", x"929b5ea8108e6f14", x"6f06ff2bfaf17c0d");
            when 22833947 => data <= (x"300543f81cc1d705", x"83c243dbdd173bdc", x"7e1eaaa68707dfdd", x"dbfad41a914b5378", x"6d48c7cf54f55606", x"fcb7c798f14c9250", x"9a390ad6f2943915", x"d556e80ae7182151");
            when 6276937 => data <= (x"5f20fe3c1f74aa55", x"c8c2e50b9ac6d7d0", x"900bfafbade0551e", x"79846e762eeef216", x"ee9d260a630d68b3", x"633cc16eeec2a169", x"a252f635b7578347", x"6e2e3b3228ea06f5");
            when 11980327 => data <= (x"8d3407020a25b708", x"21fff3aa0a732a4a", x"bce07a6bb92a2ab3", x"4edaf4430304583a", x"0624da94709b7bec", x"6e8ae03ad943671b", x"2ef2180716ee97b7", x"4deddc12c4927654");
            when 17328551 => data <= (x"2f5f8d54b1258c7d", x"c697efec5929a35c", x"ba99bd24563c1b60", x"fb612c0668437a91", x"df92f33339b51d22", x"2b7ad13c2008c726", x"b99103a1821d1d35", x"9a0dc27e4e96aafd");
            when 27418029 => data <= (x"2780cd4658499193", x"fac811adb0e2c156", x"29e11f0543147462", x"98dee78a7b4c4099", x"083a737dc6709961", x"3b52d7969b594cdb", x"517105a6fec0a67a", x"ceb2c91d982fd37b");
            when 30166253 => data <= (x"76c1dec806776b90", x"a99055c5cc830248", x"78495432f92b03d0", x"fe1cd2055f26897d", x"333553c2fb3556f6", x"6a7b188c4515b9df", x"d515f0d7c3adc631", x"cb149a0eb102cc8c");
            when 10454177 => data <= (x"048fe65aececc06c", x"c7d089d8cc51f345", x"9209a7a006084af9", x"dc5002907ba75f9d", x"5231b2db624d6adc", x"7a3712a254068118", x"51acd00c4db81996", x"3292e4c12cecb691");
            when 32008871 => data <= (x"878633310d3a5d0e", x"d7e576c9ed52e046", x"eda87f918ce44961", x"9f5efc063a68ddb1", x"ddd2175ebe9e19f9", x"d4c5de659d7b4645", x"91202c7875e8051a", x"57d602ae83899244");
            when 14742252 => data <= (x"c8bee9b3f1bb367e", x"bbd04c18362ae17e", x"c1626bf66b4934ae", x"b67c3ff65bc29adf", x"b6c408d93d896d67", x"972068a3ca837324", x"702684ac17cf429b", x"7b23dafa66152fc8");
            when 29734139 => data <= (x"c2e50779e05447d1", x"b0c47a144c82a85e", x"406afef0fb19a5d1", x"2dc36b10606bcfb1", x"6f3fc9c7e4fc0868", x"f0fb99892fcf6d9e", x"5514375e8c35a8e0", x"5a7f27d97b7c4094");
            when 11236501 => data <= (x"70b29fe5d8f93a37", x"deea89597bbd0e94", x"3cf538bf50f28043", x"0d99d0eda34e92aa", x"99a71c1039884167", x"26872db5bb0b9ad4", x"fd1309408f97779a", x"ba564d7a84a928db");
            when 17028127 => data <= (x"bedfdaa10aa2bafb", x"63ba423989c631bc", x"6f966ea34c0ba837", x"c8540f76a7c06176", x"59edbcbfc922a656", x"db3fb6abd0c1469b", x"ab29a30b160351a5", x"0b4898d863ab80d3");
            when 9180034 => data <= (x"a43fe2ccf27b60cd", x"1fe689b8dff5168e", x"7f796bfb2e791c5c", x"f31900d50a26790c", x"f189eaae6f072262", x"ea180bc856d4aac8", x"aaa92524f1c24645", x"967fd3f3bfc7bb19");
            when 32697467 => data <= (x"ae843e57bb81f047", x"72cf4f8f3eb60fd7", x"0e3f4ea90fa8627a", x"214584d16d6875c5", x"01f8780d9b100dc5", x"50b056f3d7cb6b72", x"bff21384846075d5", x"ccf3819d4187d1f5");
            when 6597488 => data <= (x"0c690a00ad674a71", x"1afbb449b9125af3", x"8d042ae2650d3be2", x"a54a94865ce5e580", x"e2642087d1eb0e3a", x"aeb727bc52f79e7d", x"43aab23027e5df35", x"085713c347f687f5");
            when 19496915 => data <= (x"a0fd4c4007c0f3d2", x"768d1e902d1e058d", x"eac76d4f2936ade8", x"c600edc0a73229b4", x"64518758d658616b", x"a6dd70a1872b7fd2", x"04d99b1b0c3d2575", x"2f317129e269aac2");
            when 824881 => data <= (x"f16c6ef246926f46", x"bc4cd73f43a9d637", x"2da1fc44a354ade4", x"46731ccbb7163a87", x"9fb63812126ae275", x"5d9de7298a5a13d0", x"f84c0b1ef3638cd8", x"25075b8a28fdcf37");
            when 16895587 => data <= (x"b21ecf7cd0a3c4b0", x"eb891be8fe9a52aa", x"5f79f662afa7ef9a", x"dfb0ed0b167a4d60", x"b109d55d06b7943b", x"6a8580ffaed6064a", x"d63f3ad58ce609d3", x"42ae62549db5b319");
            when 577080 => data <= (x"51bfaa39ce5adde9", x"5adfd4e73799ed9e", x"aadc0312e5ab15e4", x"1bd70674bc6433ce", x"f73c5d7092caba38", x"7ec3fd1d29b5599e", x"102413c7becc2d4c", x"c8ba8a5f35e0d570");
            when 9645822 => data <= (x"abd9b76acd67b94a", x"067bb8a9bd2464dc", x"e95b1aefbbf86f4e", x"3643f8521eb2ee16", x"9409b12b10b016af", x"b20a33c1e0ddf00d", x"7273e6a5fb4e58c0", x"08cc37a412e838af");
            when 1528341 => data <= (x"bdbf9c4a5393af66", x"fb984b242e2f6d1a", x"48b2566e6293c2a7", x"99110a6962d5ce26", x"87b4b4b765fdf904", x"93f29486e21c0325", x"21a02c43756eca65", x"0eb48b10c016dcbb");
            when 6099330 => data <= (x"983ab3a0fe2d9e5f", x"52859d6a4244c3e6", x"8a3cef2ee55b7302", x"bed2051ba1afd8f7", x"b5ba27be97706014", x"2584a6960d82d667", x"26c1c01120c60a4e", x"91f5baacc5f26660");
            when 33295516 => data <= (x"66b4c960ceea3c98", x"5004b1e47784d8d2", x"6092a8b3e83b3e0c", x"0dd6bf4980132b9f", x"6f6448d244e457ef", x"e0fecd705dfcdb1b", x"dc85d180fde02d26", x"c3f4623443f2cecc");
            when 21291453 => data <= (x"9b1d35135f799281", x"709deea7b70e10f4", x"69eded3bbd892a86", x"4e81dd4de9dad24b", x"d3d7cb130199e7f0", x"5e490cf57c6e9747", x"feda3a4b574228ad", x"e9a6cc71b9879a97");
            when 543051 => data <= (x"6d60c6ec4c2749be", x"239bd93a4cdcd720", x"a493031a47ceffcc", x"aadfde42930c75b2", x"1b24326fff034afd", x"2dfb285205e776c4", x"ac5a5f68349c1bd2", x"0ae7691c2a2066e6");
            when 3943837 => data <= (x"04d7a0be7510e68e", x"dd53c556f0d07d70", x"ac790632941a5935", x"8ecb5c3ab35bd541", x"7f035ec6b3bd4c52", x"b64c0e011d46cc05", x"408db1b628b20f48", x"8e0fa43bffe91374");
            when 33793778 => data <= (x"8bdc90c60f094009", x"232e7b946d343c1d", x"1c767dc4cfdabaeb", x"561f8c58e4a668ae", x"e0e3837fe0c6ad64", x"3efe3ee8c46ac9de", x"2bb681e9b8e5bb92", x"2456d8de75754dc4");
            when 31915882 => data <= (x"590336cb70f5d425", x"fbf234c09fbb650d", x"f67965dfc57303bb", x"9d4c27651a053d06", x"f5e927af6baf5075", x"5fab9969ecdd41e2", x"482d759e9c761651", x"29411060b19732e5");
            when 21315735 => data <= (x"edd558ba8b94164e", x"b027e152ff9ab9ba", x"e9a47c5bd5493fae", x"9bc7a2ad3b10a73c", x"4507a9a09b07d8ce", x"1089e6314ac624ac", x"31f0d96b17b6c090", x"7eb64012914468a2");
            when 7496538 => data <= (x"235c672594753444", x"47c146138aebddb5", x"987009c7fafc277b", x"f697fe3a0f99456b", x"51b7f52e7a602a89", x"8ebe854635bde0bb", x"1e058800c4368fee", x"2b55fa609cf9801e");
            when 9322650 => data <= (x"286b13c18ba76eb5", x"485190cd0cdaa86f", x"6c4ab2e5fc0b9281", x"d8353ad973462409", x"9fcc0f2b85007ce4", x"927d7fb8d1524b53", x"78942fb432f15bc6", x"0208ad6c7eef0e5f");
            when 4930740 => data <= (x"b932eef42a64e1f6", x"99cec71cf68557c7", x"17b9eb015049f7bc", x"534d71e67363150c", x"a680ba03e5090664", x"e3a122eafeb54f15", x"08a427cab69e0a32", x"5c5aafa21759ed0e");
            when 14649331 => data <= (x"ebba47233e29bc3f", x"59006f4c17859662", x"6ecae84fea2a12c4", x"de908b621714feb3", x"7713e6a75c35e632", x"5a929a33c9f7f4c0", x"6a8a61e0a5380588", x"310ce44c74cac97d");
            when 9408121 => data <= (x"993c84b2e343c515", x"07a7137874e51362", x"1f85d1e98f134bb1", x"b38d7ee92b2e44dd", x"1638c4a97da342a6", x"41a996065c3507b0", x"56c67ef45d81789c", x"800ebbf3d6e817b5");
            when 10078691 => data <= (x"d2b9d7dc8c88e913", x"d67c5013ac91c961", x"143f8e9e0e9afb00", x"14bcdfc83ad7ea41", x"44311536d8546cf9", x"af5b2c064078423c", x"876f1c9c42426386", x"f728716d275f5f4e");
            when 4098896 => data <= (x"c919225191608325", x"ac10784a132c09b9", x"3d2c1469b84a2e4c", x"8ac150bd152e4dfd", x"248a530637d4dc98", x"8b0fdee4a978bf1a", x"835a7ecbdfcba467", x"465f070cdd5fc14b");
            when 3304152 => data <= (x"82e310766df4aa9f", x"4a7cd4b3d43a2811", x"3d0eeadcf4014586", x"a878f0d09d5e81e7", x"22172547115659da", x"0dea0e9121a22eb2", x"bcd822887fbc4508", x"3cb439d0b2e6ed3c");
            when 19165978 => data <= (x"00a3e727cb232468", x"ceefc3c0caf6fdf4", x"685c49ec392f82db", x"1295cdab1f57146d", x"36eb85ae9177a30f", x"a8a22e38bbcdce47", x"76d75725cf3e36e4", x"6f92d724eeb4734c");
            when 27343270 => data <= (x"98f0bc3f9dfe8a97", x"c5995cf09f92dd1c", x"f70d7937bea441ce", x"112c3b001e3472ab", x"ef06202e4a55dfc2", x"e5b7ec6bf2881bf8", x"0b7fed58ff1e38a2", x"ea02a594c088f8e7");
            when 5163788 => data <= (x"dfeff5430ccb212e", x"17a183621cbad812", x"61a881dd225a0526", x"3f9c7c52c3835a26", x"f42d4c7d0cb2c029", x"caa32ba12e459fe4", x"5204d9841649755a", x"729908b7ce3c3dde");
            when 19870876 => data <= (x"5844b831f2d00b93", x"cc66db26cf27ff45", x"7c5eeaae3ba11975", x"b409b69cd53ba213", x"f24273dc5718eedc", x"0095c90e862dc88c", x"97d1f398a11d8ef2", x"a04f69b94bc2d3ae");
            when 15434791 => data <= (x"fa20e08e8c6bc40d", x"f3a8d2016048f5b9", x"6a7f338cd79cebae", x"5bf84bd4bc5e4cf8", x"12ad1307859af67d", x"cc869823a0875709", x"d6a94a05fedb20ce", x"a39bbf5fbc1ed74d");
            when 13317605 => data <= (x"bf630284b83440a0", x"04daae8abca38f32", x"9ca3ecfbbc9acd9a", x"523b9317ae340deb", x"c378af2a4b23a99f", x"768f3fd38e89e15f", x"4dbc09c793e1d516", x"55928cedf1efc13c");
            when 16724014 => data <= (x"983695f8d354a2ff", x"9f4c2d0d2f5ae073", x"ce93f4e098841545", x"d093dbe4d1f572e3", x"ed964f5fa6717711", x"dbc154c1cc7fb2c1", x"51e85421d53adbae", x"349afc94d18d9bdb");
            when 6063887 => data <= (x"c89576f2618f3f29", x"aee238a0c2127b6f", x"ed738f59199cf82c", x"2b3cd9a96fddf2a8", x"627f6ec311cb91e2", x"f37705ea4f3b8c61", x"9cf3556fd624e23e", x"f4f7cf261469f299");
            when 14942383 => data <= (x"b8110d949e09cdc9", x"5cf98d9ff3536dd0", x"87237eee7e3becb1", x"0146d81a88e6825d", x"12cd9991141cd5dc", x"2d988aff510cd98e", x"d7e5089d7b6b3706", x"66d091bf3205fd37");
            when 19334386 => data <= (x"1771cd3a41dd2525", x"26e697675353c086", x"0aa771b5d666ac15", x"30f5d153de1be7a0", x"5f2792c4b10424ea", x"7ff97f13f241645d", x"f2ee93399ed0c957", x"cec82fce880a3395");
            when 20583617 => data <= (x"ea43b6378162c23f", x"f7637077c4a9d3f2", x"8abe60d2fc10aa7b", x"81e82aa292917c28", x"0b60a6ae1da72253", x"e121a393ca9964b9", x"16a418dac06ca54c", x"5fec5ca52a21715f");
            when 10684455 => data <= (x"1f479019943a64ae", x"bb275dcfa9040a27", x"b69c0ce7af2e8437", x"db9e462e36999822", x"14910ad84f0b8c1e", x"49a33a911425f9a0", x"d8a2d549ed55491f", x"af4cabe16b3e7f4c");
            when 24231314 => data <= (x"6dac8b8df6af78eb", x"75069f00244024e1", x"a8e30a9013672fed", x"6cd4729859661080", x"b867ac9de8f5e360", x"f621b130ddbea3f8", x"4eb238e943d207af", x"97a0d29f04466b73");
            when 15326458 => data <= (x"b6a7abbe877c96ce", x"48e151b44f89f18d", x"3d587be02e5a60b8", x"2d2924d01dbb276c", x"2f6ba1abf4adef70", x"bdcfd87c08445d23", x"e387dd5ec8d00139", x"70bf11d22e8f6407");
            when 11065975 => data <= (x"175e8f950f23bf28", x"6353bca8d3558b88", x"53a1f1a5b46d228b", x"2238cd08914d7c3b", x"12c74aeba625df5e", x"27cc7c0f643bb8d5", x"5c02415d284ef9b8", x"8202a0683fa2e631");
            when 32655456 => data <= (x"de9899ec1a456221", x"f4d29d9a1f1177fa", x"d9edf01fe35ed1e9", x"1762be0539b063a1", x"a386a31977a04efa", x"802961ecde5d84ab", x"2020617ed265f496", x"818339fc92774d5e");
            when 2434013 => data <= (x"74cedcd58353c57e", x"fb519e8d972eb226", x"2f1a8623ac8ae4a9", x"eb02d260ec73c22b", x"94823c3ef56c832c", x"4824ebed2ced1398", x"04350e072fd49984", x"b6fbe5c766a31218");
            when 18052571 => data <= (x"6e08b96952c2efdd", x"321d456a0c872f5d", x"3bb79f69b786ec96", x"80fd891e6b448b4f", x"5914888760f1705b", x"912d3f5229939b2f", x"491947bdd3706b51", x"4f4e7a3edbb0887a");
            when 3753546 => data <= (x"f5c46bd73e31ae91", x"b3abae5041dd4e9c", x"a1dbbb1b20b839b9", x"6d7b7cc6d117ff23", x"f81d7ae2f2adad29", x"d750b75bfa07a428", x"0eee0eef30c95c55", x"41837500b5a5735f");
            when 5661095 => data <= (x"8dd9b7b010210b17", x"66f270fcd814460e", x"6770ffa971ee3749", x"a94552536d4b57da", x"4552122f6d454243", x"c09fad4498e5c1c1", x"0930ab2ce5b81016", x"0e3c36d9220973f0");
            when 4508047 => data <= (x"49b9c2335b4723d2", x"571e8c2cdd67cbaf", x"05f33ab0d801166b", x"03cfcb923ebf982e", x"d772c7f8ab295a9f", x"76a7882d2073058f", x"de4d572b16c79772", x"2d7c49f506c4c747");
            when 4957389 => data <= (x"75111135bc018326", x"5925b4787ec9ae5b", x"0c97f59370896dd4", x"a846a690bec85d4e", x"59240e67ce47ab7f", x"5d1ea1cf18961c98", x"53aea4caed92f6b8", x"36f1b2be94523823");
            when 22611811 => data <= (x"236454f52264ed60", x"acb2b95d37162c12", x"52b68fd516c1ce12", x"f2a19b7bbfd1b84d", x"fe9efdfc7d3670ce", x"959fe76d33073cb1", x"a2ff221e77bd6c51", x"be3abc03afccf08c");
            when 21852436 => data <= (x"6d343e485be85880", x"d6636aa7d1b09997", x"14b75db564c1c794", x"b3821064ea1fdb2b", x"bf4db33914873020", x"035953f47209be37", x"1b95b621d9e0e5b6", x"440ec06df16d8168");
            when 26698395 => data <= (x"1c2b85c1df7d5ab1", x"0a7e06c374404509", x"5371da42365a4958", x"45d16e8acd7af47f", x"4f04e0c374a09d5a", x"2d61567025217494", x"98028e21c5f888b8", x"a54fca025d2f078d");
            when 6625496 => data <= (x"a0aa5745cb56bec0", x"f453b2f7196bd454", x"0f26de058124c47c", x"482f69acf308a4fe", x"c4963611a3cc0245", x"aa7b4ee2ddb077e1", x"08bd4254abee5436", x"72b742c74eca6e12");
            when 24630373 => data <= (x"9368085d175b762a", x"69939653b985b01f", x"0a391ca503772410", x"ef743ef797b3c1b1", x"7597bff34aed8774", x"d75d0f7c4eb38ea3", x"95fa1561230b0ae4", x"c842f44c0d16a497");
            when 17306873 => data <= (x"c659f4829149ceb7", x"72e070780023be2e", x"f512ddfe8bf71f5f", x"ce0c70e0eef300be", x"af70111086b340a4", x"1985f3982755b531", x"494d8c50630778ec", x"1c57880a6544cc72");
            when 7077717 => data <= (x"ae8042e202b313c6", x"aba38f6ee9ccd353", x"15ccf2494cf86270", x"e499698d3574b860", x"59ce4517b8afc006", x"b2060a0f083c0356", x"4b3177ac7821f1a6", x"e4dfeaebe5a014a0");
            when 12619358 => data <= (x"6f054a26dc1e8147", x"38606c51510b44d3", x"f4d6db94c860161b", x"f0e7afe445db42f2", x"a20c98810b16f409", x"7a8dfd9943696c92", x"777ebe41c0ad883f", x"02117fb3499748aa");
            when 23643675 => data <= (x"315f92a988ff5437", x"2c5c2be794e880cf", x"a05e6caf7962b2f7", x"42550848ed378944", x"46f941bc5332051e", x"110c948424319428", x"94e19a80773a3135", x"8b37ec492bebbce3");
            when 15785845 => data <= (x"fa4ad4d1ec48db78", x"1562356a99b58f3b", x"c9787df54265b377", x"7d13c974d14ed279", x"b1f8b7ecb87cbcd0", x"cb55120cc6a94fc9", x"4b13e79cfca619d0", x"5122b15afb5616c7");
            when 26615893 => data <= (x"486ff5b5b25cb313", x"3ff34a06b203277f", x"e041822d6976a5df", x"7bc8915ec78763d9", x"05d9d38ec3b1357b", x"39b787c48448c4a6", x"612c8e24e4c060fb", x"1cfe00dd42b51333");
            when 7797923 => data <= (x"9fc274aef9e2d210", x"edc47aa8aaae154a", x"0bc10925ffb03718", x"73d2572fa31bb750", x"6a1df570fe232bf8", x"7a03e6b0c320049e", x"4b617f6a51b3311b", x"855ac2eed1000132");
            when 18183308 => data <= (x"0f65e7aaa0cf62af", x"d2cb68ed7c94b33e", x"b1cf2368962928ca", x"9458c3026ce1ec25", x"a96451f356f6f486", x"dc7afea13f8474f8", x"39ecee1b64a5458e", x"f8771d0aa3e6f17b");
            when 22192446 => data <= (x"a0ffa57251469837", x"93a0bc03674f6399", x"2454272c09b62804", x"df3506370a2af973", x"d297ace719b96a9b", x"b4c12e265450aa49", x"99a227d45fa6d515", x"f695d4432ad80621");
            when 30870327 => data <= (x"800867eea819c5ad", x"e8010f1b360158ef", x"8f4874b21d46c2c5", x"d7a03f6f2bb03fd7", x"63f2c40339fcbc7c", x"61159280099c32fe", x"56a515e27e40074a", x"9e456f906e721f30");
            when 21875404 => data <= (x"36b8f3348987858b", x"037a47d2dbfa8f9c", x"7bb28cc46ce8e85c", x"bd910f6d66d0cb7a", x"1113e960223df166", x"717e9834df8e4cc9", x"4bd2be8d66320524", x"bf217739e5eaa5a9");
            when 5783221 => data <= (x"6714442d9ae8136b", x"282e884280c7219f", x"2a42a5fcfdf5c95c", x"5e3daa7d6ebed43d", x"c6b9677a5d3238cd", x"fbd15c4277dab812", x"3078a97d6725d1f8", x"1ca99dea7cbfab86");
            when 15029793 => data <= (x"a64d28c545d7f936", x"df8a696958d4f624", x"4e5d0569be7c5754", x"de4435bde16b3546", x"7c18c31e4c0c6dbc", x"b5dcc1a5a3276b48", x"6a1ffc1ab93fd247", x"98e5c3f4fdaf697e");
            when 27110767 => data <= (x"dd3cd252ff6ee36f", x"b3aa160a29719cf4", x"7ffbcb9d0bdee7f6", x"822746a9dc2be36e", x"dd92179c7eff4bbd", x"3441ef5e9336c5d1", x"8555cfda3d9b4520", x"8ae9b72b8a1d8cab");
            when 32460130 => data <= (x"31696648a33933de", x"990311ff71460c4b", x"6eb27182b19a9597", x"b7c15a38657d822c", x"a412a80c23f8c2e0", x"48e5f39d4ff85212", x"993ca654b79f4d3b", x"3d53b97baffbad79");
            when 33989135 => data <= (x"cd706a792c271988", x"d4d2a234ec6710d6", x"34075861366f705c", x"4857a6d0fc050e48", x"8a20b1045539b72e", x"690ab31a195c99d2", x"933c8b1b131d3a44", x"8efb50ec3b955c5c");
            when 27573985 => data <= (x"138b2f6c11d68dc5", x"e3a58750f60c7376", x"1b2afc229ad3337c", x"55bcee2c6c85d236", x"bff779d28aa58adc", x"2dd11e5926b7783b", x"38243fba5c92f119", x"a8aff790189f6ad7");
            when 20734789 => data <= (x"eb4ddaaf972ce9e3", x"804ccbc8119d4375", x"3734e84d51d384e9", x"7dba77cd8c93604a", x"86978c71739447ea", x"551d259edce764fa", x"05c01e60cfea9860", x"daa1b7270a769c46");
            when 30302775 => data <= (x"7885e221a60db6ef", x"2c78781a2c86e42b", x"2bc653fe6c139545", x"18e58c8dcc6544d0", x"f3553ff530bea974", x"e19603835255d8bf", x"fb19c459f93b2809", x"a448d791b25883fd");
            when 5047451 => data <= (x"1894a74188629786", x"9dfc90114b82dc8f", x"e6ec414612ac319a", x"e6aed9a062d2bedd", x"287120e330ff2780", x"716d4e1ea6e98a6a", x"67ebfdfff33da06f", x"03863d5e190144d3");
            when 9272949 => data <= (x"dc39b2ef7811d60f", x"0a6c250b916276c2", x"a8921c5f599b8c8d", x"6d655025cdb337c4", x"f201cdd0d96a2bed", x"255014ab76e968e8", x"c179a35d784fcc14", x"ce5ef901f177ec7f");
            when 3646244 => data <= (x"fd5c518bf07f649c", x"2d381bcb0d3f361e", x"3c52db043f87d3d2", x"495840898e16761c", x"991b09a92022aa42", x"0b40546c2fcda08d", x"40a07fb296a70c51", x"1c9ad4881e81f5ea");
            when 32984063 => data <= (x"c6282f78cdfe24f5", x"21397eb80f0e4189", x"78596c64c9beaaea", x"87e10d36b3f3ac69", x"b117be80ca26a3e0", x"caea89c26ac7e05b", x"34f12be41ef71394", x"1c4438c02e03c273");
            when 10499406 => data <= (x"6180326802ffa55c", x"a85880d2c9be1b20", x"8269b9d86e589459", x"9f735e343ea7b4f3", x"0ac7c13a319cf78a", x"a66e781f08662562", x"904e3614e4d81acf", x"6acd6d5fa5f6e137");
            when 33059976 => data <= (x"ac1e3a24c4b7373f", x"12c8c6d747ca8025", x"c362c799df83b404", x"7bcd05939f4fb186", x"54710cdda789fd91", x"4c5b6f875a048625", x"8b48982415f3709e", x"ff5965b94aafcbf7");
            when 20886463 => data <= (x"5fa1a84005fb882d", x"ecc8807820e93e04", x"5e58c920233d2f44", x"f8f1398a0c144273", x"c75a7bb1814fd215", x"9ef23230a552448f", x"8026036f5323fc8c", x"4d77f4bdbd6413ec");
            when 19088721 => data <= (x"e648c700f98b2039", x"d74b8ab63ccebe21", x"951de6f9bb077abe", x"fd8a56fc863b263a", x"fb9d894175f2e6e1", x"de9991cfd886b028", x"672813d8a182605f", x"4cfb1385f36d551c");
            when 23603795 => data <= (x"7b23723cda36fca4", x"2c9a6db3e1db6739", x"108268e9b5002bc0", x"0c35f5e0e272aa41", x"657c50da0eec7c0b", x"2b1576455d49a885", x"efc539ba5fa339d7", x"05467e4612377863");
            when 21452558 => data <= (x"6ecfec6b3136d98c", x"ad3bafa6865bdf9d", x"15371a1650fc8aab", x"16d6f27e332d268e", x"c66016c4b93fdc3a", x"aeec74e3ea71395e", x"9f8c9c2c68b99355", x"cdaacd4337a2b6cd");
            when 16889937 => data <= (x"8fa1c26eff022fdb", x"809b84a8cbc18163", x"05d50d37e371a2d7", x"daff982131bb4c72", x"a94a8126e38bc777", x"62632fe275697cef", x"ca0c2cc8aaae8905", x"3ad9d1aadf3314a7");
            when 16255045 => data <= (x"ae38cb2bbed76aee", x"80be961e98bb58a8", x"d7d2c6c19a5a84b2", x"3c8b2ab72ac5bd72", x"52c812b54493eee2", x"cb1d623264091ef8", x"3ed48ff967f61b6e", x"767bf5002f67b1f0");
            when 28763191 => data <= (x"d7f6335857ab008a", x"822ec2ea7c4eb381", x"398970daa120c0cb", x"83e71dfa8957c075", x"046964dde71ae29d", x"1d9d277c0f2fd8e0", x"f5356b53dacf7b4e", x"8e13fc57be87f1bb");
            when 5347204 => data <= (x"8745c0d17a22d741", x"478697a1db3adaad", x"d9d9b253ba0104f8", x"be994205213b3cfd", x"90f7daddafb143c2", x"880dc69634bf7d17", x"90e3c44eca6784ac", x"3206ef2fcdb864ed");
            when 5922431 => data <= (x"d5f1cbecf1ea3642", x"4a93d1a135aa0730", x"7b21cabe4e03ac9f", x"64e3e847588ed615", x"a34d692a2ce45670", x"cb53ef6d4e3bf121", x"8f8251736f14f1bb", x"2652f14f584c8fd9");
            when 13164287 => data <= (x"feae657c92e8b20d", x"5c458b1960031f37", x"f39905b53aea4446", x"c3db66dfbf9b6612", x"3dfab3c69564c152", x"3193e62f19d1f511", x"639badb4a669314b", x"ac2f17fd494c30b6");
            when 9295545 => data <= (x"8b354367e772cc59", x"56d95428b9294686", x"dbf861d5a2aca13b", x"c69cee4a6887e903", x"5f0e590f442185a4", x"f58b3a862a2259ae", x"26387cff6c39a40f", x"5b4db05cc7040d4e");
            when 543247 => data <= (x"a9cfe672d37c8d44", x"098a9dd2d4ff155a", x"e7609c1aa0b8368d", x"b7bd12193c4f2175", x"c43139ac7fe68358", x"c54327c62c15f2a9", x"1b08d7e2b1ec4bed", x"671be5b6c6a5389d");
            when 6606940 => data <= (x"91ad74a00925ad24", x"52e516c748e785ec", x"f797efb9203afd63", x"486cb521127e10e8", x"74f10e96cb96df43", x"a7118e80181f6b5c", x"584584aa1b8294e3", x"7fdae458d6a14f46");
            when 19348799 => data <= (x"e5ac6e76a427eac5", x"df3073ca452dabfc", x"4770d29d16ecfe60", x"d340cfdd6592b28a", x"a2360ea7c641d790", x"5622890ff23db0df", x"681671f1604bd900", x"a247890e229e7ae1");
            when 25098202 => data <= (x"55f1596c459121e7", x"6d07e176f47fc2d8", x"263d0da129d383ce", x"251e7ccd4a62e7ff", x"5b374817542bfc4f", x"fc5a418d5d5352d9", x"8f95cbd6502b888d", x"bf7c8b18c1760c65");
            when 5979247 => data <= (x"071d566184f04720", x"bd0ecde45e855995", x"870e6b26c5404753", x"087c362db827365a", x"37244786a17c56a3", x"5fcc079f2c24dd4c", x"dfd17464712ea81a", x"4cfef3bef79d5e9f");
            when 18678307 => data <= (x"5875f99f2e65a266", x"6aa8dce028552d3e", x"af385f6ea0870d70", x"c107f6c4900d8388", x"556f3ec22712220b", x"5a4b1dac1d8e0ac7", x"9ca709a5249f22ce", x"e0159593811f0783");
            when 7338335 => data <= (x"6be50fe423a73894", x"72837bc2e46386bf", x"fc5c53a42d1e0ed0", x"1ed0a99d8f220012", x"351bb8e446956eca", x"06b0cdd6011b3444", x"274977822d072d02", x"c099012c16f40761");
            when 2404810 => data <= (x"43e4db0bfc869b5c", x"0ad1692767521299", x"f7f23a3a2db440cf", x"ad282d6ce745bd16", x"ba49f4bcfd27a1b7", x"7811b1117de4aa58", x"1cb9d6e50dd44939", x"c86c69c2fd50e7a9");
            when 33739621 => data <= (x"ceb266475ca158b1", x"7cbebf835fa8d12d", x"bf84011a42485ba9", x"28ff0b630b5e80ef", x"e001e0d51b895167", x"0cc4dc6ff1e180c1", x"a50f2239ffda41fb", x"eb6a44ec58a43d1a");
            when 4199338 => data <= (x"8291ba13defb5700", x"9f024b0b99ae7568", x"2312d8b7b575563a", x"513d047df9828c96", x"64df26bd4f62f8ac", x"166fd1844f508b9f", x"811a2cce5e9d409f", x"148ff3fc9467786b");
            when 765239 => data <= (x"093bad40d178f934", x"54e75bda9214cd5b", x"2695a276d379ed01", x"05f22dc65b9428b2", x"0886afa4827761ef", x"39f213b438660000", x"b1a0b331cef4e606", x"ee8613206d1415a0");
            when 15452190 => data <= (x"7e4818d781b938b5", x"2051f97691e34206", x"1d1f8d5c9c4c3695", x"f02e505deb6a8c7d", x"233d73ab99e51c67", x"35116731beb2a18e", x"19bed0154b1aa345", x"aac9bacf07e7fb06");
            when 32651599 => data <= (x"1adb721edb77cb36", x"02d1d44cb993b79a", x"3dc3a42a6933340c", x"86e17a852c285035", x"07a2350da162739a", x"2cb5bc5a0dc7d8c6", x"a4c76eda6c19d819", x"cdc3fb293c63f5b4");
            when 23432710 => data <= (x"4dfe3e77bfb8e470", x"d3423a6c04a00e79", x"c722e596f01b5fd5", x"28acc9094873f7fb", x"15def368c1d724af", x"7c5a4c483b944896", x"16ab33c5f610a585", x"3b759a3c212a99b2");
            when 1012323 => data <= (x"6726de8bf445c33f", x"92df405755f0a47c", x"7bce3600b848be0c", x"153984590cffa9ef", x"0f5a916d7693c478", x"9e8981e0f9ceb200", x"7992e5c4895f8063", x"255f3d49d7fa7052");
            when 30441174 => data <= (x"152a43e690f1e1f4", x"388ffaf675d11874", x"f5cf83c83f15bd10", x"2cbcc6f0c07e673c", x"8209742550800f28", x"81a2b3477e2c9c9d", x"a8f37e12541290cf", x"808e78c6b53aff45");
            when 6581436 => data <= (x"bf407006b31543d3", x"39e1bec26e886aa0", x"de71257fb71fe498", x"a948fe75f47ea723", x"ce1995593a7d21a6", x"717dd98b24265f59", x"04831c87a374d8df", x"f2d57268bf387ea4");
            when 12557836 => data <= (x"78b3e10b86ae7085", x"4b2080e28987612e", x"7e533c8248eeb6e4", x"5233108110cb34e7", x"75f465f7caeda90f", x"5fbe911f290079e0", x"b5a32afd3e351569", x"569dfebf46042344");
            when 15580991 => data <= (x"65a2b3a5d6b8e977", x"4bc5d9cefcd14735", x"48691ab151e8ac7c", x"b136cd9de908b2e4", x"91d33b69176cbd06", x"bc8853a2787f56c1", x"9cbc9689aa1f1ff8", x"488c4c78d1bf6157");
            when 679244 => data <= (x"a8d8d8911faa1bdb", x"20f009a9e9fb509f", x"c77c15e4760ec89e", x"e61ca5213d4ef2fe", x"adcb5c666b6e8f2d", x"f944f018f0d9f8bb", x"b063963d0516a709", x"648b478ec23b121d");
            when 6240668 => data <= (x"fb6aa0916b978f83", x"f67b12c87cae1294", x"982a20d67ccde3b7", x"e9a5e21583596586", x"0e83465591199567", x"396a13d1467528b0", x"a22d8b03e78d8ae5", x"c35e0d7a3383b6ef");
            when 4626700 => data <= (x"3693e2729715440d", x"392ce3e358e9d814", x"7d8e1c130367f206", x"b9b1018bc1276b08", x"39b4fbd132e62fd5", x"64136818b2de9edf", x"824f06525ab1a1bd", x"8a842e418ca451db");
            when 26248657 => data <= (x"58a164b9b7e14b94", x"72aad6e4102507e8", x"44599f8bd70d9c27", x"758e020e4af31216", x"8cd7dd44979392ca", x"bf4e42d9c947116a", x"3d0f8026df503b9b", x"710479563b7e96f0");
            when 6083821 => data <= (x"74d0d2513b3ee499", x"45e3cc48b1c4acac", x"db0b5e576678118f", x"256d0d734e014b07", x"8a1aa1473ade559d", x"cb3f6552514f94f2", x"d7bdbada68bc46bf", x"0f6935a52287225a");
            when 31197142 => data <= (x"b0a4c5aa2cc931a8", x"c165bfec1af3bbe4", x"a55976ab0e759eda", x"191a681dba9ceb75", x"525014fdba6f6fcd", x"37bafe2e2363f89d", x"326145b35bfb2148", x"e488e76c0f4a022c");
            when 8617929 => data <= (x"d2adc570ae6aa1fa", x"109f3150f4ec05b7", x"9ff2e635981dd0ea", x"69eda549f3593856", x"bfba26d06b3bff81", x"a4767ab148d84196", x"99632f03d68309f6", x"bcfb648348344de3");
            when 18678321 => data <= (x"f38f6abbf794a38e", x"7c368feb99f50bec", x"47f7c307b0f0df2e", x"a8d3035ed5670bbc", x"93d695bb92042d0d", x"64c10831472475ca", x"27e0e5f83bd802ab", x"a95a4bd55cc2b19d");
            when 13881360 => data <= (x"e2bed22421ddd6ad", x"590a2987dc1c313e", x"8c2a75b5188567d3", x"97361fd62b256e88", x"9cc97d5eae3dc390", x"67643b876d81fcb0", x"e244aa91123cbc42", x"b927409594da5441");
            when 22504299 => data <= (x"b75b196acc59fb4b", x"e10c6dd4917df52b", x"b10e7f8657f7edb9", x"32aa805c26a4fe07", x"55e528f52ae0c2c9", x"75694b58d8456c9f", x"d514cdf866a6c204", x"cf135625c6898b23");
            when 4307680 => data <= (x"9d39d21a27012fca", x"79817ebb3deee7d4", x"d77e4af4cf332895", x"953ee7cb747e9dd0", x"5b5bd6efac12d5ae", x"9ac350db6506c5ba", x"b5b0997f9d60a541", x"9209f50a7c030d94");
            when 16010042 => data <= (x"d638c16370a59d00", x"c2061ae28180909a", x"b157d712f942f36b", x"4a441b5562b18ba0", x"503899e211f5b55a", x"a5576976ce71be5f", x"08708aa5cb7f75b0", x"19505ba2221c23fe");
            when 3180353 => data <= (x"f93a6bdeb46de69f", x"295c605980101f64", x"ab23b86f6d8a0943", x"b9f6885823486a6b", x"3fe67cd6fc212c37", x"342da5d43733e3db", x"135ab6b7020c0f87", x"81ac94239e5af92c");
            when 10109779 => data <= (x"eded51cfbbfa66e1", x"90852b20fcb277c2", x"40d56ff4f6c1b964", x"2449549bbce096c9", x"4ce794ab6e10a948", x"177662add78b67ab", x"5560958c7fd5c2bb", x"f9da4987b9a4049a");
            when 19354483 => data <= (x"ccad6f215a1e4ef4", x"034a9b0df16648af", x"49de96d54ccce9de", x"9360f0fb123a4600", x"f8b59fc7622c56a4", x"5bbe5a2d360a9636", x"510f3e6cf9964ce5", x"eef5070a4fcabd6e");
            when 13102218 => data <= (x"f5893ad5a79bf114", x"301dcc804cfd1061", x"8edda5ebf17dc131", x"b1742814758558ae", x"7c0d41322b7d2557", x"3478ccb5d81a1dba", x"351f219d1fa99b9a", x"e0aa194e68867b18");
            when 9468230 => data <= (x"2d17fa3058a48aa1", x"89b816aeb246267e", x"f660b9c22b4eaf32", x"9054c37c37d3d57c", x"d55be506602464c9", x"308454b7f4a92966", x"0565888005b0b4af", x"407ffbfbdabbd119");
            when 15358020 => data <= (x"79422ef15c7ff886", x"6ff236c822d25f32", x"608022ac4be9076c", x"efa937837d4d05f3", x"8add4ae74ba83911", x"5bb0c47503f20122", x"a18bc536c4612932", x"9d8f7e49e7f45461");
            when 9610847 => data <= (x"8c8784e850801a0e", x"11116e872959b78f", x"fb3de28d501f0159", x"dbe07bbf4fd6952b", x"cb0bcb6c89dbd978", x"9c1652b3057620f6", x"d31c5df8d1a3e46d", x"afdea690b7803d1e");
            when 29960349 => data <= (x"3f2cd7ee8738a040", x"bab952b7735f6260", x"cbeee6bc1434d4da", x"944dc4ee1d1eb238", x"28bac4cb497e4de1", x"15516d6d5b52a420", x"372eddbe4e668569", x"e2ffdc548246ba7b");
            when 19703837 => data <= (x"ba6632190f89a647", x"bf54780900ebeb28", x"e5e41da7c3ea9fff", x"655e78b8f55d806f", x"8051ab4a9bc429c1", x"67dbeebd1d63e7c3", x"d521455f446614fc", x"d4549d26b9c2f9ea");
            when 24283236 => data <= (x"5277dec96538219f", x"b750023b998fe247", x"4cacd482a82c3a90", x"ba63cde9e91ab24b", x"6a54db5d86b764f4", x"619934f3a3aa4380", x"2a08341d067dfc9a", x"84e9630df7b77ed6");
            when 27680284 => data <= (x"bb6c1a7f78e91a75", x"c8a85c7f7d951a38", x"df841b5dfaef3bd6", x"0020a7760dc69474", x"2d3e19aa58b71ff3", x"848530aa3ab1d7dc", x"98a4082292b5cada", x"8d9fccc85ee9b04d");
            when 16460005 => data <= (x"72528362cd513670", x"273ca44cf4001bc9", x"1373d6dbe6147039", x"4e9dfa4302610131", x"9005c6ed53bc0223", x"5e3ffdb99e130d7f", x"b38ed0fca171f9e0", x"16e8cc929ac3b94b");
            when 32777317 => data <= (x"6d0dbe5617feb085", x"bb0815dffa77dea9", x"5a796ad058f024f2", x"5520e01b27cbaa85", x"edc05dfd4a094593", x"05ad97ba14f3a098", x"e225a998c4c6ef3d", x"76b64b5cf7ec6195");
            when 25436432 => data <= (x"1aa56df33a5454b3", x"4b6b9852b5dec1ae", x"c5426d0afe5304a0", x"e8c357aaead6b5b4", x"1259e6fe8d4fa7e0", x"0ed1e1850748ce92", x"5fafdf4298cf0960", x"b6099d9ec2bdcde3");
            when 31821693 => data <= (x"9b2acb32cdf2fa24", x"cae43f3e34956f1a", x"670ebd9f85ad8129", x"6e54de9a1b294de7", x"c339816bb0733c5c", x"c22d46056442cf79", x"937b401ed29362a0", x"b29289dbcad92a3d");
            when 33764629 => data <= (x"bb0472cf898675d4", x"8e8b72d43c0ae42a", x"27f4f2a2e4db4304", x"0c7fa2136b3289d0", x"e5a885513570382b", x"123e570399fc341e", x"81bb8d40e84e1412", x"5e293932ae1b7e05");
            when 2442634 => data <= (x"0d956b34b2b3b621", x"d38069adce4737d7", x"15d968f27ed0410e", x"ba47694e1f93af24", x"2b8981cbd436e402", x"7a11ad28819e8fc7", x"929e957a30561a8f", x"1793fb45cc8bdbc1");
            when 4650468 => data <= (x"0ac49b25b39b30dd", x"c76c9b8cb4487bb3", x"96491e4ce2d29b6f", x"803cacd78cba1ccd", x"03e7078408c8e3e2", x"11789c911c2a59b0", x"aa823b880d3d5d4f", x"bb9c32e0c969fb25");
            when 17397371 => data <= (x"5894af80f8ff9acb", x"6e3ad73d10534079", x"1999608e2b33d47c", x"f5db2b21092a1cae", x"319f9b26821f360c", x"9a116818f8b68c42", x"b2ecf165bdbd1d96", x"948a547c332ec89d");
            when 23449231 => data <= (x"58d9876f973d365c", x"9a084a484d43ee3d", x"8f55a98b4f7813b7", x"9adfb9bf4548de4e", x"92438dff83e04c6d", x"7b4da042d158183d", x"47dae789cf95a35b", x"b4955a56fd5eca37");
            when 32405020 => data <= (x"6f57aeea1eb08eae", x"d8e914c54ecf8825", x"944b5d974354363b", x"520f6086daa591e8", x"6ff9da0bea0e0c1b", x"9c31ba752cbdaa5d", x"66c4cda166857826", x"7d109ab2fe62bca4");
            when 33263988 => data <= (x"31d17ef1c3dc8173", x"84b700549f775b25", x"a0bf3838afb3b5a6", x"68560b9ff43d239d", x"4f2db0a8bcde0d4d", x"dc7c945783cfc48f", x"0adc10e59a291b5a", x"19afa2f9ba8f3a4a");
            when 23774893 => data <= (x"c37ff0a4ac82658f", x"c012cea12921aae7", x"5430b6e48c51cfe5", x"e21e8d3a915765dc", x"d85a26cc944b865f", x"6af34d2cc5a13a2d", x"8176289657696903", x"b38e25c030489915");
            when 6700671 => data <= (x"b461ef8dfbbd8e08", x"c4f29f7a9bc63770", x"28f91a8ff73e1da0", x"0361272f1a9ee0f4", x"0a5111979f5633c3", x"740fa41675367361", x"cc21a9e859604777", x"1d6e3ef12b4b380f");
            when 16210389 => data <= (x"901f1d995939076a", x"f238752d0a92425d", x"2730e894dd4e8247", x"0dbe346481952ab2", x"3c0ace6427f7d5bb", x"faca22ad584fd55d", x"ffac9cb57db9cd83", x"1bf93146874c637d");
            when 10885161 => data <= (x"d9b46b7fc76167ec", x"869e0d7e7f12c60a", x"0a771fd1521d3ac0", x"ad1c03fd6f742eba", x"9720ba60c9b7171e", x"00a96f8ff776f42a", x"13fe6dc0f5b4ca54", x"e5005a19e764b6ff");
            when 16754922 => data <= (x"d51c3df5a439e42f", x"fcbda1522301b4d8", x"ac166740106181c9", x"3778f06e42e227b1", x"e261bc44aa643d5b", x"b41b472a7b8fa5cc", x"e607f457a0d4f7ed", x"10f33a18e9e603cc");
            when 10821038 => data <= (x"fcc83febb5ac9831", x"c7fc1df1d577f05b", x"4e0ceb4dbd40fd5b", x"949470f061f1665d", x"53016c3772634ddb", x"8542ae5e4cbe47be", x"c8d529fc4e7de181", x"e42f28a175e7daad");
            when 19474925 => data <= (x"294d35f807b4b8f6", x"39300ea7bb165cd5", x"12d20da38fbbcef7", x"39b4f37310b5fab7", x"3e73d65dfb691629", x"1b5241724709b9eb", x"4738e2b1eb454502", x"5736d2961c600b17");
            when 18307073 => data <= (x"fbbead6122f574bf", x"3fc24294a502557b", x"5a78598cd4d588a7", x"61de23d9c6febdfb", x"eebab4d410b40412", x"405cacfd5a00441d", x"e7609e887a27e6e4", x"0da30c1b028f1003");
            when 5762716 => data <= (x"2aacd486c61f0aa2", x"39d51e55d8485ce9", x"1189118d96605def", x"08088b000db63f66", x"027d9c1038811381", x"b4d8d32ae51fbbae", x"e9291f5c0443c539", x"25fee741603b8015");
            when 13181321 => data <= (x"0190a864f46c6b2f", x"c5c9f5e7464f78a5", x"b153297a80190364", x"5d0122d8ac39b758", x"2b37654cd8d1ab6b", x"3fbc9c9316f3017e", x"22bcbe2104c6e7a9", x"b685e2d022a7e123");
            when 11740609 => data <= (x"392ccc8cad2e0bdf", x"a426bf9b7d72159a", x"5920433887a68293", x"549f9e8f1d390f3d", x"4ad439c920c0664f", x"7b0e4e3c0acaa238", x"482e06d7280dd35e", x"423e1b1bf80ea040");
            when 15047731 => data <= (x"7c404a3a80c91d8d", x"6a2693e0aef93339", x"1a376f0d7cd6b7cb", x"3342cfea4ac666df", x"11c03a9568159a67", x"ab84e5bf8a0afd36", x"2d9f0f0987dd4205", x"000489b17c1fded2");
            when 17916156 => data <= (x"003b473e00bf41ac", x"e720049fa74e343c", x"6ccd3cdfe06bd364", x"71e2e1b2169b486d", x"e938b64441d51f11", x"d5b2ab4a2c306ec8", x"c732b0d01841bdb9", x"04d7297bb45b536b");
            when 33809147 => data <= (x"2287a50daa44aeb9", x"ee33bd53f0fa76cc", x"ddb443f096231f9b", x"d73e0f1d64874946", x"50eb4470391cb09b", x"e786e63a98290d91", x"ad461827575692e2", x"b2d6b240553d2e9b");
            when 29496695 => data <= (x"68c9c0bcd543ee21", x"47c3e9c365f9af24", x"800ed6cbe29dabdb", x"3b53c0a4f0542fcb", x"3a582a8c16261706", x"efa9c523fbd113d7", x"84bd1ab177a74064", x"e4c0802858ed1989");
            when 10825167 => data <= (x"0a20afb9462080db", x"4310efb49940757a", x"b471acd9dc8b9ceb", x"01329aae6c1a9a72", x"a11fa191256b9651", x"5ec042b1ea80f0d6", x"b2003b097a0ddc89", x"0dbfe219097608ac");
            when 27913982 => data <= (x"1a6f0edaf9f1105f", x"9252ea75c6ee4b51", x"bb3f5d829e5bbeb3", x"d0710b2987e895c6", x"a6eea4de954ea887", x"0fbcacacff3fe024", x"326ac3e2c3e69895", x"87938706c9d4d831");
            when 3191943 => data <= (x"74be396f43ab70f5", x"1691e3dd727533f0", x"65697264af904c10", x"c6c47a86e4287c2e", x"effec41ec3f3ecfe", x"b9191de61858d4ab", x"cfb014d38c51898e", x"ed172381c2ce24db");
            when 29107630 => data <= (x"8fe886ec83e4bf6b", x"9d4b624edc67af2a", x"8686950cf16411e0", x"47b814971336bfe9", x"a991d5ad59a6b634", x"26d081a5ce6c2b43", x"41bb8ff7de0face9", x"36b6b4f669aa91e5");
            when 13844024 => data <= (x"8a8b6caa5990f38b", x"53531eecaa4f37c9", x"9cc3ea844cebebc3", x"1654de69d0533fd9", x"833791ae91d77286", x"c4f0d043810d7b9b", x"8c839678939d63a2", x"fb5f61f873e1932f");
            when 2645057 => data <= (x"8da0ac8c519fc225", x"8f1dcfd3a9e99462", x"5a30ac07596ca41c", x"1bafe258a45be430", x"496da09c2916dae5", x"2680d406450941ac", x"3b14857048834667", x"b3acda22952871b2");
            when 18861445 => data <= (x"5c46e44042a180af", x"cba182d1746326fb", x"4cfd332afeb53402", x"e045b10ba7e4cf75", x"3fdd27a625241860", x"295279604cecdf4b", x"1ede4bfe17fa3c8d", x"93be9db720697dce");
            when 15081030 => data <= (x"81dd8f5297e193bb", x"249065b2bfc2bc7e", x"f2695c7b6e0af036", x"396ed577663c6ad5", x"94409bae1e84079b", x"d726d47323535864", x"16eb3fd5bc6d4cee", x"11c9e970b5270d7e");
            when 11213990 => data <= (x"b8cbb46370319287", x"d80b4cbbd9d72142", x"2d6dcacfba0f46ee", x"c08118b6f80c77e3", x"f84496f0ed180fdf", x"3a7b4843229336c7", x"93ac1bbba8689062", x"25fa8bc421fd9864");
            when 15838912 => data <= (x"19f541aaba86ba78", x"9f283bfb8fb163a0", x"2a42da262a9ab7b8", x"b0861aafa8dd63b4", x"2c12c584748c25d1", x"e82d84e5fb26595f", x"a1eb1011d65f5088", x"03d00973e0a47499");
            when 15367977 => data <= (x"988701d725cfbd3c", x"98c66a0d65d932a0", x"7fa5683813c32ae1", x"bbf53d1251f03105", x"ade2b36fb14462e1", x"0ce3a6855a45dd8f", x"63d9fd7f4c96ff0d", x"21d1705e0a2d403e");
            when 14904490 => data <= (x"b84be2fab1c1e39d", x"af5b1f01d65fb16d", x"148f9304f9061835", x"748ccb4d4d56a848", x"8575fbaef2baaebd", x"9b1827edb7f64f29", x"07141ac8c227c0c1", x"34e4b7fb448f8c73");
            when 8007926 => data <= (x"00fc1bd5b8bc994b", x"fd96ce9aa3529954", x"fee576a817682f00", x"ec0e497711a9e4f2", x"fc36e4230caf2a58", x"0d59ba7973b5f4eb", x"fb3287976abc5274", x"1fdd65fcc4e39681");
            when 9407439 => data <= (x"42d54d1457cf0d91", x"92e6854be669355e", x"6a6d50fcc06bc53f", x"a292c3337412ad0c", x"b8982fa2a0e207e3", x"805f9dfd37ff4ce1", x"6bc8d44b33617427", x"8c99cff50b00fa33");
            when 18180418 => data <= (x"500c15aa0dfe7db8", x"76feef02efb2ecca", x"fefe82e518122647", x"218df7e3e4e06d37", x"7a033be679458c51", x"81d1d59251a42ff2", x"c91a32da2507efd6", x"55cb810f5b5fce75");
            when 28376232 => data <= (x"ed51fd8db462ed13", x"90ce9cf760070b83", x"cbca38a4ef005e0b", x"dfe6147cff0dea12", x"14726a5b8c88cd1a", x"5acd44b1baea745c", x"20d147b89b5d3dd7", x"2cbef4de516b0557");
            when 7789908 => data <= (x"086abc03d87c0981", x"2100be9af239af73", x"99415389447d31a7", x"4d05e36bbc0e03ed", x"a29b0909008b5e3d", x"84c7c60e847c3170", x"66895cf50b5f897f", x"4eda52cb9a32ebf8");
            when 28972808 => data <= (x"94bfc06ce39a81cc", x"5a004184053efca7", x"02b0c178de11f009", x"b064924f677db1fb", x"e7ee4fdc3492fd72", x"1d56c2c81ae82a8c", x"cdb6461f4ad58b40", x"e6dc51a65d1c8015");
            when 22632814 => data <= (x"18e133596a828edc", x"0d5402c7a5511390", x"fb0bd96342b14466", x"d92813332247c99f", x"08e0138c8930424a", x"f069eb348a12f1c1", x"015c99d9b96c96e3", x"4134cccaabf26aea");
            when 17160394 => data <= (x"bb10ae5624f74552", x"9629436c5825c314", x"cd8834f7391595c7", x"fe991ac5dce8a4ab", x"71e26499abff8ae9", x"6cf997362e372fea", x"3a5f505a3dc148ca", x"aeeb89bb4e4329c5");
            when 9162461 => data <= (x"f85a15ac757e4dce", x"d3958a949fd17449", x"46d659660ed235e3", x"954e8b7cf80f564f", x"62490b1b12b12815", x"76ea618b0de1495e", x"655f98013d87036f", x"28a84ddebba25fbb");
            when 18637262 => data <= (x"b0f006bb40a78aa1", x"8db44797c4f38ffd", x"65377414687810e3", x"8560b4387000dfde", x"df22a6e2b3c01b23", x"657fcd47a9f88656", x"a3a6adb5dc0f7a52", x"ec6a66d7ecaf451f");
            when 16359356 => data <= (x"811e4d96f3b3bad1", x"045287253eab5ece", x"4993d5264a840e70", x"0b19feb6ec9d7d0d", x"e01dadd50992428b", x"c6c2a4d174960a1a", x"56062f1174db3a61", x"483e938a8ec15064");
            when 7575595 => data <= (x"b9f50193a9f02ec7", x"f4177b3dd0430395", x"2c6c50d1e47da22b", x"c47bbdc663c081bc", x"4b075ba937fb1019", x"c5ae0c3f910122a4", x"5bad2cfcfb2da260", x"f82953aa73ee7a24");
            when 1430074 => data <= (x"a661e9910bc27ff8", x"3136878449cac9ac", x"197b0f7b0564a963", x"5a27b33fdea40022", x"b250fe417e053d1c", x"ecf185d853adb340", x"b85fd280368ab619", x"1022bac58a53ea0f");
            when 9366695 => data <= (x"dca989cf04405cd7", x"0420bd2017ddb782", x"9473a2f34bc7f78e", x"6ea70119c70f15c0", x"3ada210e4aaec3e5", x"1ae6ca3261f3f9af", x"e424f51562bbf404", x"7c572298db0c27a9");
            when 15501211 => data <= (x"fbe6099a2c9ec7ca", x"c1d782f095a3b3ae", x"ed78a48109b9040e", x"26ad4f58ab4b1243", x"2aeb69a1d8b9865b", x"635a4bb4051b9f76", x"7c7de27ac43622eb", x"31b6a638a9be24d2");
            when 2694534 => data <= (x"49238703b949672d", x"264aec6720a688f8", x"a5224147594e0f93", x"2cc6f2106bac9b78", x"43820065deb38996", x"6bad19012e27f648", x"86e6301c29e2162e", x"639e83d50f46f6a3");
            when 32400022 => data <= (x"68abf8131c654b45", x"b86d1ea44c6c4a1c", x"99540a1260d8f980", x"0beb00e0c321ab62", x"d51105c597c16ad7", x"fbd995e3dc4056de", x"ce8a93e4d3a3c1a1", x"82e64f7f8f0a30e6");
            when 17175473 => data <= (x"f557c8907f782191", x"ce9ab4d1a08d1b8f", x"93fe50fd2ee990f3", x"26f3d9126938ffaf", x"3ba679933d4f133c", x"b00d361aee1fb54d", x"c5512ea0ea78240e", x"ce7eea108aa2f715");
            when 32157558 => data <= (x"a49ec055d0505070", x"8bc405f1416e8f0b", x"4f018166247bb66f", x"c60ad130d68a415a", x"3e58777099bea2fe", x"7d26ede612c58470", x"06089adeb6e424d1", x"7cbe4915efaec237");
            when 26634022 => data <= (x"391eb19682e16c9f", x"c0529eecf6da0f19", x"8a2f449fe95e90a6", x"aecb53dd0fc61141", x"b1954af5c6f35834", x"8255142836622bc8", x"773b6c0f4c0a313f", x"ac4ff0843dcce63f");
            when 6818668 => data <= (x"e33cf0abd6ba5108", x"6c5c3ea448d0c0fc", x"efde96581e625da6", x"e420a019ccf8dbcc", x"b8de2a9e6af7c406", x"4e688b8d259f9f03", x"44697e1350c926d8", x"e9a0c8241e9abd2b");
            when 21966036 => data <= (x"c22c31d7c3c06e6b", x"c1ef17b38ff81429", x"3816cd3cd903335b", x"a09bf493b4abe9c0", x"6a20792204a95155", x"b0c705d5b8ad4208", x"e0c8efd622db2261", x"a308df8d47399ff9");
            when 2377318 => data <= (x"f61009cd1b7dc138", x"df2d52126c6b1c46", x"99e74886636d8b29", x"35379b775a82a6b8", x"69967b7f96c24aef", x"d126dba011aa4181", x"79aa8b0b5fc7069a", x"65a5493e208f92fb");
            when 27171804 => data <= (x"a05f91ed9a8318f0", x"f32d6dd78cf939b9", x"2f621248e98d3cec", x"bece11ff217b976a", x"64be39dfc745410c", x"ec147e6d4f538827", x"bd584c4f8be06348", x"98bd3d2a5c48849d");
            when 28656803 => data <= (x"1aee35858cdc2322", x"e4cd0b388e0fcef6", x"9407264a52ee25bb", x"d5f0f5bb64ddf038", x"86ff0539d7d7dcc1", x"71c253ffb5ccb69b", x"00fa1510ca625af7", x"f0616c660e516643");
            when 28423071 => data <= (x"bbda09fb5f498e28", x"d17eabb67ffbd7fd", x"c546e0c99ab9885e", x"98a11fde52c4d4e3", x"cd65791a3fcf61de", x"4a24ac4c13a021c1", x"9104b6cd36464615", x"651da54d9358f171");
            when 21695436 => data <= (x"2aab7b99f09e17e6", x"ced7f0cd154ba42e", x"c1c36835904bab3a", x"3f9b5786c50d58b9", x"1fcd43457b053f4b", x"5746b220fc1c1661", x"d9284ffe7be8801d", x"daaaa218792f4467");
            when 30502925 => data <= (x"f75d565b21cd33eb", x"d92b7e2bb40de87e", x"b271e1e1e652a585", x"defd3f3e1e11d2fc", x"2ac998665eabf2b1", x"1db84231b10e9ad6", x"b0a6499957c162b4", x"11f686d0d1b9faf1");
            when 33364760 => data <= (x"87735334117ad8fb", x"0116961ff325fa77", x"7d51db4b3219423a", x"593129deea1998aa", x"e521d72cb01d3a49", x"afb6d902dff4fa6b", x"2852db9b318024b9", x"8e2b7cdecfe43027");
            when 11533355 => data <= (x"73977073681ba8ff", x"29deac23f2632a41", x"3692258faaf5e952", x"62eb3328a1fb2603", x"7e010d8bbaf13ff2", x"35c148b3a5548187", x"86f83c69074d80ce", x"a1f5216de3264cba");
            when 18852106 => data <= (x"09d7e97cf8051c96", x"151bb1f04bec4f6f", x"443322667019708c", x"ef5e1d64c92f9df6", x"631538821ba511a7", x"4b00010c5925bdd8", x"c6374ab03dd61631", x"5fcf084041ccc941");
            when 30253065 => data <= (x"f2da18653ebde54b", x"d7b2a76dbf8b5606", x"d8e141d4f0d044f5", x"b78a33f07d89789e", x"a471a477e45c51e1", x"04e95da5e10c3ac7", x"54efde9ff6b647f6", x"379edf7c91101a81");
            when 5807298 => data <= (x"b933107a6c8f7849", x"8bcb2bc1a0b0cfe2", x"ef3619f080bf0256", x"16a93a753be6e8a8", x"ee5b219559aec79a", x"1fd733f99e2c487e", x"97da8514f9171098", x"4e2b393a7a664c5e");
            when 4169798 => data <= (x"c295631453e43004", x"256e0526d8ca0421", x"4747965540ab27ad", x"9d96c42dd90e15ba", x"d63132978a5b1b05", x"cb8450d23f567da1", x"43aae4480038cec3", x"14f7af8242d685ca");
            when 11024805 => data <= (x"a43b9fda6262ba54", x"255319d8aa4cce97", x"50e87fd7d0047fc0", x"d27e536b6e78b8c2", x"9ab300c0f8c6063c", x"e7b552f274a07d5a", x"1c3336b2713e4717", x"871b4a7e419022c4");
            when 5132370 => data <= (x"a72cbb01e849f548", x"b357ec2504cc6fbf", x"e8d90d3db2bcb443", x"6d24ec8ca57b8bc3", x"7329cf0da0ea669e", x"a9be1c45dfa4bef5", x"77c86646246fea56", x"c539e781126c0945");
            when 10461288 => data <= (x"ffe9a79732c0011c", x"34708f5d279a30e7", x"f190433de435cbe1", x"e9b58dfc67d06dcc", x"0f6fa310279198aa", x"f0bcb29d0ecdfe28", x"8e792b50ad76c1bd", x"306871a6513c5a45");
            when 12018612 => data <= (x"75ffa05c6af5dc1b", x"7e3ea195c0d8851a", x"540a009341fab0f6", x"7a2e982ca53ad3ca", x"dc4e91c1d8b0ae2f", x"d1e9ba2527c37249", x"00edfe2be03a7ab7", x"f272f547f68979f5");
            when 30792832 => data <= (x"45b167089fc58a65", x"e7d4744662356dbd", x"78ed481505b9b665", x"51c7ec7efc63d195", x"d27e7479e9de4bce", x"b478571123afbc7f", x"2389edd1463dcbda", x"248480982b33e3ac");
            when 3710806 => data <= (x"dc8a92d7a66c32af", x"19c31d0e0730423a", x"f6f7af7bec585006", x"9eb0f84f285e67f7", x"311ec71de9b3fac7", x"41c5808887cb4ff0", x"741ca52c0608f38f", x"37e9165499930057");
            when 26220330 => data <= (x"741846c50d2d7321", x"eba3cb8abdb6445a", x"2bed2dc571d81bfa", x"3d69d88deb1ebf67", x"bd3c556d9d6323bf", x"44cba9fcce9dbc4c", x"c10aa2ac3196814d", x"756f3633734672c8");
            when 26942966 => data <= (x"259779f1d983e1ca", x"937296aa002910fe", x"e3fe1d1638d95396", x"4003fdcbb9a7596b", x"3d537424893703e5", x"494aff10b5f3c74b", x"9eb3925b1d09aed3", x"66b3048304cd6c5c");
            when 22618841 => data <= (x"80a4c807f0c1575e", x"42823816a5ab0829", x"ca65f2438d50598d", x"6644e5e76684fbba", x"08a46918c3844161", x"34cc0629aad93f34", x"40458c7af4f55f06", x"f358372162886e7d");
            when 17700634 => data <= (x"f79e9a047bf6ab47", x"d59339266b89e99e", x"e61f5c6fdbaba1b3", x"6d068d06c37d7c38", x"5ca8160418bac80a", x"814a36f3efd51b5e", x"5cff1a0eb8321fae", x"4592d6e0851a03ff");
            when 3970790 => data <= (x"240aa8716e06999e", x"2f9acb76282c8d57", x"3f2fdc628222f057", x"27609d120bcdb855", x"4acc12c2b0311440", x"4bfd730417d32455", x"3a9cf942916c711f", x"5eb234282dc64b7e");
            when 3718507 => data <= (x"44791bd7f2d054a7", x"a528f36a9a71f19e", x"18bb8f180eaafde6", x"da3949c39c6611bd", x"9f90594ac17ebc62", x"8b277a025e5123ac", x"009f11989b7033b1", x"43cb559aa58449da");
            when 17168069 => data <= (x"494993758be2b271", x"738730fa764e2d90", x"392496a926a18b83", x"f9d437d415d6fb1f", x"4295b9d8989e0b50", x"d32a5e67f35e4f90", x"065c70683ea79c09", x"e4490e2d1ccc0bc9");
            when 13155571 => data <= (x"4b94c7b645fdeeef", x"505e0b94bd036c37", x"2043238abb77edf3", x"4808b398594a6e39", x"4f721c28cd5ea033", x"1ff61a81ed78d7be", x"68fe6a4a2c4e3b0e", x"67b39cc43c452bdc");
            when 8432775 => data <= (x"ce8ed4632a53ff6a", x"996e1d4cd1b05ea6", x"b483d782b308207a", x"bff19fa665dceed6", x"f7f50007b72eb48e", x"3c8ec21a310be818", x"bb236aeebfc11b7b", x"b24541d2662441c3");
            when 18913640 => data <= (x"280280b0dfff679a", x"925bf8f72ccbd838", x"27a4a256a5e8a825", x"0ebd9808ae491583", x"edc6a7129f79fafd", x"89a2d6f1806b0a92", x"c7bcc2261a3fca41", x"a1b17de3eec590b4");
            when 12743252 => data <= (x"cec77d83661c0d0d", x"c318582080674e36", x"9a12f6066aa2226a", x"cf99044c3397cf63", x"aff892e70836b638", x"eb5c6acbca7cd0c0", x"bf967e39f14ca0fd", x"ad2ab62c8642b9ac");
            when 26002121 => data <= (x"80194750db795c65", x"0af0f2b128134610", x"8d088af3b1ea8f14", x"73ed106d8d223b0d", x"000a5eda2cead80b", x"ebf0c128d2b31831", x"12907be2844f3216", x"842f3ea0c580b874");
            when 31927211 => data <= (x"f6d0efd3a60d2d8c", x"87294cf2bcd1c0f8", x"9e2b16a91e68be49", x"51d2b2fb75ed2dde", x"2bc0519fa16fe705", x"0cbcab0440843c51", x"9a9d0c459e1f2854", x"e0f6d3f643cb7e2a");
            when 26472753 => data <= (x"8eb2511fda17b1f9", x"153f15473761f692", x"3c5d6911137db966", x"e0918e9ae6dcbdda", x"16af4dafea107618", x"15bc3dd592c5399c", x"ae0c4dd3b34e1df5", x"876725b80f564025");
            when 922122 => data <= (x"263f14d984ead2d4", x"caf71a495947783b", x"c12662d18efc4977", x"a19fb900cf7d4d44", x"819a30bd98d85db9", x"14436c169c1dfecd", x"c0fbd75fe912678f", x"44629458b9a2842a");
            when 18608754 => data <= (x"791a7ee39f2890b6", x"409c25afb0132374", x"70363b890a92b8cd", x"8983062ae02bd92d", x"3d7c1ec302ff8192", x"3cb3ae8f757d8f10", x"9028fac09930f9c0", x"40d7b4361ba2cb0c");
            when 20748160 => data <= (x"5dcbeae529098423", x"3129c6fa10e7589e", x"050f6a054c72394d", x"b382f4d9b616038f", x"f56497e0c198bce7", x"5215bfa50e66d139", x"8bd23f8838864cbc", x"bbd749f2730f54c6");
            when 4615235 => data <= (x"dac280d2665da103", x"97b6637e63d9afae", x"e70825a8906fa9cf", x"bbbdacee85cb7b3c", x"2d71b9393204adb8", x"6f2942d4c89a22dc", x"4f656d8a4a947291", x"b79f2ab004b58992");
            when 30717364 => data <= (x"1e98c04a239a5315", x"be72a142f2e22ff1", x"aeb17c26d1215ac0", x"af5c0ee85654f2c6", x"563cbbec1f776a83", x"c8a14e30d78142f9", x"6a80a7d8408857b8", x"b16983c3c97a73b5");
            when 29628526 => data <= (x"e0867c0890f2ecfd", x"42a0c35229128459", x"ee69f2ea6798353c", x"16671ba309b871c7", x"4ba069dbc9649dc9", x"dd4302a3868d4f11", x"79d4c60cb10bf881", x"6ef118880c5cdec8");
            when 28578268 => data <= (x"5c07fbb689e7c472", x"14f797aff01a7aa6", x"74fdb43666e7bfc9", x"608fe906c122f25d", x"b919b1801908ab7d", x"60045861406c29fe", x"88f7254a3b449f87", x"9abd3ef64eb88bf9");
            when 14823988 => data <= (x"7fcfc8705621010f", x"9dc3bb3cbe97ef16", x"e417d9ad2f673b87", x"600afcdd129d2148", x"249ba18e4414a952", x"07eb1b2b151bb3e3", x"5d3f5a0041fe8620", x"7b773f7a318a1c0d");
            when 17747190 => data <= (x"bf3d5b7156e63d30", x"9a9ab9b24e050674", x"91e108ba3816ccc6", x"011d0be6f4340d7c", x"422b139805e04881", x"c20900a15d4056ee", x"4462fa23601416a1", x"676bd0caf49e95a7");
            when 14663149 => data <= (x"48610263ba393741", x"a1e4806b43b747c6", x"1cf81094fdfa347e", x"a3f0f29c254dad1b", x"c0f6fa0710f9b8a0", x"0aa16b2e5df5c1f7", x"b39e85ab687fee9e", x"d8d1b0e85207e72e");
            when 23457177 => data <= (x"5ed0ecfdb91ed50a", x"76c183f550cbbb7f", x"1e2aeebebc4e5c13", x"f29281fedda9f9ba", x"bd35cf54d7d01cc2", x"6af2a1b4a2cdb7d6", x"e3cda937ccd84dc8", x"51c292ea8ef0fbeb");
            when 28413938 => data <= (x"18d68e2081116284", x"750a471f6ddf561d", x"2ff09f6dcbbb0c09", x"c0bc1a8875cd993c", x"ef69db8d8d3ba1f2", x"09c07f9d19dfcbbf", x"4f2e42dcfd3bb2de", x"9f2ec328b68f9fd1");
            when 25333889 => data <= (x"0011e3f13e0833db", x"21d8b28bf2de1f35", x"1a0b12bb96f291d8", x"5400e30cb7b14bee", x"eb4c037442e5d6cc", x"e5426e77cd1d8bcd", x"6627dc9476ba8dc6", x"648d88a16fb16837");
            when 29927220 => data <= (x"3fd0e4fc29fb8047", x"aa985d196f968eb6", x"ac5f48a81931268e", x"c9f05991fe816d5a", x"3bd11cae596641ba", x"1b88a2b767a2bb80", x"7d90640892689773", x"23890e704ce77c41");
            when 28112745 => data <= (x"e9ecbb312a9b850a", x"c34037ff3d644351", x"a3633372c927c317", x"5ae00f08cddaa97c", x"4fb5418b64c79a69", x"991ea92d8370ee7b", x"041501dce2d05a8a", x"48b03dffbeda9a4c");
            when 14587321 => data <= (x"590779adbbac2eb2", x"5eb3f809ff19ff8d", x"20cbb5b4487e6f9a", x"e37113ce980f445c", x"53fde6bfeafc0910", x"df2fd46bfb97abaf", x"f11fc47194b0192d", x"63e5bc9fefdeec03");
            when 19910573 => data <= (x"d571cca1fa2238b6", x"3e914701bdddce2f", x"a409a95a68e914ab", x"bc529bc89854ef5c", x"bba4fe97c5d0206b", x"38c19b94c2386ac2", x"294aa2b6d6173f74", x"0330f785618cd927");
            when 12779902 => data <= (x"7af3475ae8de16db", x"c240c2f00fa402a6", x"f270ed8f95b1af07", x"7ae8dd18f61ee958", x"194495ace2ea2a7a", x"74c3d138241fbaf2", x"c1fcb2b6d951f5dc", x"0ed925a15a88f468");
            when 25599394 => data <= (x"9ed2033cf3c1d19c", x"71299e2d77c672b0", x"a3febbcc7254c06a", x"9e7e8cc783f9861b", x"08c70c2e24941e3b", x"08a6c56561ba05cb", x"e4dc2304da698ffd", x"954dd217e0024309");
            when 33512159 => data <= (x"f147f823eb599f4c", x"e83bdd19a02bd5eb", x"aa4ad6e374df0030", x"b9250ff62a99a46f", x"c25b4b7499f4ade6", x"9975813b64c4c788", x"ecec721e88a517ac", x"c1af84ea0abe5828");
            when 13124041 => data <= (x"f6128a484eb291f9", x"4550c93f46ee8057", x"8c0c9f7af24f2767", x"40059c445543209e", x"ab98f46781d30615", x"f72d328aad684c7e", x"57204829b19a5fcd", x"56160432faca15d8");
            when 28799780 => data <= (x"c0481a9d936ee3d6", x"2562857c0b22ed28", x"1355d3d3de3a9fc5", x"1b386f3cfb5e1e62", x"3e0c3887f7ff5452", x"f0815f4565fec5ea", x"acbe2207a37c4767", x"216f65c7e98c0362");
            when 4740505 => data <= (x"f12494c7975692a9", x"e59ebee161bea5ea", x"ef2eb0bb102e4800", x"7ca02ad2e8052991", x"6ad90f0a2c835389", x"32088a5d413586f9", x"1c300eb41009ae0e", x"485e0e7660d07a6f");
            when 4782733 => data <= (x"eb4442783048ab82", x"5d33209aac0d5088", x"1737f343262bd193", x"dca2c586ec5bcda3", x"2f4796d8f892106b", x"614c053956965fdd", x"6ffe4fcec93b629c", x"39215d377947b957");
            when 15512377 => data <= (x"02666bffbf7104a2", x"5f471faf0db482f6", x"6a4f53a1cabcbf91", x"f4271ecc516e91c4", x"885994c7c36e79c2", x"6474590488c7043d", x"974b9b34612b9bf2", x"6276878c50acbeb6");
            when 12284340 => data <= (x"fd739f2a465d911b", x"3ac795be2b6972da", x"79b439637069ba3f", x"946753781b696e9b", x"2e05cba76f979d45", x"522123cfdedae0a4", x"05018af36b79b91d", x"c8911cd2f23fe6a4");
            when 24268432 => data <= (x"0e307b8e7954c26d", x"8a57f6aff29afa4e", x"99101c3cfdebea16", x"88400128eb62165c", x"1fdbe416116b498c", x"0c4a45fbb302c4db", x"48283a45ade8f03d", x"98d00cf338495dbb");
            when 31861040 => data <= (x"3723b2c689deead9", x"69157253c7c792c8", x"24529652cab7743e", x"40a2498946686cb5", x"1d9fa30731dc6b1a", x"41aef3c4cf87d25b", x"d32d60ef98e35c3b", x"a34a2ac6ff22821b");
            when 12326825 => data <= (x"982450e04d076660", x"ae3ac38145f4d145", x"cd8d59e268d10ca6", x"5dd4d67232a39a7c", x"8379a3a2d172f0e8", x"fc6c536eba7fc73f", x"7607e254cc1296c2", x"a943ae99293c4866");
            when 4383518 => data <= (x"cde3997c788da698", x"b9b8bc8078b0dbef", x"79fbd8d52110fba3", x"30814e924233e98a", x"375b07bd36644e57", x"4213607c7fca0434", x"a3e4aed9617eb722", x"0c3132fcd93eb520");
            when 18815310 => data <= (x"7cdb7da7a9561797", x"0c107afa49539674", x"b4838931c07bfc66", x"dca8b30c5b60b353", x"313d01993003d1fe", x"323d5aab53bab468", x"051ced901451a0d0", x"c7de52022a99d232");
            when 7162494 => data <= (x"4043a175983c207c", x"44a89c84d4797ac0", x"00428a9c72ff314f", x"d7f4cfa0fa38452b", x"91067bc4331292fa", x"e3a19323c3088c3a", x"d630f02027dcb67c", x"730b32de4e6a2d53");
            when 5620685 => data <= (x"78141bb24a691611", x"0bde2b90ce08b1e5", x"8db361033742a487", x"e8bb6dcba070e925", x"5ad324bd6f5dc1dc", x"fc8c00c149a22fa2", x"337c5eb843eb2032", x"e1d920a66343d6c2");
            when 23693687 => data <= (x"86a743492cce8d14", x"9ba920780c06554b", x"225508a582c2477b", x"3ce733e2e7fa4af6", x"d4243c5306ef2c0c", x"c2742ddd157f11ae", x"79a889b5d155375d", x"d5a9c3cc5de35f74");
            when 20064704 => data <= (x"84a578afb3c967d4", x"09b4de9f2d68ca27", x"270700b06a1fe00e", x"4ae8439e1354c6ad", x"ccc4c3b23aebadba", x"d9b13d62da7331b1", x"30ff7cfd613a9820", x"d9a1cca56608e293");
            when 32277081 => data <= (x"3687e906514a236d", x"7c688a28f718c502", x"f581fd714211e5ea", x"63ec767345967162", x"85cba57c14d3b4a9", x"bd3710e22710002d", x"85b3734663d49118", x"954d2c5997b3854b");
            when 4975841 => data <= (x"3414fc668b178ffd", x"8b288928226d35e4", x"3e7d3557d5b40413", x"d224ade02fdb05dd", x"d89d761bb1e488d0", x"9aef09b496a2f205", x"074c640982fc09d9", x"3305a2d39b203699");
            when 10254710 => data <= (x"707621984da45dfe", x"70ac339e4102ca75", x"ee240e4b1064c4b7", x"e1c21add9a4988d1", x"154752c4d874182c", x"97c5e640f65b170f", x"979b5272ca7b7c37", x"f835526dedc9c76d");
            when 26277840 => data <= (x"51186deca1d1eecf", x"a25dedd1aa2ac63c", x"11bda6cf1cb46091", x"a2d548607f0eccf7", x"71b9cb1f13d0e2b0", x"db4f9597f7cb6256", x"ad17d4dcb8422d8f", x"261465d66d44afe5");
            when 20191512 => data <= (x"166bff0983e3702b", x"6ac2f650ed3cd5a3", x"aa976ecd2139f96f", x"68b9c8fa0291a20c", x"521c367b562925a7", x"2e46131162e375a4", x"0db4c3c101c336a6", x"2b57ccfe1b307b1c");
            when 22418355 => data <= (x"33b4ce234e81d118", x"c6544062c437ce3b", x"ebfef7d2e3d32c48", x"cef77678bdf80c88", x"f5bd01f01b0c4656", x"c36284f378ec157e", x"9ef36131636dd40a", x"21f1f999f92c282d");
            when 15180832 => data <= (x"a38a654da954a710", x"9db1792f6ddcce2c", x"5cc3537e3d7c8c6d", x"1340aa0dcc9bd24e", x"819cdc3059219b55", x"1255f83e9278a300", x"03d59a9e848ac055", x"9753e1c475889969");
            when 5366703 => data <= (x"1645f447437d3970", x"fc10a260c97c346c", x"ea30acf31b9208f3", x"bb02cb17e2a99899", x"f1a6400c6fe6f30d", x"6c8dbdf4cf5dfa27", x"314a6f81c7c05a90", x"600f095b10584148");
            when 5626254 => data <= (x"c0cbb60e54dc2867", x"8fa9cbc35bbe41e5", x"994a97c7755688f0", x"77e3b3cca0640a20", x"b9d31871b3234a08", x"91d7c871ac5dd6c0", x"7e605cd095c619a5", x"81fdff9e6b032434");
            when 1328331 => data <= (x"57dddbaea6a120db", x"e5646abc899c4449", x"6b656a49b0a981d9", x"d8d09756a58f0f1f", x"80ac2159991a2ab4", x"5ab65791bd07814a", x"63c9c1ba9492fc52", x"3b850c85d9375a57");
            when 33911898 => data <= (x"7962f0bf0af563b3", x"4a838ba4872d95c6", x"549ebdb0b1d0a112", x"3b38d963cdfa8c71", x"4704b39129362909", x"270929d37480f970", x"0aceaed4e2c18d15", x"81882396720bf6cc");
            when 24239254 => data <= (x"b910936246f17698", x"943265db4eaeb765", x"ea5a4171983387b5", x"e763989208caaa6a", x"e2c384759d1479c1", x"d637374b443802c8", x"6613ffa02389e0b4", x"303def38195b7e8b");
            when 23175301 => data <= (x"8813c92f8f6726cc", x"e25c9c5d3900305f", x"0e82805836cd1fbb", x"07254df1f7d869a6", x"dc05b2dcbb5404f2", x"eb9c2f045e90d564", x"c6f788812016dd06", x"c5e780d3284cfe3b");
            when 10948442 => data <= (x"6d63a0459422cdb1", x"6029c83cab5f84f4", x"f04fe8689eb6a0dc", x"757295c27e5955a9", x"f375a7f80af26094", x"2c6de5bd8ed8227f", x"f578cf23fd65bccf", x"76878af6e47733cf");
            when 22010011 => data <= (x"b243579116e7f2b2", x"d29ece2a99eacb2c", x"c386704b446a0a1b", x"c6dd7cfc89e389d7", x"c2e758d562026bf7", x"6988335036902769", x"fda34082ace573b2", x"cdbafbbc9d9f5df6");
            when 3785324 => data <= (x"36359307ad69c42d", x"f57bf6b2bbd74ba2", x"d11b5171c5d38df3", x"c68de76fbbce5121", x"b9ca63423310b3cf", x"19693d69f9151296", x"3c5ed6109e13285b", x"c7da6ed4c293ecb0");
            when 30413279 => data <= (x"136082b104e07da6", x"d62ef9ce03eadbb1", x"2b826da74b0068fc", x"9c6b929b5853e8a4", x"368fc4e3bb336cc9", x"7496a4abc225ec46", x"7c8a2dc49a66946c", x"9822ac7ea391a787");
            when 19933879 => data <= (x"9675ea678874b400", x"a2e64f87c88ad98c", x"b29cb69dfac382e9", x"21c87165fb677a50", x"fccef2505f14a72b", x"6de9fbccd8818807", x"499d7b67811ac081", x"814c294da12b9a1d");
            when 5806629 => data <= (x"8de720a45e68d92f", x"5e66430e345c1fc5", x"51b3cb44b4ba8e07", x"9da940b7f2c766a6", x"838b11a0ba45ad39", x"f8afde091cae45f7", x"f24a363380745fbb", x"eda579fabbb9b913");
            when 2058109 => data <= (x"d02097b5de1c3db2", x"70affe37b46eef5b", x"257b4bcd505dc6c2", x"23b1c2e5b4d9b861", x"6fb3b16fd931a147", x"fcab7132babba072", x"8f7214baf5af0564", x"586242ed075ec47a");
            when 19569675 => data <= (x"36a86dc3e1723b4f", x"00a3abeb7c453f2f", x"608126b82c47f79e", x"dfacf794fc188fc1", x"e59b0dec79e83dbb", x"64424fed1ce78d37", x"b73f522241cc8573", x"db864ce4ba3f6bda");
            when 20138374 => data <= (x"8280f71373af66c5", x"cdbb1057b6b8ad28", x"7bb59746afdad103", x"12aa7402430da7d0", x"f9fd802f36674d0c", x"4b4d3578505f33e1", x"ce8e85be2960dd75", x"c4a3d47cedfeada8");
            when 16029004 => data <= (x"d108484f6ec83d8f", x"237f2363cc60fa80", x"5211a3fe9f188732", x"7e94ec055ac5bf9f", x"70245d4958140838", x"f6d50f9549cbf508", x"f112619a7cf6f19c", x"8f79ba9a5f70d196");
            when 20817410 => data <= (x"9a3eb62750cb164c", x"eb87e840f47c8945", x"410a0748eeacd918", x"cc1e7b5d195a22f9", x"0af650d8c7a1f90f", x"77e5e6e714d31a27", x"9f3aa3018e827869", x"520c70b9fc55b915");
            when 7204642 => data <= (x"eb43d95214f72a94", x"fa93391996ff0662", x"6f124804559fe525", x"ed3c8d941a337329", x"f9b01b6dcbb761a7", x"16425a7c4ed96105", x"c0d443613dc5017c", x"33d1935c4c097d75");
            when 23876328 => data <= (x"3776db0870245dc2", x"be0a6c855542a247", x"4cbe9b3421cd8373", x"ccfd59e19ec5893f", x"c7ba880cc2739886", x"dec084958a249400", x"20e896330e610fda", x"d1c52c98671c07d4");
            when 7169609 => data <= (x"8a9a65a143fb877f", x"b31947c3afa8389b", x"20509de465028096", x"7b08d0a5d70b911b", x"d6f95b4b4bfea159", x"2a4233230921b6a1", x"51fae098bf1c0056", x"6bcdcfba5c2db93d");
            when 11932496 => data <= (x"313a3c51861cfdf6", x"1a9e3d1ed2f01101", x"d6cb18080428ee69", x"9ed617e60d69eb59", x"dcb2b1d4795ee287", x"8f037b4024e9acb2", x"941a55dad2665493", x"87f2e3d616d64af3");
            when 7613127 => data <= (x"b19b9231d511e8d5", x"c6328e2cdc92a528", x"4d00f9b1ad823ac2", x"f76dab50b7e2c5d8", x"0aece130f5800524", x"8d8637290b9500c3", x"20bb9cd9749b09f1", x"b84410822fe14944");
            when 31203718 => data <= (x"d0d7e547660ee606", x"ed62094409778f0d", x"c500cd2e39ca9211", x"24335a3e0028e000", x"9ee42957c800f271", x"ead0c3921c1060fd", x"103fb9a55a9ea71e", x"e78131929f704fc3");
            when 15759311 => data <= (x"975dae126b645625", x"70f97546e4be82ac", x"888d083c4ea5edf4", x"2cdee3a71dd61295", x"65b3f9843a3f8e5b", x"bab51e64f73f7f8b", x"7162707901960c58", x"c831e76b01c3ef1b");
            when 24394909 => data <= (x"7628cdb05ea7ead7", x"8c74beb7dd2319d2", x"a97e684372004e16", x"1a0f4b5e7e31552f", x"6a03ae0f097d6820", x"b4e71b4b17dc9e55", x"3eb1cc61d92294bb", x"cd80c28ef1bcc436");
            when 2603384 => data <= (x"7a2428224200f2d7", x"d0fdc81aa91f65ed", x"2bcbd37b7db4dbc0", x"169a32ef9f5f637b", x"d58bd1279542a0ce", x"bf8e069e584795a3", x"485a2032684780e2", x"6d0a519ddb0084de");
            when 18340900 => data <= (x"c43d2bd9a3e724b5", x"371b9b2f90e32481", x"d713b0ec2496fd54", x"4059c7caabfc6caa", x"452fdd179b1ec903", x"8f3e8497dff2e52d", x"e9a201748afabbe9", x"313a543972929aae");
            when 32958070 => data <= (x"83508555f3741fe6", x"b536f3679e6510ce", x"05627fa49ba9cb0e", x"cd3cf1bb71bbc297", x"0a90a2f1005f1059", x"6b4feed637c794aa", x"86cb6950327257e7", x"a16293d3be244c41");
            when 29530635 => data <= (x"44258f98290ce2e4", x"bc38e6e92ff737ff", x"9dbba675990e6f20", x"bf071f5be5e2b132", x"55d2dfe8ef7c969a", x"aca50f780ca2cff8", x"00d678db7da6995e", x"cd4922cf36a26865");
            when 23111645 => data <= (x"4d1c891ba82e5ddc", x"888722a3aedb38e7", x"3a9c8cf269bbad4b", x"de7ee301433a8765", x"59e4df891e326c8e", x"c2d6e35dc9e6ea64", x"fb01ce53749a1f8a", x"7d5e31b1252f5a96");
            when 25231317 => data <= (x"95114bbd7011a60f", x"52e65ba15a873886", x"399658354b8a0a41", x"9675ee775263d685", x"498ceff8456ff457", x"560451a2535661ac", x"bf3e56f34863baa6", x"aa65684ddea5e5ca");
            when 26559449 => data <= (x"f6b748acb78e9990", x"60e385cc0f918d02", x"94956752c1e9fb81", x"05c179564cb0b35f", x"5a677397c87ec4e3", x"2bda55f6f4569a39", x"4aab4f0d53b4ea10", x"fd6f1ec2129c9621");
            when 13902274 => data <= (x"9f1c1d5eea80a9bd", x"a39f3778840b6185", x"c56bf7a10c7293de", x"864d656593b3eb7b", x"a4602e7e1cbf12b5", x"787e867e65a1fc9c", x"ade7ca3f18459b6e", x"e25c0549377f1a5a");
            when 986854 => data <= (x"a67513283d689eab", x"7b08673fd5205f05", x"6fbc7b53674e2121", x"ff05bfd5526e4d73", x"8a03f7eb6db43d80", x"388ecf81ac060d74", x"bc2d47cc63a9dca2", x"c09cbb79747be079");
            when 21910450 => data <= (x"357ff259f0a2931f", x"585cb25d8421dcbc", x"a3f0d3a0f23b0093", x"87e2a2f8063470c2", x"9e1d227a0c5f11c6", x"0d052780c878845d", x"1a76a0198292736d", x"c90fa72b56fc9982");
            when 13771815 => data <= (x"c6ab10b656982b8b", x"3697e1e5b421388c", x"02c507b39acf1821", x"ce94d3a435f66ed7", x"bc82fe61a69cf071", x"194f7cb686a56d2f", x"6d2360b4d4b5508c", x"0d8ee1acb06eea31");
            when 26897305 => data <= (x"cd85fbaef320d321", x"ed3d11023560f61a", x"788add41d48f49d2", x"c65dd89c61bd73bb", x"96313f257fa48027", x"211f18f85719f80c", x"4d0aa20bda0dd6f1", x"814523296cba77fa");
            when 15640695 => data <= (x"b9f9be6bb0fd8503", x"db774a95942c51b4", x"45828ed3f4f27ef8", x"a8f749b0efa9fc29", x"d3a928868fb7f341", x"69024f151b4bb24c", x"74aeba925bd8a6b3", x"fbb4d9c6b8b0246f");
            when 31103371 => data <= (x"93e88a96e9061a4e", x"0fea6868026bf4c7", x"302d19ed60142776", x"8615eac9d82dd986", x"2921312145bc23b8", x"91527acc8bea074a", x"cd61f9bafb55f074", x"5f668634725cf211");
            when 17918383 => data <= (x"0bf4e8b9ddc23e36", x"1d86449a3beac4db", x"6701252c28bc5b92", x"303d83fa2199a5e1", x"fdbe78f2b38e286f", x"0cf7a2cbd646fd64", x"f1616704b5f0c9a5", x"8bad1b19f81198dd");
            when 27460113 => data <= (x"69aafde7d5f508e4", x"442d520bdf448a12", x"c86cae09371feeab", x"5e9494cf1b88ac22", x"3b93e06dcef2a8c1", x"053f41aeedbf74ba", x"e9cdf3c32df6950e", x"dc52f20c30332f2c");
            when 13878656 => data <= (x"3a4fae32422bf9a3", x"9235f8fb75f5b74e", x"1a371b6b7a16baa1", x"bdb85d5104987d53", x"fb8242086f252d89", x"0a64acba720d59fc", x"bf93b144e00c9fe7", x"3fee9cea266693de");
            when 16095424 => data <= (x"ad9253908e5f33e2", x"24f4fb8574877c6e", x"80a908aedd754fe9", x"8d5ed550d173c844", x"f618deaf1ca65b14", x"732a01bdeba45bf9", x"4d69dbdd123b15bb", x"73eac732e25042b1");
            when 27015309 => data <= (x"8a72396009e49c90", x"4c3911d195fb2b3e", x"bf6deda0ddf7a9d2", x"d272b0a06f07572c", x"9e9c441d6a5b7185", x"81afed7a642c318a", x"e8296551f2fc8e6b", x"ca9f1148b5b93586");
            when 14405745 => data <= (x"916a137a4535af74", x"ea4f030668b7536c", x"3c1ce4786fa58f1d", x"26b6ef10d396627e", x"b1570a21c3ee90dd", x"96469438d6bfa8b9", x"98173de28f3ece59", x"833a728ffd9a6213");
            when 21035281 => data <= (x"e836bde31b07ef59", x"e64a61955db0535c", x"2ef79b9be7e65d02", x"761ed1b2e7afe3ca", x"c13466d99095a3ec", x"c4715766478f8a28", x"08458ef5a94947ce", x"da52419848eb432a");
            when 11069245 => data <= (x"856f24bca6cfd697", x"0e34fd770b800e13", x"1950d5f01e967a0c", x"920aa1c38aa8c49a", x"4c5037195c10e4be", x"319d71f9c3b2b61b", x"e590e92bcbe6bf6a", x"da6f4abc80405559");
            when 16933030 => data <= (x"a92455171a0e46ac", x"e5e4cb34fd5e8ef2", x"aa21b5643148719e", x"8a7a3fa7115a7b8e", x"702abee603b61bd3", x"82e99359388da566", x"7e9d12e854bc9fda", x"2db06db2fe0c872c");
            when 24940995 => data <= (x"2f03d9f4d14767b5", x"cb0904b1606979a7", x"a4b9a3fd80144d37", x"fcefd827b028431b", x"739c754d5e9a9a7c", x"87980459c8225f1c", x"99d692124720f1ba", x"255e644fd49fd287");
            when 3833212 => data <= (x"576c7060529cd78f", x"6522e88a6aa422c6", x"68ff02788ba4c899", x"958369afa35a0632", x"ff9e448bcfec2616", x"707e4d5ef3e29dca", x"6db48908e9207d97", x"e845bfda65f5920d");
            when 21939950 => data <= (x"044f563250d2563d", x"6cab069f91df6639", x"8bdb29124bdb5b6e", x"33307092f2951006", x"aee9acce2f6cf2f8", x"3f922459ef4fc4f8", x"d940d09c0b7becd7", x"f2f199a0a67f2cda");
            when 29356376 => data <= (x"d221f554321dbaee", x"dcc8a69c81d75e34", x"2b40f2c2d303a87e", x"771cf78516476fa3", x"96f46fe6e7c9e47a", x"a12a78d52b474eda", x"ace1a3a1037ea8cf", x"5f0e15c6f8eae51b");
            when 1593151 => data <= (x"2f55a32e5d2aacea", x"9a6b71e4ddd2635e", x"dc96be5ec88af99a", x"705edf7ed2e8b8a2", x"ce2038440c03302a", x"2e9e3675f0f0a45f", x"c4c0235c8e929eee", x"0aa39e3890c9a58b");
            when 1218164 => data <= (x"d734ec2d34d4281d", x"7b6a836d7937dd8a", x"e77675ddb57082fc", x"fd16cb1315db0352", x"3632a01d3c62ace2", x"a442c604d574f277", x"a8b254bc9dad53a3", x"de49e71ab623b052");
            when 27533705 => data <= (x"8fa1576cffffe4bb", x"1d06ad986d84ab51", x"e5f8293cb15a9fc3", x"65181a04526f2889", x"9e1aa713a066f7d4", x"abdc6fcab30be4a3", x"288fd434e0645366", x"4268760f8f8e0025");
            when 32458169 => data <= (x"dbdbf5c05de8b644", x"5d66fef36e93893a", x"a710a8aec3626449", x"b48a14ff94ab685b", x"1cc2dc6ce3e8f026", x"0afe5e95e39edb15", x"9a8b76572f5ffede", x"8866a8701cc7fc1a");
            when 20282992 => data <= (x"b8fc993e45d9e9e9", x"da1be682f7cdbaab", x"ac11abf7461cb603", x"cedfffc787d65675", x"a6b441a852e92256", x"dc533696c96ee2c5", x"7a52e686767b8f1c", x"08581b236e5a2f53");
            when 28380056 => data <= (x"8000ae4f5a4e2adb", x"f6c0630270bdad93", x"cda2aafd06f46c98", x"605b9c8c39a1f579", x"3f87ba7a022f6ebf", x"cf3e8cfdfa23261e", x"0dfaf8c93fd6f9b7", x"0b4bdb9e9e22b73c");
            when 33501274 => data <= (x"3dfca3bc48830122", x"fd8221aa7b25b1e1", x"544e0562803cc96c", x"6866ab4bf753e604", x"a829b28e83afe198", x"7f154e940fc40b92", x"d18579ac8c870418", x"ff3920f83ede6bb7");
            when 20479494 => data <= (x"2906b53db41e97c5", x"2ef67c15f3aca29b", x"aed99ad7c0b98e27", x"8ba513ffe2b0c962", x"8cbed334cfb0b3a9", x"cfd4f739ffdc07b5", x"943ef71e596f2fd5", x"b2d7324e24f496cc");
            when 4374171 => data <= (x"af7c867e2fefbd9c", x"e0a71f0696bae8b2", x"ffbd76b24caba8ce", x"fd0c64ebeb9c1e18", x"841a2bc55b8ae244", x"560593b5e72cb4de", x"e11b93a7a62dddc7", x"2cd67045cd79e13c");
            when 17183063 => data <= (x"f0eac9ae6f7e881e", x"85851a261e38f4f0", x"c167b990ea17b954", x"fcd3d1db259dfa64", x"06f40eae7e1a90e3", x"dd09083ac30a4439", x"94e7efc88273365a", x"eccebcc5119b6ad2");
            when 5760656 => data <= (x"5232afa1818f09d1", x"3d0844febdd097e3", x"e4633fe03ad8781d", x"a517798922afde0e", x"759dbc759254ca47", x"80352443f4b0ed32", x"c195852b2616967f", x"389861ba8f72b173");
            when 22646499 => data <= (x"3f1527d6b0deb43e", x"9088161cb1ec597b", x"28cc1b38b9a744d2", x"26ae25bf770134f5", x"9b16a082db5adddf", x"a03b19848bd14835", x"86466d79f5e66693", x"fc7d816f9b88628c");
            when 2827617 => data <= (x"b4dc5897cc7b704d", x"358154227050da62", x"3a49fffdcc04f775", x"0fb943f81ccfff33", x"f851fd13bd173c15", x"e4b2fe62677196c6", x"4ece33819c821533", x"62ee176d43564182");
            when 19010594 => data <= (x"14ab7d082bbe1910", x"00c7e1feabbc93d6", x"5fb7b4730576cd8f", x"e09ae71a56a93ed7", x"249b782677bf55af", x"cfeda2b85442e09c", x"55f062498a5b4b19", x"d2fa06c12101168b");
            when 27738493 => data <= (x"829516a94a98c44f", x"ffa73f1a87fb85bf", x"9e4c4fd3b3c77a3f", x"d7a7516293742aa0", x"be8ca2c484585f6f", x"ccdbd8b0722d9b8d", x"7e04e194f39a96ce", x"cfbfb980b2770516");
            when 13506823 => data <= (x"6bf11bab94001862", x"054b22ee788d2041", x"f92763a67c319d69", x"3cdd44011ba275fe", x"d626711aafd5bd13", x"4d006efa5fc4cc7f", x"965ca17530089417", x"061e98314bbd4228");
            when 22678552 => data <= (x"6dad3c00b3b9be3b", x"3f35130b5705fde3", x"51c5712ab7fa5494", x"820bddffa76e0abb", x"833d3cde38542cc3", x"32fd3b2b8c82bc02", x"3f2f4abe7fb35158", x"c1d905456d240c1a");
            when 6076020 => data <= (x"2a1f28fba13dc42c", x"a85b1b52af5b17cb", x"5a546fa9f4972f4a", x"b7aa90ca7d787a2e", x"2c9e8f92d8c5d4a6", x"db53d5c1bab7889d", x"de818fb929e79329", x"a25f7e6ad719f017");
            when 13891454 => data <= (x"c775d5fd3c3287b4", x"652fdce25f5f5d14", x"cf09fb48bf2f9f83", x"342e7a734b9a8136", x"c86b6f978ac6db6e", x"1933278a98323ae2", x"72674746625bcfdc", x"a1e7599268e7981a");
            when 4683158 => data <= (x"681771ed93be7592", x"1706c0ef37b6055a", x"16a1923e2b4e1304", x"cb1dd4f6d7d33763", x"c61fc74179e5ae42", x"212e9fd69ce61baf", x"127aa4cb073d4cf3", x"ca8f188a6f52fed2");
            when 2569668 => data <= (x"1fa1a65700167358", x"3507599153925f13", x"67becfe30e8c08e0", x"5397728f1b7aed3a", x"752284686e3b2a69", x"eb5683cbe51a8c05", x"737446e08b85ec73", x"0d8e55222728da2f");
            when 5460667 => data <= (x"4fdbc69a8ebf48cf", x"4c40694d7931eee0", x"bbd4d46d7859a77a", x"fd109fdfa0a55de7", x"10a70de0831992b4", x"2e4df7ac9c2ecc61", x"f587b8f3b4140c2d", x"38088fd9ad7b3aac");
            when 17010987 => data <= (x"72ed58eb7270e9bb", x"8f86d2f8c46c7c25", x"acacc6c419709238", x"8b773ea858d6b5e0", x"503f59f17c75219e", x"2b863fd8ff8cf992", x"590e0cd71181550e", x"37bd0136d4b7780e");
            when 6595712 => data <= (x"2d19e9dbb4ba6f5f", x"a8f53bc921edddf0", x"8d555522519eae37", x"c28ac850ceed2834", x"31ebf56d339a7f1d", x"d08b11ae3559ea8f", x"9ce487d979083458", x"5743bc8d60374291");
            when 21246521 => data <= (x"20f9bc6feebc513f", x"12ab1d7f967faafd", x"dc87255260f9878d", x"b5cf9558e1bf39d4", x"22ed17cb40bc7984", x"5536ef42257efe2e", x"cbd64f7ca5ba48bf", x"0414b22cd0e45d53");
            when 30592952 => data <= (x"82114e1faf894d00", x"1bdc21fc32685e6d", x"3b722a8ef00f8bdd", x"f5d80408281ce3f3", x"4bc6171b9e941e29", x"9a955af2011d3a86", x"0656e84bd094d55c", x"95c2b76ee213cea9");
            when 5908036 => data <= (x"6b0298aa4cd577c6", x"9ee676bdc47d86d4", x"9ab246bb1a3fc186", x"cc91e2419e36f3a3", x"9b938eda37bcbbbd", x"4c8895964f4c921e", x"645d88a54a97f6fa", x"a13e76a13d35e6b7");
            when 31649165 => data <= (x"3fd03ccebedf9d52", x"85f8071e4aec9a8f", x"362a2378185aeb57", x"066c53ce34860cde", x"8714dfdb21c59847", x"0c333a77ea88a8bd", x"1de965d07eb25a09", x"8dc34f3b5e3017d8");
            when 20861522 => data <= (x"a68f03d3723291a9", x"dd3d5ec8e7243e28", x"48922e285cb1653a", x"394b0c55fbd27d80", x"df6bba15ae424155", x"11a0482da5aa895e", x"df29916c96d73470", x"c6a8a8ec82a39a53");
            when 3734749 => data <= (x"d290f06e3d5df008", x"ad0a36105e1888c5", x"d6847ffecc9359a9", x"dd9766b99f5754a3", x"0545545e116d17d0", x"2e63cc95834fb86f", x"5c942d632a7dc8e3", x"60947a25261c8e57");
            when 11305506 => data <= (x"d40374fe42aae25f", x"6eb125dafb86e864", x"2dc71b638dadbfbe", x"0c4a8d67438fb91d", x"ba9524129188e931", x"9553d0d86dcace44", x"64de003cc1914171", x"414772b6c7c63381");
            when 18182879 => data <= (x"941d572a2b9ec167", x"963edab4c4ad066a", x"398c980924a507ca", x"05a32af93426ea04", x"7b3837ef98dd41f0", x"ce0220a5dcff57e6", x"a285e84e3070db01", x"4c511023a5aa347a");
            when 29563094 => data <= (x"1878b03f6e2bacb6", x"0156bad8c564fd33", x"ade67c2d15361426", x"fe655faadd355ee0", x"04eb8bee755b357a", x"c526ad604deaf0a9", x"16e347a0f4c80f8b", x"c8606fc06a951e0d");
            when 11196508 => data <= (x"1545633c0b8bde49", x"d2c33ac34f72689f", x"6f2eb8d1becb70ae", x"0a0c7d592f7d1542", x"29829d29048f3f1b", x"daa6895db02e2a52", x"6946d3d7a0eddb50", x"0bb057d56f0131f5");
            when 22169532 => data <= (x"c927da59fc1a2444", x"f1400d2e7d5293c5", x"1c3c41196d9e3313", x"b5023e8600a8c22b", x"03be977036dc52b9", x"40d29420af7dfe1e", x"537979a5bf966383", x"e59d3d86025a02a9");
            when 10236971 => data <= (x"85fb7b445d00078e", x"e05763e5d52fc4db", x"947159aaf7cc1561", x"a390dd9336422026", x"6e89499beea92b6c", x"a99599491c35cb30", x"c1239292c7c76f65", x"894748c742c10d44");
            when 21690524 => data <= (x"61a2da62caaebd18", x"801c8c4fa548b66c", x"f01391343b969003", x"b08c57a8694d73cc", x"3c50a19e4e865e2f", x"2ee0203632210032", x"2fa00b9f5f7be1b2", x"0c910c1a8c650e80");
            when 29473689 => data <= (x"d57ba6efce1786bf", x"38e5d0f561a784c3", x"0ed1fd7e3a40fea0", x"90deaff8036633e7", x"0744b7fb5027ce48", x"3d18eb3e5f15257c", x"7bfad00fcb9a962f", x"8953845338b77797");
            when 959133 => data <= (x"9b8c8fb90e3552d9", x"2e5e01520d9007e5", x"574ec45f9d1f0611", x"2996a4ae9732e51b", x"e71a0f21723f28d6", x"d44e7316c7cb2781", x"715ff5b7eccf7120", x"729b98cfbfd6853d");
            when 24861946 => data <= (x"00927b07125e2aca", x"3a3fea6fad23d706", x"67e69ac46eeb0488", x"8607d6fefcbb56df", x"985e07616a6424ed", x"ea46d971104f0912", x"3883d47262485ccf", x"b89b33a2fa1b2286");
            when 33948465 => data <= (x"4c3b1dc19e0360e6", x"bb51933d7065b801", x"48888964e97eb39f", x"d4fd2f4d0a716229", x"583e848f51ead036", x"b8012a4dcdcc170e", x"9fdd4655a3da179b", x"8f32aca8fc6f58fa");
            when 18739081 => data <= (x"198d0a46e10e62d5", x"5460ad8a38026bc1", x"19296aeb4f606376", x"4f50b7cff0c8b7fd", x"4397c7d05b8bfabc", x"fe35b673499d2fba", x"fb2a453f57c5548f", x"8369695a866eecf6");
            when 6628057 => data <= (x"5504fbdcc66463ff", x"e546578a704a5710", x"0814eb84dc26188e", x"41e874b96383741a", x"2d8929ff0ecbd5c1", x"1ad1daf5f32360cb", x"fe07fe2aff432fe3", x"18543f16b4cc9eb6");
            when 13916750 => data <= (x"93445de7edbc0c5a", x"f808fb6030154059", x"60de7548d95687e2", x"60e6c7ff09a14736", x"11849093557f60ab", x"3ef62ee3e19932f0", x"89e137fbe364c5b2", x"fa25f9ed6b69de34");
            when 32221547 => data <= (x"c66f1dcc6b5b6591", x"1c73bb7e7f424540", x"b4f51a7e22bf04b4", x"6219a3e45c952633", x"750664a181aea671", x"c84a632933b72dfc", x"2f95b9930fd3a5af", x"63d2a1bb39506355");
            when 29493066 => data <= (x"abd4b8067b0e5381", x"3b12e89a5a8bbb0b", x"016d5bc3140e6424", x"a30d22f65c4d1f0e", x"1713572ced52e303", x"f6cb1811005251c1", x"b87214cbcaa9d12c", x"3c000b306bd9b6f6");
            when 12100164 => data <= (x"3d4140d882238f64", x"e3159199163821e0", x"dbc88b206128005f", x"b0e9a40722c544d1", x"986ba5fbff006478", x"059fb2c8487f7f70", x"b1d9767b2ee9164c", x"74c756f2bda9261a");
            when 29267473 => data <= (x"987addff01cc4f34", x"853d43305b977a23", x"321205aa93289438", x"261c4174ae4583a7", x"13f1a13e0d641f79", x"dced0054f45c5970", x"e87c441c1746f96b", x"4f5df49dee610d27");
            when 3256671 => data <= (x"d3ee717f35f16f47", x"21dd17c43ea8cf90", x"2b20031c9d3dfbcb", x"7348d426ec8fa587", x"41b8a93380e97eed", x"5cc26a8b4de625d9", x"c551e72a7b074113", x"5dc7fcfef7a6a258");
            when 2485423 => data <= (x"d84cb533189b75f1", x"40f25cef9f4ef545", x"fcd45be7a9e0240c", x"6793761f5b13dc2e", x"06cad01da975f2fb", x"9843e2080005936c", x"989f015d1e992982", x"99f5ad0769e39e16");
            when 33486486 => data <= (x"991fdafd284ca062", x"0f1e613786ab0e95", x"3ebbeffb71dd0464", x"24e88ef87f062144", x"3932868c133929dd", x"54556c091074aacf", x"51bf4578b4e9c60c", x"8125db0ca70eff25");
            when 1866409 => data <= (x"bdb15aba8e4dfce7", x"91f9804fa87529eb", x"eef7d92982d5509c", x"1fb2cc1909b75c2c", x"60d16e3cbbf0ba36", x"b3d7ad2f7206345f", x"98a797ff3b2a8c50", x"f996fdc593c83466");
            when 10983750 => data <= (x"54bc404112c700d5", x"662fd78f1d1f637f", x"ea4f3c193249a58f", x"8f1b2bfdcdd14e8b", x"8474c4ecaf48d2f5", x"d213128d0c15ef19", x"a18c640e3534cb28", x"035ce8e026ee5080");
            when 27472094 => data <= (x"54fdbf7c8daec11e", x"ee7e7dacf1c14307", x"9ae302f185e2868b", x"d160e71fdef8b57f", x"acb1c378a4c17cb2", x"a41bc8ea6def53e9", x"a667131562cd36eb", x"8a73c183ce724cd8");
            when 6122152 => data <= (x"3cc7290f5c3f04d2", x"1c508b85d1cc5294", x"c0f08ad17e2a9191", x"c0cb3f900a5a2f34", x"413841d25620f8df", x"22b8f6cd442c5994", x"fa4f4daf32ec0571", x"cefa79489c75d6bb");
            when 5159242 => data <= (x"cce8f38f84aae660", x"aa9ad708967899f0", x"239da54536088753", x"79f61773a7fd2dd4", x"3e0b1678358416af", x"36c13235245a1e6c", x"8a3072f643a0fd97", x"4386f20c98be89af");
            when 19503244 => data <= (x"85de236ba7beb7ad", x"16cce5eddf8b23e8", x"b05e39561d48175e", x"0526fd9560c1a812", x"a0f8d1430dc589b7", x"c3ee675dc4302736", x"312224d537630088", x"43605a8c102b2433");
            when 4119931 => data <= (x"f603eb9a8fa2a400", x"8917695003ab953e", x"d124e963ec9a1f38", x"9f0ec9f931bdac6a", x"0703a4ca86db591a", x"9451aeb9630e1c04", x"0ae7fd17e63f9c6b", x"4526fa9da77514f3");
            when 24868124 => data <= (x"810c65e5207b3801", x"86a2dda10bdaa678", x"b9a5f0bb6cd0e177", x"03adea242f2e0633", x"47590a4ea8576a37", x"e74ab166ef64e6d4", x"1d6628ed0246f51a", x"d93eb968c1203295");
            when 21851234 => data <= (x"8486f5257dd8745f", x"c33f732790f0072e", x"6600d543720e8152", x"bd2649a929bf3b76", x"93a13dfc780ed75c", x"4c45743c01093c58", x"aca6803570899fcc", x"4d63088e4bc0616b");
            when 4128752 => data <= (x"2898e3fe3f0d38c3", x"b278d3933115b2a3", x"29bc50d99becc99b", x"f71071926a780919", x"6b55abec7c242b32", x"b5bdd46082ed1f97", x"96328f44c126747b", x"e9076cb982d053af");
            when 14912631 => data <= (x"7b34bf25831e91de", x"a91d69f33c5d80e1", x"ccb2047e2ba7da3f", x"747535d40b7db698", x"f161f94b6dcbe800", x"3ea656a8bc25ed8e", x"9a3bab5be37061e5", x"813f8d17d769436e");
            when 29584576 => data <= (x"b5ab4566d7a7588f", x"f84034a719a56a49", x"3957d24b82e8aeca", x"3f026ec44417c29b", x"cf6ed1c8f246e8e2", x"ecd575747e2a53d7", x"530e901717ba91b4", x"c44304fc1692a9a1");
            when 21832975 => data <= (x"78f11cf4b017dd6a", x"b36c15567a18824c", x"31d3284a7f85552a", x"2e69d6678b229c71", x"be2f64dca2a92fb0", x"71370a5ce37b19ef", x"9aaf09b2693cf4a6", x"537f9d6685ccfce8");
            when 11490989 => data <= (x"3f0a437e5cd1b98e", x"be02328e390862f9", x"65177702f6d517ba", x"c7acc500336fa9d9", x"5d75b68f89d48064", x"cea80d456ce20ed0", x"f54efdd280a3a5b5", x"8bc123e4df9a38f2");
            when 13571025 => data <= (x"29026993d6217160", x"7ead78559606b8cd", x"da685a970c0dc8c1", x"b079684860a9965e", x"97a8443b30c2abe8", x"eaf54170ab402d9f", x"57d12ca0dcd81af8", x"d3f3ff11094d4de6");
            when 20615589 => data <= (x"9f851661a4f31007", x"e176bbd50154afa6", x"e210458768da7249", x"d270fb7d5c4b5827", x"394f5da245817a0b", x"84b87293113bfde4", x"84a607b89bbbb704", x"2c2df870228023c2");
            when 684546 => data <= (x"e9b1ce2fc45575cb", x"5ea8b0a6a26c97f8", x"00bb5f8ce870e9dd", x"8cfdf741b8072ea5", x"37f5a46bfd30d46d", x"b62acd895555391d", x"66954b2da84f98b8", x"828ae019d8029353");
            when 7422398 => data <= (x"2e8e680e30fa3d2d", x"b830391176860d30", x"9ccfd227dc29573e", x"f0394bac52d60ed0", x"b1c087f66bce8f89", x"b3680e13a4d13c3e", x"cbddb813685bdace", x"f5d0b4f7a9cde86f");
            when 30944631 => data <= (x"c64f91a1de5bcfd5", x"511d056dd64e1b94", x"fcd98eeef52d4222", x"30ebae6aef1e7648", x"67dfcfabc82388f6", x"7b4faf656b6384e8", x"9a7d6cd1779a22e1", x"e69c0cfe6a27981c");
            when 31277720 => data <= (x"98c602c98f352d43", x"9c7d9f29457fc709", x"1d0e06cb4c171f41", x"11418e9034d771ca", x"a547162001dd3b5f", x"5927617914fa44c0", x"3fa6235e0d95a21f", x"7d4b008d81e86277");
            when 1050790 => data <= (x"fa281b332137d48e", x"11b2691f012e9408", x"d298571dde3f873a", x"061051c805d20b97", x"4e683cebeaa1c8a5", x"ad84d69f1cb5a241", x"820b0ca21c8536c2", x"6de0d31d0501a2ac");
            when 33019604 => data <= (x"99785e2e05c0f272", x"2232f84d7d97ad66", x"e7373a3340eb7b39", x"87aab84821eba2e9", x"afaf21603133edaa", x"3efc28025b455f98", x"281089fddc9285b4", x"953da32ef1d90472");
            when 19000039 => data <= (x"93e0625fd364e273", x"1a992e68c6955bba", x"54190a977f2fb9e4", x"b8f034367f88fb7a", x"9a6aa31ebf7a89d6", x"97e0769e491495d1", x"badb8ddeb9d71706", x"8af55aa5764a0840");
            when 16741202 => data <= (x"bc9c6292a3cacc7b", x"1178b04d07360407", x"3b102ad7407e4860", x"fe4c6baf23d5dc15", x"3986741ba2f43b6a", x"bfafc0241c6e8940", x"8e4bcf9a1b0faea9", x"142c8ea6a4b17d1f");
            when 7447376 => data <= (x"cc6f0037f575f262", x"0e9dd2ae1b89e9e6", x"b026c147fe7da375", x"e74b3ca756aca48d", x"6b0aa66d2742df82", x"0489605d851c124f", x"076944dabbac6e19", x"851a6db91138e164");
            when 23758228 => data <= (x"4d437c4d82f673eb", x"07dd18e348600c11", x"82ccb99e7559e126", x"624e0003cb8731e2", x"dc941d967071cc18", x"6bfe481d2f55d1f9", x"06ece133652d6371", x"0b8bcdd337c11bf9");
            when 17949179 => data <= (x"5fb1cbd0dd667816", x"91b380d2908dcc39", x"a26b59639c23d07e", x"8dbcd95aa6180f04", x"556bab40b81b1842", x"f4b719fbe0e0747d", x"734604bb3fa51a72", x"1af2f239f54a3949");
            when 30658277 => data <= (x"a446c672a26e2141", x"c1a18c59a32680ab", x"3f1cdd085897d750", x"9b7abd20f6c5ee5e", x"9327526996d4d2cf", x"47f2e66f456ba21e", x"5825311a9f9ee75e", x"89c926b1f0dd650f");
            when 11982542 => data <= (x"93579e3384848996", x"f070b77f5f9bcab2", x"2129178215f88347", x"8293fa249cd7a936", x"2747201468b838fd", x"8ce16e1ddab568dd", x"ab4cfc6446487832", x"25de285fa14fa4d3");
            when 14703796 => data <= (x"339f8d844f95e09e", x"d4add84b1d4d1b17", x"ab0804847733d8de", x"a06295d53ba2ef8e", x"ff97b58f1f7dd081", x"328c644d8edcd1d6", x"9ffac19372aee662", x"70764a9e257eb50e");
            when 13194677 => data <= (x"d12025365b2a4701", x"14d5d053f763e570", x"f01ca19f6dc1296f", x"d876a81c4883ca0d", x"a19bafce7a900fb1", x"5df38ecb9ea4ce0c", x"c63ef8305beb4f7f", x"3c9a0cfe90f8e3c3");
            when 18594426 => data <= (x"1939811ebd8d886c", x"90afeb262ceb956a", x"3114b68c4574c218", x"45dec157cb4d1917", x"6fb6348e049fea65", x"7bd22072e9718efc", x"ef860ef450931122", x"b45c18807ca90b6c");
            when 32360945 => data <= (x"378bf4543979dc27", x"cde55db4c1195720", x"307a161f00a31281", x"8d4c77a4ac7bf01a", x"eff347a86c08bb35", x"1093e92e78cffc7e", x"b6ad17b41a05aea3", x"5e6ca6aa1b9408e5");
            when 13210918 => data <= (x"115832f8f536cef8", x"bad5824d039489cb", x"20eca37d45d80294", x"220dbfdac397cb86", x"c0cb04f01587f927", x"cee269edfa7460b1", x"71e3adad14b9e980", x"8eff56eaf1d5e630");
            when 963042 => data <= (x"cd4845d55618b1fd", x"d6c2e485d34f9779", x"125efc453f662011", x"f6e0608659341b7c", x"0392627f0f69ca99", x"b0de6529ff1b1e77", x"8ce5a93d56fa9298", x"b7c2396e1a4747c5");
            when 20478581 => data <= (x"508f7e78cd9e6505", x"912b4cf6dcc131f3", x"1b9fdd519dd1adc6", x"632dee6ed91119f8", x"483ebdf6666da28a", x"53f97192cd33111d", x"c4fe66678fda80bd", x"9234ce3d81d78e43");
            when 21825770 => data <= (x"89810a4708f4de33", x"4df735390d9ab25b", x"628510b69f197e59", x"59a9aa9938b2153e", x"f399612d176bbcd4", x"56278a5deafdfaf0", x"e197224f0bd5331c", x"822f67058bbe6bd7");
            when 12938910 => data <= (x"dda0934371935e7d", x"014b534b78ffd600", x"bfb9c523ec8d6f22", x"c48feea90bc7f493", x"41e65440c5deab57", x"871ce19c1f74302a", x"1d1e0acddc5eb65c", x"520f8268601ea896");
            when 25642197 => data <= (x"541b448614916c8b", x"5033c58e9b9f2a2c", x"5d9879394291e2c7", x"f14ac997274f2a0e", x"50dd753343a32319", x"a7be5a4f57bf56d0", x"2388d4b49533a973", x"aa1160a5756d06a8");
            when 25346952 => data <= (x"281aa3177ec32e9d", x"e975ba77fbd1901a", x"136477ffd5ab49d8", x"b8b9182e282e2fc0", x"159ae55a788d0ea4", x"fee67f9b548067e4", x"ad0d14baa9e73c82", x"ad965197b6798340");
            when 13502749 => data <= (x"f089bf03fb3c1711", x"f1e748cef0d2f0e4", x"976310518cc8022f", x"7a6b98d1a1bb5105", x"877b4cfbeb5f907b", x"1be306fe42550b79", x"45b5e14276d1865a", x"95ba0394c8d29aea");
            when 24638157 => data <= (x"40e855cda59d4612", x"3b69383c05aa56cd", x"c0066c57b9eeea10", x"cb3a95743aeec48c", x"9962fc2640760266", x"5c6c2814b20914f9", x"a26df1e806d7a160", x"fbd8ea105d33c217");
            when 26774692 => data <= (x"65c2190c929f5788", x"3e9ddee607f84d2d", x"7120c5c83969ed4a", x"081f7000fc888133", x"47d191f5e8d7897a", x"c1baf66a9f90827c", x"93add5d7fa63584b", x"37910c5fcfcd9576");
            when 12779088 => data <= (x"d396cf43b9d64fa8", x"cf72cb2091a66fbb", x"60b31589fad27fb2", x"3f94521a3ceed8c9", x"149958f711f51285", x"d6c3289a4daa9fc0", x"abcfe67eb0d4671d", x"675e87db18c988d0");
            when 1508124 => data <= (x"e05e903b52467542", x"238b00eccfe5979d", x"851b8d104a0f937e", x"7e522d51bd7e7514", x"5220315c32ee09b4", x"4e5711c099fa7ff6", x"59df71fbc6c2525f", x"76cf4ee7dbfcd595");
            when 29083191 => data <= (x"28d83e67a9fc0e1e", x"bbaf860d7422bda5", x"ea2402047844db59", x"c56f74bd1c29c2b2", x"5fc59e047d2183a1", x"cda37296b629d735", x"b07c058097086b49", x"042540e2fd778d71");
            when 29374490 => data <= (x"fb283f991145eb60", x"2f60a982f7536eb9", x"665aaa849c718208", x"a9f554a4dfdbd262", x"4f25a19264dc48df", x"a8b4501f34b93508", x"b0752b35101cd822", x"dd17b946e29b7d09");
            when 18211084 => data <= (x"dd7a4496490dca99", x"1c342d9d2baa2e46", x"c9ff304c4d07f680", x"c5d72c2fac2c9181", x"937c3cb59f2eb125", x"b0b6a969dab396a4", x"4559d9277e3ea357", x"9fb85b36bd0e9c0f");
            when 10644522 => data <= (x"9cc0c5a428de0983", x"75f09f9190487ddd", x"d226ecc96e3798d5", x"a3a0cefa0f0ed84c", x"d849b06056f5d664", x"7039a24d84c28bc7", x"bb4a0e1a3c668c66", x"c90deb97f6df6d43");
            when 24770566 => data <= (x"7ec21d8f29753c27", x"b6af24ca6b4693fd", x"1ce6f4ff70b0d640", x"055ad6dcbb64bd55", x"d6d0291d5f040179", x"935133a1e9c83b0d", x"61f32aaafed7c7f8", x"be62e2632aba26b3");
            when 23214847 => data <= (x"10cef0b2ce3c5a86", x"c4c25cddc6fd70a1", x"720580e6dd186bdc", x"17ed93ce330b6fe3", x"7ebabab25cd68ad4", x"e54e89ee181499e3", x"5aa458c389ae4efb", x"273b7554b3524a50");
            when 8557801 => data <= (x"7ac7b52f5e3aaa27", x"c8852b8246cced15", x"f0ec1d8c890d3b89", x"01a950f889e8a8a2", x"ed43975857d867c2", x"16f18cf8a9b93fcf", x"e1efbe9c3b45c1d3", x"b306687febbfe227");
            when 16833554 => data <= (x"3da07ef5a657c450", x"3ebac1f1a673ad2b", x"535461a8f89b4a32", x"92d62c36ba303135", x"13969b59166eed93", x"e5baa4a57d6439a9", x"7e7dbfac8713867e", x"1b746d5ad9767f6b");
            when 31226190 => data <= (x"56df2bae6f9cd3d0", x"32a778e210331bc4", x"9758c6ab1a05fe09", x"8a910f30c222d816", x"397df8a5fc30ffa4", x"07f4e537c45d8c0a", x"bfbb0584a0f5178a", x"3ae06715bc416c0a");
            when 6117467 => data <= (x"e2af9c370379da32", x"927441029dfab61a", x"9a705b465c0a7b99", x"1254eed2ee96f0bd", x"8633a3b46f99ea0f", x"5c3baab7e76ce404", x"e1837f88c9869706", x"ed34c19a36977f2a");
            when 22744838 => data <= (x"ade9c54359a22e1f", x"1476aadba2ad4cf8", x"3c981f4248741cac", x"58eb553d76b6d1c0", x"790d1cf2164a8ef8", x"348823bc8899554b", x"dc5b1b86df69d66a", x"a4d3668728693e1b");
            when 20127083 => data <= (x"22e6e6aac022958e", x"83b128abca55099a", x"611537759158fd3a", x"0c68ce3b7ccdba8c", x"e4b3bfff84d19303", x"728ee0ccc807d546", x"6915f94cd9db4f31", x"d5c48371c03e637f");
            when 27940218 => data <= (x"5cc87186522bb5a8", x"2c7e990e9a117f71", x"1433037322b89c5d", x"fa4ec9ee1968a9fa", x"08843dbe1d7f197a", x"5602df717d863348", x"dc67cd4df6714987", x"73d2be613f19d9d1");
            when 23368947 => data <= (x"44307bc5b226cbdc", x"7fd3c538d8bf4f3c", x"56c3105361d07e9a", x"215c9b40d96c6837", x"70000eecda15d277", x"7c14573f6eae9d9c", x"e728bed2ff85c4a4", x"e11d5e2321b3df3d");
            when 25191734 => data <= (x"e4c403f1b300b3bd", x"dc241a9e7d4c26f9", x"1d811e1d753250a4", x"25cbc7f07a451c97", x"01d17dd89d3f0ca7", x"b2645597131d9c10", x"bf3b9a756e1c8dc1", x"79b249ef57aa27e9");
            when 8469504 => data <= (x"4d7a6168ee9fcea5", x"d45438933b52b387", x"48b24bd96e142dae", x"00d8acd902a6fdc0", x"f2b150b102c3de2b", x"f56f02546312283e", x"4bcff63c14eeff20", x"11cfa950311a1df2");
            when 14700752 => data <= (x"2cbfe2f98d370ff8", x"bd8bb1508e09f777", x"515970324df989c4", x"1d22ae102e287cc8", x"cfcaf8ac7e082047", x"8ce2793db2ddfd70", x"01e16dd710b7abb6", x"de45a4a4add01508");
            when 14763498 => data <= (x"6c77235bc0cd423f", x"5c1658f248b02c40", x"1618a02d4a65377c", x"a19dec4689b36ce8", x"f17bcf3bddf26815", x"510490752e02b410", x"a9247d324e0f7e4a", x"26e910f534dc15f8");
            when 2254443 => data <= (x"82c16bab51748541", x"fcda9cba66df0c1b", x"f0bbcb38f29b5431", x"a786adb29e766c41", x"3178c48454bfa20f", x"3db398c5c805c1fa", x"d5801c11351057a2", x"da930c34024feaa9");
            when 28779538 => data <= (x"73b9fbe06459b53b", x"8e7851b8b0995095", x"11e3da273e5af897", x"468cb204a4f363dd", x"6d477260bb4f2110", x"7f56e1d89dfa6e59", x"afb09f0064a1a143", x"164449ba65bd5b82");
            when 24809532 => data <= (x"01015af0435e1c96", x"daccb0f0912e2b85", x"4893a9a4f351145c", x"f24f7fe89b0a1f6c", x"a61b0b61de89ce42", x"d380abcaee49f264", x"0b577185fd9180e7", x"463dc988dc0b32be");
            when 2587595 => data <= (x"5f89397a73b8cafd", x"1b7dfa04d180cb8f", x"76572ac40246d268", x"1bbad60f12bfaa39", x"1e47e2b1aea1c799", x"cc1f3f7b1d8dafad", x"34873fde0784d806", x"ed23d9c015d2600c");
            when 10818416 => data <= (x"14df38964c830379", x"ede8cd49e3f93868", x"fd4833766075e1d7", x"ede87774d4adae95", x"dc99788f92a97087", x"5468ee6742c0025d", x"367ccf4b1ce0d682", x"87810f1897217696");
            when 12150964 => data <= (x"a5c72d5b2094560b", x"dfc6fd14f68365e0", x"a90b342992eaa668", x"eb96b1c2db861b2a", x"fe0e3afa3aa9bdf8", x"e47d213cad33250a", x"4e1163a2a5b9cf79", x"d7e3967fec7a0159");
            when 29329674 => data <= (x"6076fd1f0efe0305", x"f5e650d945d6f84f", x"a5d506a7e0c38e50", x"cc4bb8f90f0cec9c", x"bf1fa70c84678a08", x"54705f01f9d2e7ae", x"c3316f4625d84740", x"0548c8a74d97a4f8");
            when 2791611 => data <= (x"5a8527223a454fe0", x"7c5261d0bae8c0ec", x"429a397b049f96eb", x"27797fd4bfad3124", x"c2260100e3d523d5", x"f619176da9f19762", x"7234afc252ba6924", x"9b2817df02de62a7");
            when 15606129 => data <= (x"e745be335a684045", x"e9d0ead9aeb866a6", x"24715b41f9c0d50e", x"d0d4cdfb90150ee9", x"dcf94b16ae1ddf14", x"02c48a937f63bdf7", x"286a4b52c04e4e91", x"6d48f060f068268b");
            when 23755388 => data <= (x"0fcb91ac842ed876", x"a6708134e04fc978", x"b0e71b371de33314", x"091dda404e43b5de", x"99153582b3c76449", x"a1af1dfb835f297a", x"ac9b0ec2c85017e1", x"a39e38ca49d4c975");
            when 25898380 => data <= (x"cc1f6a18e57565f5", x"8bc31b902ade79a8", x"880992852212c573", x"339091d9b1f66d50", x"a117bb09da0efef0", x"adfd10febd33068a", x"cd6b7149035f0e10", x"78dfafc2b70d8fe2");
            when 18298379 => data <= (x"61fb79b067b55e99", x"465d36c22e35c86e", x"2278c690e2049319", x"4872d4f3df569b1f", x"34cb932bd278732c", x"4ab9b21dac2e295c", x"9284a6d250594e9a", x"2433f7d7fd09e2f3");
            when 24561934 => data <= (x"1d0d0f2850abcbe3", x"3cb15d4cb7f67ff7", x"df3d0aefaa411c77", x"5dce82437723db80", x"75ebe23704bde34c", x"26184a4af9f7f746", x"0e352595c4ad07cf", x"e48968f63b8e8e0d");
            when 7999364 => data <= (x"039a0ecc780aa22b", x"da8d457d5b8d3927", x"2ba1b7f56ed096b6", x"cb47f826644f2359", x"9eb087a333925ab2", x"2e474fcc29a85182", x"99979b7c14fe8a02", x"b982d5d73cdcc0ba");
            when 6296496 => data <= (x"498f0d6f52ea1481", x"2442b5154d6ea273", x"2f330e6dd529a654", x"18553bbdf64d8915", x"d484d21408478e7a", x"fb397c665d360ace", x"d9225973a76d64c2", x"ef4bfbf721be415d");
            when 27317259 => data <= (x"2be8f8aa040f724a", x"e00bc4188bcdbc16", x"b753d889c6cf2fe8", x"e20afba5ff2a1c79", x"2a9421d02e7b3fac", x"9900bb96ad9b4b1a", x"7984150f95631cfb", x"95d74290df393283");
            when 2803830 => data <= (x"40f63dae1db46244", x"8e0454aecece77cf", x"2e635e85a577c0fb", x"da99f88bfa8a076f", x"cdd8db8232a9849f", x"b162e5db909b7734", x"1bb52db15ec12a68", x"d9c9ef65906dc3f0");
            when 30062060 => data <= (x"f977981f8ba6b21a", x"94bdc839f05904cc", x"bea7cf8836ed4663", x"e0b16441690acd89", x"c96c5f22d4733489", x"66943999dea5fab5", x"2862024d656a4bbf", x"e9575624d57c8da1");
            when 13735555 => data <= (x"bb1e34a77c8194c4", x"412e34ca1a931ff5", x"643561a8658ce8e6", x"a4df79286756746e", x"29fe9d3ba9d098ba", x"c673e09fc888b268", x"c77a7cf4ee1fc49d", x"b23ffb1d63e2a696");
            when 25628356 => data <= (x"fab51aa3a1e7e8f2", x"6b3590e0709f0fc4", x"c5d3ed6685e3a030", x"b3589a6bfdcdb3c4", x"48c1c2e04834c76c", x"821872de286b2fce", x"40cab1efb13488d3", x"12eebe545ef5883c");
            when 21533778 => data <= (x"8ca94135921b7532", x"80c7fdeffff458fb", x"c16694cec5a51dda", x"8bae6a5977f4c9f9", x"19dcb381ac0be419", x"349a21b8e68cdcbf", x"fcc96d20ebdeb380", x"795b2366461283cc");
            when 30065732 => data <= (x"1b793d0ede1b0e6a", x"ae6552b55d75fa4d", x"4e98430a6db00682", x"0a849ecd1a9537a6", x"1a5902c548efdfc4", x"a344ff4c2b52b06b", x"d1ac649b12ded87f", x"e64db53445150936");
            when 25767911 => data <= (x"67ccc09d653c3e6b", x"e9f58f2f1cb6beb1", x"7109cdd941874211", x"ea18574eb4fdeff1", x"282b0909577676ba", x"ec1947f9e178d43a", x"be6e8db5273abddf", x"7c2acc3612c6b7a9");
            when 32654977 => data <= (x"b5f8e6603ec20799", x"e717ac865eaa868c", x"a35ac8551826ff83", x"9e020b9c3b34e5df", x"e19d73355dabf158", x"35fd30c93281fb31", x"80007f8b485921f4", x"0d9956fb4f668f88");
            when 32871099 => data <= (x"283b8a8ca87fdfc5", x"a03e8bb447b2dba6", x"a63edfeec0fed675", x"8c101733184fcd29", x"a32b9c1810512328", x"93e606e5ec72303e", x"1a31ca82ad9afee8", x"47f76bac6beecf75");
            when 17624298 => data <= (x"b3a9e9aa04c57226", x"27cdd343f193bbaf", x"46d1c67714ae9d06", x"5af083a1110eea66", x"d695a344826e1c5c", x"c8b6e6e52f739616", x"44bf1c9f546c1c90", x"fbebc9776acdb6a9");
            when 31343581 => data <= (x"bd783d0cc9772117", x"10eaaf64883c319f", x"2c5aa68d5308beff", x"141a243705f1ba22", x"0de0a880ed976962", x"12d345c427451347", x"a7303a520c9d22b3", x"58aefc537ee2f4e7");
            when 31094760 => data <= (x"86855bc242a14245", x"dfce50e0ccf09d8c", x"1e7b9ba7dcecd128", x"1e44c4094584592e", x"3097ecdfc5056b19", x"3034827124faa45f", x"08837f2e3671497a", x"d8bc7aa03b93b707");
            when 15599841 => data <= (x"a987890d29377fb0", x"48a30ba899d148a8", x"3f7c566265c41374", x"c167bc09383f164e", x"2d995bd7ce4db7ff", x"2c6f05ca83ffdb68", x"3c87d2d4f17bc591", x"b30379eb5fda2254");
            when 27148338 => data <= (x"c4aec27d82ef2e21", x"5a2d14371a89359f", x"5169f6d2de778ca7", x"15bfa26b6c71554e", x"9a0c419174c7fced", x"f3dc7eccff9a60c7", x"bce1a32df8799547", x"0642e41fb52a7961");
            when 544753 => data <= (x"e7abbefb0d51fdf7", x"7c61e4238546cf5a", x"f3799155febed3eb", x"5b9270a8c8bfe034", x"2850a3f4540655e6", x"1be223c5988c7a4d", x"b2455565a5e3eb14", x"4c4469ff0aef051a");
            when 16338610 => data <= (x"2557e6fdc1eb7091", x"e3334c9d038262ad", x"2746ffbc6288d780", x"e5726e79699dabf1", x"5993e81324168467", x"1513bed56810ece4", x"2319049a2851dfc9", x"83706a3cfe7ab272");
            when 28454356 => data <= (x"71f16c9d7825054b", x"e5101d2052450ef3", x"b23df2e362c30a81", x"3d4897e884be088c", x"eb246059e4e0d941", x"e84d8924fa697a96", x"7364a8e4e5f65d6d", x"56ef52ee85a760a3");
            when 30944651 => data <= (x"619cf109a1ca5b7e", x"fe3e02d2cc50fd89", x"6fef9155cb8378a6", x"8354ac31e9fb7aa1", x"92c450d0842087da", x"98c12cea08b86895", x"ae40c627efd48fec", x"2cf9ac3923a1803c");
            when 27427309 => data <= (x"461c86caca7f8ce0", x"4dd9529a2904acf4", x"d6466f1433d88cab", x"2014cb8dd4beede9", x"181e0d102d84d75e", x"7e681985f0fcecde", x"3542ff117ec6b6f7", x"841e9f983dda1bfd");
            when 27143630 => data <= (x"71b49804dbd22d5c", x"46bd6a56f6604926", x"9cfde6ffa5eaa841", x"ba7fc35804cb661d", x"9226454fad2c0689", x"a5aff74e7bd153c5", x"e78d80ef9ade0193", x"17933e927fb3ffa7");
            when 11870931 => data <= (x"abbc4fc45629d3ad", x"f6d46e5510fe764a", x"16b554237ca67e70", x"62527f72d66ceeae", x"88bec20a23dbf831", x"ad7bfcdce90e2173", x"c110eae133edd585", x"a5221acab67e83d0");
            when 20526387 => data <= (x"d1452943f0c23386", x"d5592ae3ea15697f", x"3e4837c6cdc6180a", x"8a1a28c66eab0d6c", x"6c30d9cbbc995e05", x"d3ed706882056068", x"31cee89c841d7a29", x"1902d33c641499c2");
            when 14007541 => data <= (x"a0e4e3e837d93156", x"d67feacb4be86659", x"516d003e452c700e", x"fed18b05359797d4", x"b38a3dc6ece87a95", x"af4540c7dfa0791d", x"8acbbe8896770484", x"5baca2a42441c97e");
            when 29217919 => data <= (x"14693cd6324d284a", x"e1264b19eb3ba584", x"96dd82e33f967f64", x"f62f58f3aa93fbee", x"17b0e7173dcd94fa", x"608bb7ad95f142aa", x"c49cbbf6068fa102", x"3f84858ab7ed6919");
            when 16358847 => data <= (x"d3169adb1606f3fb", x"5f7b41e256190a51", x"ce54fc1fd1b62bb5", x"18e17587f4360919", x"05436a72ca5d6a89", x"0415ec7cc6b0b347", x"947868b2df18a5b0", x"75b9a3e037d8d923");
            when 12233952 => data <= (x"c056bdebc63b88fc", x"209768941b60dbf0", x"e734e709448d8530", x"f2e1d718d055783c", x"eec489aacf32ede2", x"deebb48ea3533b12", x"5951e09c57c1e47b", x"0c8baba0a1baca26");
            when 13597657 => data <= (x"c4ab49230e3c7db6", x"4659acdd27c3ae8a", x"b12eaa40505397ba", x"6759c41ade5cb78b", x"37543a57aba7dda2", x"a496e41d899aecff", x"12c4aff554e57beb", x"79ccfb01a4dea2ba");
            when 22637426 => data <= (x"de8df48066ada41f", x"4dc2dd9726635aa9", x"4add211e1369c167", x"81bcc210ad8913d9", x"2b4e2b8eca8f4bfe", x"cfa406e59eb81270", x"bbf58fcce001cc0e", x"84a260ab6e45a780");
            when 29676087 => data <= (x"5e84921006f08d45", x"f9bed6ae260291cd", x"940467b7709298e1", x"7c15f587a1162120", x"23349913a44a0949", x"b9dc1066d803728d", x"fd67d96d22bf2093", x"835f847ea4e12f14");
            when 14374829 => data <= (x"fe6547fc04f65c88", x"4ac7fdb6eed8f4c6", x"9da10004cfe4bed7", x"13ad50e340508e56", x"867a8958062e02bc", x"edccb6df6c7250a1", x"a04b7cb3329026bc", x"5b7d4002a529ead6");
            when 29789539 => data <= (x"3514c61a7d124898", x"a1798e89552379a0", x"51e925afc5e94216", x"fb469922c4125e36", x"c0f56fe395663ff3", x"8ddad26b7d4de8d1", x"38cd3570532dac56", x"5d2af6156fa25c72");
            when 30425002 => data <= (x"e7872b312b06b9e3", x"2229a898897fed69", x"f354a7132ef7f4ff", x"25d4f4adf030f999", x"a7e9e9224e826846", x"ef5c3d41bfa823fb", x"91d07c553f2239d8", x"9e3401ac82764383");
            when 6822293 => data <= (x"be9ed10d633ddc08", x"9bbcccac8932cd1c", x"4886fd828a25efe4", x"cd05a0109e8c88fd", x"b38dd8dab704720e", x"00754304c06a6f91", x"59997a8a9891c7c5", x"414660fc5a8340d5");
            when 26441788 => data <= (x"648678086306decc", x"e1d1da442a71562b", x"f04bc7f6605ef4b1", x"1553ce11a30015ee", x"db1a126f9997d363", x"9d274e470f42460f", x"64c093e8fa594b45", x"b3913d415b72afae");
            when 11338978 => data <= (x"2c9235398087f33e", x"1d4d0b4aa6bc260d", x"bc778fa6892f3885", x"7b997ced8d3796ca", x"ac139c88c83dbd2f", x"de1abe21361003ff", x"1c86981dfa242053", x"e2a92e337d359411");
            when 7607719 => data <= (x"a4fd56756f40d4ad", x"ec9fc740e785664a", x"5bc3bb13d0d999d7", x"87f54bb59189d72b", x"a2fa0af6b2fbba98", x"97b402810bbbfe26", x"9a47d74dd54ff4a9", x"f3c921bde6329b7d");
            when 31553856 => data <= (x"67f626207118c299", x"eeaee4eebee71ce7", x"963776a20f0a58e2", x"afdbe2028fcd90e1", x"d838a45680e4bf0a", x"b320379ee3184f7c", x"a19e8cda79a95c3b", x"6b69fe41c95e89f6");
            when 8789447 => data <= (x"19cb401150ef26cd", x"2e776955800291a0", x"5e4336512ad716ac", x"30983fbec99f6973", x"52ea4821d0d2addb", x"7f5648a7be13f144", x"e6f4f495fd140e64", x"021c462b3a55bde1");
            when 30613305 => data <= (x"9db367d399ec8784", x"679e6ce7165b4077", x"0898e94c4302b886", x"5dca82803b5d7ca1", x"2cac4e2aead7307e", x"4fcdb9b95a770581", x"39de26722f627493", x"ec4701c6046c2fbb");
            when 18146842 => data <= (x"83c4b13355591d81", x"e7aade48396184a3", x"fa22f877e01cd67a", x"9215b4633b4aa37f", x"00fabebaf5c47111", x"87f448bf239ede40", x"ee24f3bedf8e7d6f", x"70df8914830f549b");
            when 14516496 => data <= (x"d4d45f41c5c5edf2", x"a9842edbcea22777", x"789b3d0b3ffae261", x"ff13226adf3d8ef8", x"fa9057365c4d982a", x"cedb6b13719a0c7b", x"9251a1765ac14a3c", x"488c1d13e08a2536");
            when 32590687 => data <= (x"ed3f4450aa427042", x"5998bbcfe0ceddee", x"ab2174682bfbcf60", x"ccfdeef7d9e8fd99", x"578de0751021ea1a", x"5ee99ab3da206f30", x"45c918bed1df2e23", x"0973cdcfd48aa0aa");
            when 14830946 => data <= (x"c77c0b7f07b4fbeb", x"d15826c9beff917e", x"e8f212bd2927958f", x"cb1f999880c5c58b", x"52d38421cc09af9f", x"aba9eb8f18677f87", x"9f89af1986a4fd4f", x"2867c477b2d3c547");
            when 17627935 => data <= (x"7f2c718e8fa06ed9", x"096cef055ad5bad9", x"32ddf3166668a734", x"10e051a58f795fd7", x"ceb39bb9d9fa3cef", x"fc5ba2b981a98572", x"52ebb36272e4d4ee", x"2c03a6fa07c15294");
            when 10396249 => data <= (x"4d8d0dd09e2daffd", x"1d2012976675e4aa", x"5861c400932e61b3", x"792c2801e1d0a0c4", x"d90d425ea678403d", x"211fe92f734addaf", x"b175c201e895fec0", x"d97541c60742d29d");
            when 9197541 => data <= (x"f3405c98196c3995", x"2e4d9ccc3106f514", x"c1ff573b99097a43", x"8dc2476cfe5411e7", x"ba7d18ec0886288c", x"2ecd5fd94481e5af", x"692d2f8fc75ab528", x"77d1b1f635ef6506");
            when 20160866 => data <= (x"f7409143538b8ba8", x"4f638127972c2495", x"0df10326c051e27c", x"2d5ff0b0015a5894", x"1161fccf8db5e06a", x"974f1c1c2675a9b1", x"22fd4b47fbdb464d", x"04f3bd6c3c725046");
            when 23594010 => data <= (x"e5a2f96d881a5ddd", x"b3313538a59969ad", x"8fe7ee61efd5cb6c", x"f5a0b2a6043e5301", x"6fec0a7b27209383", x"f7e49ae2381925bd", x"a574acf76cad8122", x"6c215e39736abdb8");
            when 31031857 => data <= (x"7a7361bbce4d95d3", x"dd9eb2dd1fe6e277", x"51fad5cf5720ee8d", x"adcd4078e039a480", x"7949e50b8650a509", x"46db7c3d58775b80", x"40a29bb6b1484f98", x"7b04f140486ab8a3");
            when 13448570 => data <= (x"7edc422e15e37647", x"b04eeea4d4cc1a81", x"b5c2b3f4d44e9db9", x"b6860c53a5bd79c2", x"dacea60bd66a438b", x"5e8e69274e0b743a", x"559e309832a2f8c0", x"3845c783e9ba756a");
            when 23402545 => data <= (x"745016594c693253", x"d690a5d9e422e84e", x"ce8f43354a271894", x"b59cf23ef8ba86b0", x"ee499ad1947b1221", x"bfa3f17d4e0280ca", x"636207bee50f8ab5", x"c9fe9e3d8517853b");
            when 24082009 => data <= (x"d77df1158ace0382", x"76c532545e095a39", x"8f2e437ad4a49f0e", x"8f9103c4c0d4eccd", x"713af5fdae73974e", x"809cac007b180eb5", x"e21421bae4c7e79c", x"af03df0c6adcfb33");
            when 28646054 => data <= (x"1be044b13110950a", x"597e58572fd416a9", x"538d34d77bcd1158", x"3eea89b1aecd3e79", x"45621bb73014243f", x"ec41500f8e456658", x"fb9994a3e07f41e9", x"e112b4a6e972b1a1");
            when 12285141 => data <= (x"5c63e83b14404186", x"cd5722623dab0c24", x"5ce8f5e36688dd57", x"317ab60711f18ede", x"2162e2a7833cc919", x"bd94cc1b9da2a593", x"986e24a1b01e380e", x"7b493bd307228926");
            when 26589467 => data <= (x"c97891d23c2608e4", x"c8633d502136360b", x"deafa57e0ed9496c", x"84cbac19a1d3be89", x"3c8227680e4315d5", x"bb239fb08919ee41", x"4bc960485187f951", x"1f3d03716ccb0c88");
            when 4677566 => data <= (x"362a342f28641c84", x"98f4fe0374d1d654", x"398db2be6abaa96b", x"99dd43040c52487d", x"b07b1dae15c2d3c4", x"681c101bfad411ed", x"1a0876f571730488", x"f1b8fa3b5d16d06b");
            when 5177986 => data <= (x"d0228b9638f24dba", x"9b66587f305851ee", x"19b7d1ea5a1d4172", x"bc8597ea93903836", x"cfb81c471fcc15ae", x"e6df8ac6b7622c43", x"6533a5f2fc4b6837", x"b15308ac8d489e4e");
            when 33465500 => data <= (x"48b6e4a6d5340763", x"e6c93d2e20195f07", x"507f221226ab6a21", x"4b5a1966bb67b05a", x"d735d17cdcb7c8a9", x"73fc0219ea6c6de6", x"180317be1f9b7eba", x"1a467eac76396203");
            when 9064967 => data <= (x"65be5b348993b4d1", x"f120dfc1e23a2a97", x"402aa8d8f1851de6", x"ebf62b20a74592e3", x"3d298152df07ddfb", x"472fcd330cec7b6f", x"4ea545866ee067f9", x"b34ea0a7dc3d8118");
            when 3567412 => data <= (x"f3b403a378971c8e", x"1174411cbec36fdb", x"7aee107ce005039f", x"3c9d94e6a2f570cb", x"f6e2ba4e1960b2ae", x"2cf2d0085c14d4b6", x"09c80d4c36436e66", x"c30d76b3cbd17dcf");
            when 22712764 => data <= (x"325f56fa2e430907", x"c698b75a86dca301", x"9a883c14bd50840a", x"ef80cca6eed9d69d", x"abae659d81b76dab", x"f69cb21e9dfe06a1", x"115201de11842c15", x"9d91814da88a0ee8");
            when 8880864 => data <= (x"98e57ffe93b84537", x"226242fc6d9f22f8", x"4e1e392632b0e6f1", x"4fec1870bcf18ec8", x"d98946eef6b047d7", x"aed510fdd609a0e4", x"2bb5b8294c44da33", x"4bbe5fe4bae2021d");
            when 3606953 => data <= (x"5889e3db5d462570", x"c77c5f4189b61e51", x"7be5f79c47562d82", x"f63c08c1105f022a", x"4e9a206afa33956e", x"9ea0f48f1cd11a04", x"2f3769e6f7cc848e", x"c8a5549a00272160");
            when 2748160 => data <= (x"3e79e86f58421229", x"8fd50c8888fcc623", x"8c7520423d059925", x"3a2ee050599c89b2", x"ba796ea5c593a16f", x"c6e60fe096e0296e", x"8342bd4690343297", x"b211ed596ed0ba26");
            when 13179343 => data <= (x"acc5a11439e3eb28", x"63a025f3ce1c1a1a", x"fa2393dbfa1e9d77", x"294134288cd9f70e", x"82fb5855b46ddc25", x"596f4c8a326544dc", x"fcd41530aa3d2559", x"1dae6690ad9c3ae0");
            when 1826162 => data <= (x"aca6df49505c8e1c", x"33587f9bf69fb4e1", x"5ee1ed0c6e047554", x"1b2cb2e5037ec325", x"678aab712d962f3b", x"cebb8efb0c4f2744", x"272bfab7244211b8", x"628b9789920809d7");
            when 7222704 => data <= (x"c13a38827ac80207", x"59c3ebd9c21f47ee", x"fb85436cd7a06c58", x"a94cebe5ae9aa3b8", x"053077403b1bf2e9", x"5450bcea5af92db8", x"c236a7fd867d2074", x"92c7757437f1cf3c");
            when 15427756 => data <= (x"df636820b34e2e5b", x"f753ce9fee379564", x"5de15d4412f7ff22", x"e1d5e332d44d9d4f", x"8c3c95b136185820", x"45fac48a3907da25", x"b008e53db761ba8a", x"625d04bfb4507690");
            when 25369528 => data <= (x"55d56fbb1dbe35fb", x"e30f64ee234a473b", x"11edd6dc4afa60b3", x"7a27e9c43761d130", x"4de246c0cf6aa465", x"77f6816a42786710", x"d377e75f13b84ef2", x"59be925c443b2783");
            when 32921526 => data <= (x"7e0fd94347170c75", x"92cc414a5ede2beb", x"d521f2617b73010e", x"9e72ecdf9f0b1e42", x"498fcf6bbe0fc674", x"c17ce293a2fe6e44", x"8f029a2b446db682", x"b34ed4abad3a9e86");
            when 5297139 => data <= (x"1f9cf22340478c3e", x"9849f34abce4ae1b", x"93b8d3efba760d8e", x"861b3082eb89939c", x"df4c16bb2226bbb2", x"3224bb3375e368ec", x"3941d738e0f732d8", x"544b7563550b0935");
            when 22835209 => data <= (x"92aeae2f3842f0dd", x"0e62bd2e3ebfa19d", x"c8e23f57483f7bac", x"624b8ac478553ed1", x"ac7d72bf53382538", x"c603cd0e20daf860", x"9d219e4c41ea3540", x"5f1447bc6f1ef252");
            when 1886254 => data <= (x"054e2cd2ef782090", x"f62e4b1076970f8e", x"3c6fecef99ca304a", x"dc840f36dba740bf", x"4064ad12d798afc8", x"d0d3cb872cb8c709", x"3704df25a76daa16", x"01325ec99bb36912");
            when 18410759 => data <= (x"a6a9625a2874071c", x"c2ffc2ab65030db7", x"b67f8ba738d75f0f", x"ac1f926f03681723", x"0a1600282ccd21d0", x"f74f7f17a8dd9b48", x"7e5c21247e196ae3", x"b26f78ed8b82ecd8");
            when 11765092 => data <= (x"3d9c40d203fad610", x"29d52dd4d8a1c6e1", x"d566538fc6bbaff0", x"3557b2233d65b411", x"22446f56f64ed933", x"6aba1692e2cc88d7", x"c371c10d2314292e", x"c2e124a17e69729a");
            when 32118048 => data <= (x"f8cdce92bde2f261", x"1fe6299c7a75267a", x"1b2be0e21deb6a28", x"b5c06594ee001c36", x"42b0bd79f7007444", x"5e4c9d42ea5999b6", x"12a22e3250b462ee", x"732d154a54e1126f");
            when 15169737 => data <= (x"4793f28cb4d6c3d0", x"a07a5125a2e16873", x"9bbcfd9eebe155bb", x"e483ede1166dba5d", x"e0fb8a5d1edff15a", x"0ea4672e883da84f", x"3df024f78ab8121d", x"0fe155f9f21fc316");
            when 16417224 => data <= (x"29a90a39d5a4088d", x"44e3f4818b760786", x"97ad6259881c1d9e", x"49fa1f6ac8e125cc", x"4210973f7db7a60c", x"2f869260be72d84f", x"a4af19bb121afb66", x"2bead1100045dd46");
            when 29542177 => data <= (x"b84073c67369bb09", x"38cd631deffd0bcc", x"cea0e46cc41c7e26", x"f015c99ca0e6c834", x"1f300d7e25e36d28", x"588daf12b6c0c79f", x"ce27ea882578dab2", x"74f8754d9c622eae");
            when 2876707 => data <= (x"2a9e0c45c2cbe99e", x"e35e4780a62f294a", x"32ba1f1577b78f4b", x"7476ec5d6ccaffe1", x"fabac1f1ad25803c", x"a74044e1f255e1c7", x"a603579cfabd55c4", x"559dc6afa74262d5");
            when 27859526 => data <= (x"ee1634c3bdcbcf72", x"f39a71db788ab0a3", x"d5adfc1e9b11e4ea", x"52ab849aad3b2872", x"72a443b2d04244b9", x"f3b26d3a6fb26208", x"dd42582b2b2ac4a0", x"99fb1d8c4d969ae3");
            when 12774959 => data <= (x"4962f9cfef9f19b1", x"82361b491c7f249c", x"615e11e3c17b028b", x"85079e976ebfc86a", x"9de8cc57cf6ebbb8", x"63ce7b51044a42d7", x"0fceb27bd1ebfe21", x"a701f8753cc620b9");
            when 29325852 => data <= (x"bc3e7387914f1a9c", x"4114993e56f530b0", x"eedba07b4ff3dd15", x"27b5eb90d8102429", x"944934ac57f1409c", x"cbfef3ca67dbaa1c", x"b1544c8177f8a4b0", x"a3e67a0b224a55b1");
            when 13906967 => data <= (x"adb5973b514f6174", x"d9cfc7a522e5bc9f", x"b927e5202926fff3", x"278333824b95ff3f", x"f1e3b7a4fe962348", x"06945ba0d6d94a2d", x"2f29b7ccf2974a5a", x"bc875434ca228e65");
            when 31312428 => data <= (x"6ab1fbd72b3116c4", x"f2074b865dad9645", x"56b9d9e2ec1bc03b", x"4688d1deaf35e65f", x"1431a5f726757bee", x"31e8060e2ba71f09", x"f204603729a700f4", x"febd7705d890ea1d");
            when 9130997 => data <= (x"797255b42429cde4", x"5d391a18d2138f95", x"b529394a72f74697", x"e3389c89aaa8f8b1", x"08a4b9232af81380", x"a1dff75a8c446fc2", x"2a0bfc7e792825c4", x"29e10e334a816145");
            when 17953129 => data <= (x"d1d490611b0fb698", x"6153814d2ef84b3a", x"dc427ee1078591c5", x"5a2e6d457fdd9e5a", x"19eb378e232c7547", x"dc477c4a4160b96e", x"8b8babef4e8c13ac", x"d567a3b23301dd41");
            when 18829961 => data <= (x"55e4c88d0ad6d7e8", x"fb282395a24501dc", x"c8a1ef82e84cac98", x"92b43867ae3899d9", x"9a41fb22699fcc95", x"b9c3ee061e41336b", x"9d0ec1429dbcfa49", x"4d74d1d78a4e2518");
            when 30525663 => data <= (x"dba85246b2fc2c48", x"cfa5d27fb1ed4b25", x"091fb648e83b940c", x"65d5bbbe62c77e28", x"0dd34be37d6820ba", x"ec68a10202540055", x"54d46cc1c79badd3", x"348226e7433f6b5d");
            when 1539767 => data <= (x"2dce7aaf025fa9af", x"8ec55de4b1061a88", x"f17f03926acf610c", x"8fdd81b321a8a465", x"4f5bf0e7f190e0e3", x"1d8167f0e7fde59f", x"3f779850b82f38fe", x"578cf35e335dd6c1");
            when 21140356 => data <= (x"81bd15c5ad88ae45", x"be03bc39e3285588", x"21ba110d7de8717e", x"584322b603dc70cc", x"c38ac8b4e8a85583", x"2e8faab947239593", x"2138ed287e35de65", x"7405832f2929a134");
            when 2321357 => data <= (x"c215d35ae502850b", x"2d7a79af00343249", x"8d7e8f15c3a107d4", x"a07419c52f293667", x"de97c05c66b7636b", x"f06576ba76316836", x"183e14a0b6f3f8ec", x"d4aed9e7298dcf1b");
            when 26959221 => data <= (x"98ceddb76930360f", x"1310f789cfbe83b5", x"efe6fa32ce6001b0", x"add48364260c9ea2", x"cfc9ca465c71503b", x"77ab36cdfcc95563", x"a4ff2a8281e8c25d", x"3913d209e49bfa28");
            when 14684255 => data <= (x"c0a110b5c06b20c3", x"cfcf70c9d8abb887", x"bb9baba21fe1aceb", x"ffcbb61dc721e78a", x"57932d4e0177572b", x"55280d188cb2222b", x"2057684cac99280d", x"0ce56ee63cb7d986");
            when 30405645 => data <= (x"d943246e4a15616f", x"be5493661209bc7b", x"1d287e2c30dfe1a1", x"5531f91940b340e3", x"2b2eaf20c52d9457", x"f12a26abf24237e5", x"eca21ecf3ee7646e", x"c60e766c226ddc18");
            when 31545103 => data <= (x"69f620cb9c1b5c92", x"c12633daa7a63abe", x"7209c135f88c7137", x"32f4f40b6d70be18", x"256dfa59a71de6f7", x"c84c89c4b7a936c0", x"61921648b1bbd8c8", x"8fb3fdaf6a6c048f");
            when 6973651 => data <= (x"1fb2d05b84e4b757", x"a6fbc110bef04ec7", x"a2b94efe61745943", x"5f26357589de344d", x"1735c978ff83fcaa", x"343299cbd1164377", x"2c50d48d1bbd5890", x"1c7ea94b52ffa2e4");
            when 5917639 => data <= (x"3859db97f6f3f481", x"cd0c7b53c28a5cf8", x"7481a2b335818d07", x"02c222b26dbd1246", x"cbcfb5468b1fe1d6", x"008095c56dfe393b", x"b0d73cf4f24d692a", x"f49d00fb8df0f93b");
            when 3361303 => data <= (x"e873764a3f15242e", x"3fd4d1f45d05811f", x"0980e3eb5d2dbe5c", x"53c0fac692487d8d", x"3ae717f8429dbf72", x"a421092ea5a33ee1", x"cd26ad08551df228", x"caf10ef8c642bde8");
            when 29369994 => data <= (x"dc34cdb6ea0cb87b", x"91960708ed870420", x"4a30b84304e4ab89", x"255ba5a97c1abe4e", x"abe3a15d24a1b822", x"ad160132cc676461", x"bba80c013fafc772", x"a1b5c15050863b6f");
            when 12802063 => data <= (x"78ee791964f2de0f", x"7e0fa6a19d01bfd2", x"5a28f16ec73d24ee", x"fdc47b1af0975f04", x"2ad974e14525d045", x"a699ded5999723ad", x"b9bf9d1218849ca7", x"2893df3cd8cbaacc");
            when 33250548 => data <= (x"650be030bbe22f48", x"3969971af9d7bd12", x"92c09e3b582d48fb", x"bf48930581a0b669", x"11a3cf87f20619c0", x"a1a0ab48763392f9", x"ac8b44143934fc3d", x"b80a810599d00923");
            when 10563501 => data <= (x"10cce8353b788460", x"5a0a3b443f747fbe", x"020009a5aae6d69d", x"6dd997d39b8556b5", x"b97f55b55c13016e", x"579e5b79cccd6dc8", x"092e1ec7178fde87", x"3dac6f92def7ea30");
            when 22945404 => data <= (x"58e0374ffa62e3cc", x"5bbb6a678a007d1a", x"910b546f22fde18a", x"58c2d10424d2d9b0", x"7047f6a3aa7eefba", x"9a54bdb2835a58da", x"b34060c9d2cc2ddd", x"8f5571cc8ca96ea3");
            when 6029446 => data <= (x"30d4ba7cc7bfd89b", x"22f3b2f455f13809", x"8d07ff5ebf412bd1", x"66fef771f55910ff", x"7086b6795a3c8440", x"689af8e212baab32", x"8142927efd6bf426", x"8a298475d0be585b");
            when 18150908 => data <= (x"e2123a4211060bb8", x"a7c1d85880d2df84", x"f76728804aa366ea", x"fc084f2f99799ec4", x"c9968cca84c557d7", x"f31d39b3e665b82e", x"fd6e80a4d53521a5", x"6c6933ad16a2e9e5");
            when 26386040 => data <= (x"132cdf8f26071bbd", x"91e1271eb1184f4f", x"17f91dea676ce6f9", x"bc339b117b0956d4", x"2890f8ecef1a681e", x"dc0910f5e6a18013", x"864c939278ef3e17", x"d483d330a19f450a");
            when 7610918 => data <= (x"efcad9629d47de19", x"9f178bfae358c727", x"4e3440965c09f2d1", x"18be2de35471315e", x"95ca1921ec5bc696", x"2b2f03a52e8a43f8", x"2671ff0f81287d59", x"adce6b1c60d39421");
            when 33606268 => data <= (x"60fa3b83a31b7e74", x"e3cf5cced1b3e3f1", x"e9a7c6c6cb62ef68", x"311ba57888eb2e5d", x"d4381698c891c47e", x"e4e9306e7793d0f4", x"94f37f2bc1a59ef3", x"665dde6492fcb22b");
            when 32188052 => data <= (x"e1e5e59c6f40673a", x"ad401ed49b9993bc", x"fc11f379edd8c96b", x"fa5efb2baec81ac4", x"df0f6f112b62acdc", x"56230200313d08a2", x"7d497fcb1abc9753", x"9a8606999809f951");
            when 22630742 => data <= (x"d7d496e3b1306d90", x"08bbc7d2c80375c6", x"8b5b5196c3f999b7", x"80a458f6071e1abc", x"100c4b64e4f589e7", x"b60b1bde8b7c935f", x"35a5c24ee7aa9f5d", x"1172870b8d9b19f7");
            when 30592465 => data <= (x"13cca6983523d33c", x"c78de3a84127ed5d", x"16146e29afeac8ac", x"c66d13f08ad4358b", x"b8aa86b5a030fa64", x"a5f42016f293b905", x"a02f6dad9a9b4556", x"4d08949e3b0fc8ba");
            when 13074836 => data <= (x"3810b17e1713d358", x"0645c756304640e4", x"da2a2c6afd88a36b", x"2c0291310a463aeb", x"dca2c699aab69693", x"a029fbc1c1e97db4", x"19d95b19d42528d7", x"32a75836af5e6d50");
            when 9042166 => data <= (x"db43e2322f093090", x"f8cfe91342092d53", x"997958e94525b933", x"b7a8a957c049dc79", x"9516f1dc4eda575c", x"0cc4b406e74e5842", x"fcd1a579c9368f07", x"66a1dffb361b5888");
            when 23549505 => data <= (x"71057f5606995103", x"01eec754dc255845", x"fb5c62052bcfe821", x"60be5651e5430b71", x"8e13f7d32af3d4da", x"b7005e71e1302635", x"4779cb7f9ea23844", x"e1d8164fc5e36c87");
            when 17620439 => data <= (x"755da7b2985ba86a", x"0b202da970f7b8aa", x"a810d82195d085ae", x"1f731db4969c2551", x"9a3fa55526bcebb5", x"92cfd5ce9591e1df", x"cb7f6999ca748df1", x"218937c53e55c0d9");
            when 31760818 => data <= (x"7b5a5c35f263939b", x"19e240cf2be29866", x"2218654dde82d39e", x"4b60e073934569cf", x"c5981076d80a6eab", x"129b0b3c17c145c1", x"6ed03b4d10a87223", x"18f803aaf55c39b3");
            when 29590757 => data <= (x"e40bbb903fceb80d", x"88689fa12db09a1f", x"16aec59fe55479ee", x"484f93c32c73f243", x"73950e72443b8609", x"33c97f810c02e47a", x"8ddd5211bb8ef355", x"b30659397c805340");
            when 19924139 => data <= (x"b400a48f6dbe458c", x"28c578c6916091c4", x"8cb44b64054716e4", x"2614374c2142f710", x"3627342e75f5eecd", x"cf51500d26226b41", x"0aca2a5c6a56b186", x"da377e256b65554a");
            when 15639967 => data <= (x"a5c555581d3fbe7d", x"dabd3cd5b923002e", x"9adedf13e8564985", x"b9b1366113af0fb0", x"0c8749149f9124f9", x"5e1019d4211d6512", x"72eb8e94beac3d86", x"1dc82685c95bad71");
            when 10386961 => data <= (x"ad0d177b3fbda64c", x"f596da3b72120fbc", x"d4d09b74798c3402", x"ba95dfd077802d35", x"69ed592c7b656200", x"b53f6da2a76f6c53", x"ac4392e84bbd2238", x"1c382bc0df616da3");
            when 18413925 => data <= (x"5a261038dc850b27", x"000f4642d73d94e1", x"7e7497f869518c86", x"ec95a0bb93db21be", x"01426abbb0f7e221", x"8b323f9d3bb22da3", x"77afb3b4e6e383f2", x"ab646891abace325");
            when 18653240 => data <= (x"44122334516a05c5", x"0659c4240526264d", x"45813afe413b796e", x"78a75121d62197a5", x"757ed9cd1070fda9", x"be317007066362a9", x"5190e04c61261c72", x"8cbd39ce603b59b4");
            when 23705541 => data <= (x"80db42940f11e574", x"552be0c2a5c11bc1", x"4f14fe4909d20b7c", x"6fcb279dfb5d165f", x"0c92a0da962ef6ae", x"456dcfd36e326bba", x"e7e5e4bc8bb4591a", x"02bc5d9373380ce5");
            when 17771997 => data <= (x"7af4eb78c20e4955", x"17a186cde614f0a5", x"4baf0629e60c802b", x"f9f74d8f4d158da9", x"2d5574fd42ec324c", x"17253207a96f163f", x"3778ad6b05337efd", x"12c6636a1a5a09fd");
            when 9136677 => data <= (x"5954a85b8e0c1c5f", x"05ad2b9728bae3b6", x"ca6c66210b79f8f6", x"19500b6fa9ae0932", x"dd3f3b24495f0fd1", x"fe0b4894c2d4bbba", x"c6d59bb6989eda3f", x"3baddee50d692e47");
            when 5649480 => data <= (x"c2d70183dc4d93ab", x"29919e9c2333516f", x"3245f6d81ad26287", x"489eec66a053e47a", x"ecf2da1f9a69eb59", x"5a5252622757235f", x"3c01fa57d0d22ac4", x"8824ebeaec5bba43");
            when 33653821 => data <= (x"af73132e0bd40b83", x"6f224ad00f54d464", x"7c77c73050076912", x"d6c39b5cfc620d6b", x"c4dbe78c8e4265f3", x"ef34ae70e1963664", x"5755a5f3e1c75f4b", x"8b99ddef18bc9826");
            when 33975980 => data <= (x"caedcb785990cbfa", x"770c48cdf322c316", x"02fc8fdbea2603b2", x"fcc7abdcab315ad4", x"872be6b898d7b47b", x"134c1ea204f0e135", x"1158c766af85f2a6", x"6eab98e3ad168bb7");
            when 4861685 => data <= (x"c9e5400e270abbd3", x"8861564e01c7b959", x"56b82326d08f05e9", x"4aa150d523924b92", x"436c7f4d4c4aae71", x"c82514a8557ec0e5", x"75518d95f7bda898", x"519a4a5431205239");
            when 4952951 => data <= (x"ecb08f79eb2b891e", x"11626a731492d26d", x"d954568cf6fb5c1e", x"86836b47c662d93c", x"6e7d8cdebc8cb818", x"1affc1176d0d2dd6", x"e3fe09f08a881ec8", x"02ce387ed9f79c34");
            when 15652652 => data <= (x"2255f80ac5afbf24", x"775dbd823278b760", x"7c164b731add4bf1", x"98bd8ba9eeabb06c", x"8fc84b080eec20b3", x"1c7c22a4d74ccb41", x"66bf76b0381f0efb", x"244c23d8a6ba1fe0");
            when 29131530 => data <= (x"d3c3835c25710d92", x"64092587e1933471", x"b452aa794c0b0454", x"184596c14aadcc3c", x"031e328ceaac9701", x"566feaa9b0de0ef1", x"9076c6240d30b277", x"76d11433664e7f55");
            when 24129039 => data <= (x"6c97e274931a1796", x"98a71e76d63e504e", x"7bc344fbeb6c5abf", x"2be34298eecd8e8c", x"55bbebfa0fa30bad", x"302cf471e5debd33", x"db7258d704c7bf9f", x"be9eaee49e2640e7");
            when 18584830 => data <= (x"1c81ac29b7fda1b7", x"673b177bbbdc833b", x"6e9efd290d96b4f1", x"ed2150013f30969c", x"ad7bd6c244a3cb82", x"6eda364b57e4bd7b", x"7a6adcef8fe54622", x"bf4bb4506fe3ea3f");
            when 22214632 => data <= (x"de46c8b32c9dce0e", x"8dfaf473c2da6164", x"044ecca8c6979d3a", x"dff97d212f20f107", x"40e8acd6309e4ec1", x"b7a9864f39657108", x"1c62afeaea3f02fe", x"9469fc25981ad11a");
            when 13620091 => data <= (x"36758da8e8e905bf", x"ed452a6e040ce3c5", x"46152254e9a913dc", x"b9d29d30329f2702", x"d26081916776a4da", x"fcef9591691d3dca", x"a45c7d89d70a6d5e", x"5ec16d5860ec6db8");
            when 29768010 => data <= (x"fdb24844485f117e", x"947cfcd04fbd42fd", x"07da6d0e537c6985", x"0356a24c6ff693da", x"cb68aad0d1acab4a", x"296d613d686f210b", x"61c8b471d6aa6eb3", x"a0333c979f7a2055");
            when 7990120 => data <= (x"111097c1b2cada06", x"1a0ade092c99d277", x"10411a5583bf9842", x"fb17d72612dc5f3c", x"8e14b2eb86bcfb71", x"828cbb17c33d281b", x"157ff8c6e229f08d", x"484def2b4534d33b");
            when 5956388 => data <= (x"ca62a3fd4edb42a6", x"b03f2b5540bd8798", x"8b83a0bc3dd9f8ef", x"090e1eb72666b356", x"f25e29fdc1625a92", x"fa3ac504ba150d30", x"e5924ecc1bc11dc3", x"3fa438b81d66384f");
            when 32087219 => data <= (x"bc73497e0df51fc6", x"1ac5652bfb3d4953", x"a6e2b894d8837ff7", x"e7e14e63574104c1", x"d2b267b3f4b21ab6", x"e0d91c17ac5a5d37", x"e8e49c06b0c328e8", x"6ee72db6862ab25e");
            when 17350283 => data <= (x"3a70e29daf28e35a", x"63c4e24c866f3d15", x"22492a34b7ceb7a4", x"f5dd5b98aa4286f1", x"a90f967a790d3731", x"9db2e8d425cd82d9", x"17ba7a1bf5e126af", x"9aff69cdfb5f7cef");
            when 16450250 => data <= (x"f1c83239e35d0683", x"01cafc22f15e7dc8", x"79ceaba264edd8fc", x"8ae215030a376a08", x"d233c0f264818823", x"d4b8d9235091ce78", x"d3597e5421f42c3e", x"bde898abf43df1ff");
            when 2146822 => data <= (x"443f35d07fa302a1", x"31361d9e67609d94", x"9a1a382e8910743b", x"89547aa32e6725ed", x"0df5bc062629754b", x"f46f777e9e83b918", x"ea18509b8df550e4", x"ca05319126fa12a1");
            when 9226715 => data <= (x"5fe03217eac22755", x"edf000234aacb4bd", x"74f04b5c635f9893", x"ed75f1fa1f085537", x"952415a97ba9725a", x"bcc182b7f4ba18c2", x"efbbb0cae7d1e6fd", x"de22ddd0471e17f9");
            when 891525 => data <= (x"7465e09742536763", x"2b1dce6308eedebf", x"e1c881ee94369602", x"778652fbb8fe57c4", x"8150cf9d2637f90d", x"82e34bab7f49cdb8", x"99daa05d830ff8b6", x"5b92ac575daa0500");
            when 9896692 => data <= (x"27cdcbabde6f3f53", x"33e37e438cfa4c8b", x"fd23c24b6f09eeb9", x"8da0aea876530f50", x"6b4c586938ea9888", x"2574048fd597180d", x"ff0f5f8dd96ceef6", x"3e20087132c881f9");
            when 31458711 => data <= (x"c482978b1f993517", x"0c721c1a2f8cac4b", x"21fb25df5637342f", x"e3968f6cc9d2dcf7", x"97b835a6c1cb6cde", x"53581f1267f48536", x"aee3cfcd85901901", x"cf27993b176b6f54");
            when 33261943 => data <= (x"6520a0e9c9ff55f5", x"4b3963ee701f8eba", x"6d62209abfadf9e1", x"ee22af1224289553", x"9004ac578f350bcc", x"ac74ce216e16f948", x"d8af1cd9c0a38b66", x"37a0572be0df48ff");
            when 3366401 => data <= (x"a51ce74542f4389a", x"a8997fccbea65683", x"5b1caae722a8b20a", x"70fb80d00dfc631f", x"7f0064c83f7980fd", x"d5065f90b952b5ab", x"9b78a90391fc22c8", x"14a671eb69994974");
            when 5711024 => data <= (x"97a4e37c576d6727", x"f2077f1706bc8d2b", x"0ddb565a3bd43a71", x"efff3f3f57189053", x"79bc31561a81fba3", x"530a0cb3f37cc8bc", x"f2d09f5cef9a0586", x"648c9121475a70e5");
            when 31600086 => data <= (x"bb79b0b616b27db6", x"bdcdb06b99e6ff36", x"be140778d059b519", x"f3f0483872c91a97", x"dd095b96471ff45b", x"cfcc98512e78da68", x"1efcb4fa71215327", x"9d832fbc6666ca08");
            when 30631549 => data <= (x"56c84ed4f29bad10", x"1b36ddb65e8aeaa0", x"57e4ed5aeca23d3e", x"3bb2a72cca26cea4", x"954c22df79685d84", x"727c7f0d9448f1b6", x"5e91e3faa094801b", x"92a4d490652df72e");
            when 21923735 => data <= (x"71385a932a41d063", x"428db154a3a62509", x"b542425eb4f3e4f2", x"be35dad7430c7147", x"b80f48991260cfe1", x"b072e85f9d8137c9", x"f31dee1148a94542", x"0e3f4f08fe758484");
            when 5838527 => data <= (x"aa8e70bbb98da280", x"f7fc9fb85e580004", x"7fabe56894ae8a56", x"02a07b57af62126d", x"765b3352b5d124eb", x"4bd0e0664be66408", x"15582b3d0873a49d", x"0e4248cf00667655");
            when 11339115 => data <= (x"13ffa70471d7a8ac", x"e32b5862f3b214b3", x"d927cdfb50cac49e", x"fd69e0d99b7a9c1d", x"409c92a67552533f", x"b5a074b862ab14fa", x"75f148d63ed07fd5", x"74d8c24b695a4756");
            when 29230697 => data <= (x"dbf57051231a6c35", x"c26c2b2213ea2de8", x"12f932545b2e02e8", x"3a7a414e1a31413a", x"d39cd85bd52093c4", x"2b1b319835b04ae1", x"22cd5ca92103da1c", x"7b408688f2ea9654");
            when 1639944 => data <= (x"0e34933b66805afc", x"d724fb1be73165c3", x"b3b566fa27953723", x"a6b6f2f8e72ade2e", x"7863ffe915cd77dc", x"8dc29ff44ba2fd9c", x"3302085f3d3efc14", x"54e96e83a2e8b677");
            when 2670670 => data <= (x"b1faed16513127a7", x"2c25ae5bef6fff1e", x"8df9f7f9443fce1e", x"60312a0d1c516be7", x"4024ecb766c96fc5", x"2d3d69b5e438d999", x"89530fff07c65d8d", x"dc972c8e803f162c");
            when 24697849 => data <= (x"bd863231e7bcb83b", x"3adec5438a6f08b2", x"503e0b84d3d24d80", x"0500915a35c3db7b", x"80f3acf9820ff2ae", x"c913770179afb96e", x"bfcbba646fadc5c9", x"409b004a492191e9");
            when 13164850 => data <= (x"9c70a9b18d36f87b", x"c18ac9973257452e", x"9f10356ea12ee975", x"94822f5d156800ff", x"242d0492b1922e60", x"26a7f578b26884b2", x"809fc4e3dbd598d5", x"0249e8fe44a36a96");
            when 5780316 => data <= (x"a69e08bb6f25b94f", x"aea9b3130b73f10b", x"85a0e8970add315c", x"77a40c117e6ff586", x"55f0aa1b9e512eb6", x"e73a772e2300658f", x"e3edf4f5877a12fb", x"c6154bafc616cb52");
            when 14887124 => data <= (x"f40b21106ccb7898", x"d8f8e4b88be89b2a", x"6efbf8f518e37d0a", x"89ffd715ccdf0f08", x"3295ceb1050b948c", x"758b8e6865c87b41", x"91c1817818d132e2", x"c4031505425f000b");
            when 32006809 => data <= (x"d5550a48261ca283", x"0cebde11145f74ab", x"6f4cd20d6fdb6299", x"121ad95278821006", x"8d3299ca29c00a21", x"5d8ecfe3aeaca1dc", x"f1e77b43cd35707e", x"6ea4054cb9412366");
            when 17982526 => data <= (x"f8761273904a4339", x"d3801565330e0e80", x"73f5294504031ccc", x"f5ac1d94cbb9b5ef", x"e1e9b1977a954344", x"98b77eed640aae87", x"1316f9b776a1f35f", x"720c5e66092e50d2");
            when 10905163 => data <= (x"e723f352cbb1920d", x"d7b15009058f0b8a", x"d58cf41f32704c41", x"72e1fbcfaeb6fc41", x"5d1058b19551fc80", x"709c71d145ae150e", x"1013a869d9d65a27", x"36780c8f33295bad");
            when 9458845 => data <= (x"fc7b7d17a161e98c", x"406847bd07b2812d", x"5174ef0d16103a56", x"540de7c5acf99632", x"4f90cd49a2bf1cde", x"a2ac279ac5b38759", x"cc0f540f74236af8", x"56adf9e6f48402f3");
            when 21097309 => data <= (x"4a3df6a48364dd59", x"cdf8083af4d16996", x"2ecd6d8d5cfd6ad3", x"c385c3e28e972aa7", x"4cf9ae20662467fd", x"f3d4d271636ddc8a", x"579d7b850c724365", x"9dd81121767179c1");
            when 16471518 => data <= (x"d1feae2596355948", x"5501d32596ae8d97", x"c316c7ee590597d9", x"a36df38c35c304db", x"9a193f9ee2587fa7", x"f80588786e3aa5d1", x"65edd7ab3198dcdf", x"c8a99aca4c0644aa");
            when 15764674 => data <= (x"7b652476967f0859", x"04d9ebe6cdc5de68", x"e88d1bfebfa6cbb5", x"5aed4b8ba58e2aa8", x"5757363a5db78a69", x"0731878c2ea545b1", x"4932d9c01e7a515b", x"99d665a35180c6eb");
            when 13848282 => data <= (x"85d7baa205aa3281", x"bcc616b7b917a6d1", x"6cf7437720d6bd73", x"bdc5550bf4585ae7", x"e26756bb3883d4e3", x"8a9daae07a8470f1", x"d4e0671923168451", x"6b65f5c37feb216f");
            when 15106694 => data <= (x"b737bb0432958511", x"673cb86c058c20f7", x"f34edc70d1023de3", x"5660841f60824bad", x"552cfe9ee6fe1337", x"1d67941038846871", x"5b201e8a3d4d268d", x"ee8318e8b2cd3b4e");
            when 7324128 => data <= (x"6c7ddb045e276371", x"0cc71722660b2c9d", x"159b34405de2d952", x"b222f3f8051b420e", x"915527c3646930c4", x"bd6c0848fb88b598", x"467d062c28b9bd07", x"86a8f13d4641dbc0");
            when 15219333 => data <= (x"0c70610b630be75f", x"5a5b0b38239892a8", x"00d428f18e80c639", x"827e9cab0afa57b7", x"41fa4adfc559b986", x"531a885419fb301e", x"48f8121a58668dfa", x"7758ee05b582d94d");
            when 15988937 => data <= (x"014b2ef1d41a2259", x"ae05acc73575d8b8", x"58147e25ce4f31fc", x"32b8eed894fc7eb1", x"e7dd57892df5cbb4", x"af525a729d454a56", x"a48bc39eb02e6d05", x"7b141687fd759ccc");
            when 13517121 => data <= (x"e4ebce7e3d8eca6c", x"3692e4093c1f3b57", x"04711f260e96555c", x"52611db03abdf5fc", x"62f4174d4cbb20ca", x"06cd2f982a6cae15", x"75e4726929b8715f", x"2b7164ae86e394eb");
            when 1843987 => data <= (x"830e3c5c2b799bc7", x"91dfb499b83cd7c8", x"b9c6f13eaa23bfaf", x"f8affa520c5dc8fe", x"96ac909d37c66930", x"5b093e7da79a16bb", x"834d5ab7dce506d4", x"8e23dfc4b6b8d8db");
            when 21886456 => data <= (x"a72567dc87747d8e", x"bdd69478595caed3", x"31c4d89a8314edc1", x"a1aa6afff339b6a8", x"f9378c9b79d8b341", x"698f644e65d0e3b6", x"66f0a98fa4e42807", x"3c12e5da41dd0c7e");
            when 3397206 => data <= (x"b46659d835717f45", x"2c7fc19d52be51d6", x"567621ff7ff78f9c", x"cf766f712ed9bc8c", x"d01008ccfb478694", x"7edcb79156b25a05", x"21e960ed43307993", x"90b91fddfca08b93");
            when 11101358 => data <= (x"0fefaea1383a5cd4", x"ef19a1e6c9e60295", x"b388c9e2657abc6c", x"17c0927418e220c1", x"006610be1c5710b3", x"27c0a46983f2d386", x"beefeeb93053345b", x"ae7460485484fdae");
            when 25548275 => data <= (x"10675edc7d649d98", x"1e6574a4b8d35589", x"a5a434ed490fc5b9", x"129c46e345e20433", x"b614a28aa62c58ab", x"58904883f0d338a5", x"2cf0c288ec882464", x"fbcd1d9c6377e4c0");
            when 30717562 => data <= (x"7d769cbadcdb8fd1", x"5f08a1ad12cddc02", x"696e35edf5b4ab1f", x"9b952a2b00f34146", x"3635f706f4cca25c", x"568ab56d3ca2457d", x"756128b6fb2f279d", x"5af5c9d8a7c74748");
            when 29062220 => data <= (x"0412153d252043ec", x"1882727e1bc9ac65", x"21191250c0775126", x"877b424ee976b663", x"50d607c67d289889", x"a2e5a53bd4355388", x"d8a28c1df67d55b9", x"c843c9c6b9282976");
            when 23373235 => data <= (x"7c8752d520c825ca", x"6cb7ed53491435ae", x"5d87040c89cac4f0", x"76ac452cffc49512", x"6d30e4fccd998adf", x"8b8ba5a9726f2d10", x"c477b6f31184cc79", x"d65b6f315ec45165");
            when 28698731 => data <= (x"f3da992e15dec42f", x"821dba57539a095f", x"25e5bbc8a173fdbc", x"6187dcaf4c9ec62d", x"50673370bab7a571", x"ddaaff8cc5b7a0a6", x"46908698356de183", x"39ed573b84354ccb");
            when 5483071 => data <= (x"9cb584e03764fb99", x"62099627b75c0f5d", x"67ac3734ce6bc2fb", x"0b2193fd94f48d99", x"0e5f1b9c3abfae47", x"1b832132a91899fa", x"f2f0341734ada503", x"00af9735c433553e");
            when 4991756 => data <= (x"dbb7cc23398fa7f1", x"9ead9638ea3ac99d", x"22a32aae00d3b213", x"5e4e8239c2f4e152", x"23bccf08ef67adc6", x"4e0e2161008ac7b6", x"a70b017b505a35d0", x"328ac3938d01cf42");
            when 20224254 => data <= (x"810c69068e959b3a", x"55731d819acb6c77", x"b1bf9bf62b7f4e32", x"ccc5add10e81c87e", x"a16dbfbbf4429ace", x"121f346d44a32401", x"3e8211fbdb35d8c9", x"0175f43ec85ce537");
            when 27423559 => data <= (x"d60dd9a36f3d337a", x"08d38a8a17bc74a4", x"8c6342dce243633c", x"f50d78e8b1b9b1f5", x"57ea7e2a85db129c", x"06103a3ab876c578", x"2a23021014f54a47", x"efade61bc9530b90");
            when 3019242 => data <= (x"bef7b9f3d162fa62", x"75856a11bd35914e", x"442ff8172ee1975a", x"e8aa4c40252348c4", x"9f8c41aa9b8c8b75", x"273c74916f4be64e", x"bd7c123e013673af", x"228c7e022f03c5f9");
            when 16532021 => data <= (x"8d0d7ad86bdf1187", x"2b6aaa4835a1318a", x"05ef2d104f9afdc4", x"ac0a504dd24a9b93", x"0b5d3bf18833c395", x"6a86b5ac7fd11437", x"0c4bc1433535f501", x"2be04d9ee9d097c2");
            when 4149468 => data <= (x"5c4a95ce4a4ff45e", x"3479e8476e1bc841", x"4520067fa0fe7993", x"1d63a9fef3bf5ef7", x"83fb17b95c8f9036", x"64c9396186022e68", x"8eda11d455b2f84e", x"da8a3c11b6db3470");
            when 7622406 => data <= (x"7956666691de3033", x"c633be7934657ecd", x"6a9478b3394500e0", x"2267ba16719047e8", x"f4c9b8e86f67d998", x"ff304b72774ce11d", x"b8c50872029a96c2", x"6d78b7ae9c554892");
            when 29208799 => data <= (x"09d24ea48341e875", x"4266c725d6e7994b", x"2d3644ff9e41dd46", x"2b7b86d40f195aab", x"c764343bcd3333eb", x"50f828dbefd313ec", x"f697d23e71b0102e", x"184f2de8b8f871d1");
            when 18457531 => data <= (x"b772f7fc02ab7f47", x"c20aab128579ba45", x"9120146c39255171", x"25db926150225f6d", x"d725bfa1200d87ae", x"f1240649996115bc", x"a08f1c4f4f88e080", x"cca87fa62dd217bd");
            when 18169448 => data <= (x"6060676617d77dd1", x"73a02cb468d4343b", x"ce7cb12bedfa0417", x"01bcf3d27882ee6f", x"ccda90a112ede335", x"2404a0b2ee0bf30d", x"8936065ccff5a5b1", x"7404e9007d93d715");
            when 20963772 => data <= (x"a2cfee2355a7f772", x"91d051bc9d0c0c65", x"8cd892827c4d30c2", x"2d7f81c1844275b7", x"5367fd68f485bc52", x"9c3a3f8d5854bee0", x"904ddd8001859481", x"5096c44b2d16dc2e");
            when 23647029 => data <= (x"e9fbe320c483e9ab", x"f72614b7d448f975", x"089395d846a59d07", x"94eada44d4ea274d", x"3bb06c2d7581e695", x"299e51033d3563ba", x"c6d4c9993b87afb1", x"19e3d48e270f1e5b");
            when 13426312 => data <= (x"1a788b66c93d0dd8", x"a3305b1ed564a4d6", x"9038e036edd8a4bc", x"bc51bf2731fec77b", x"600ac9cc46a2e1e8", x"27005dde0203ded7", x"967917ebd84c35c8", x"b51a2ab62fab7826");
            when 27424978 => data <= (x"c9ba90b82b9f2bd1", x"99e31c3fca5980c5", x"fea45da4b2b7d45e", x"620951bcded4a499", x"d2021fa934b4e2cd", x"1908c7bc1df7ef54", x"09e65ce87ee62a2f", x"e5f07c8df67804b0");
            when 4590497 => data <= (x"e4beefb3fdc18f30", x"a9be699cf022f8dd", x"37d88a53c56987a4", x"e9db0a1aa164bb59", x"85193cf2918b7299", x"33d8894be7d32f7f", x"1a6b60131d4c7c76", x"67f29ab54d80c90c");
            when 16105078 => data <= (x"ef3c71f4dc718137", x"d89eef5774b5cae4", x"bc5a56245c6ea57e", x"3647440e5a0f37c7", x"ac7e9481f83df414", x"e717861adee80b6c", x"9ede122e11a56e7b", x"4f67e3c0dd340fb1");
            when 884275 => data <= (x"6966b7567ea87f76", x"e46f7475d36eab32", x"7f96d8e51cacb951", x"64498f7f574b92af", x"d35c1d8ea5cb45ca", x"2e283daa2b5682cc", x"fcbc15b52db27d00", x"cedaf1c43483bfd3");
            when 16968898 => data <= (x"78c25b62e28f8521", x"4ec8196326b102dd", x"bcc28027a8e5c737", x"70b8169d929c89b2", x"5e174f3020c0cfd0", x"b3fc7827d791f939", x"4d0384c275642792", x"8a1012a3e1d664ad");
            when 19569022 => data <= (x"20d11e31fcfa9885", x"cdf29400f2fdae50", x"6b5c600cffa3b5c1", x"ef064ac18e5e0ae2", x"20d2d5e5b836eac7", x"2b8d543060e976ea", x"05e3d2ee41c145ac", x"724fcad38018a092");
            when 3392156 => data <= (x"f44717c72ac28d35", x"46c52f926a8a8f3d", x"e524c123e310475b", x"e0dbf89f966db92b", x"e99aa7448923c8bf", x"56afb4d6d509271f", x"30f18668aa3e5849", x"56dc0b63725452eb");
            when 32914952 => data <= (x"8768f59a35a26438", x"354470a3efe36ae1", x"26a947cb089bd74d", x"7d35377c5a8efa4f", x"2872fcaf03e2ae72", x"aeffcaa3f697fc9a", x"daada0f6165e4e2f", x"5c42f8311fee0baa");
            when 24173397 => data <= (x"9dd231f1eea2abdf", x"86ec307b51999177", x"b6ffa0a3e0c86a67", x"9d1b811ff6fb3aa5", x"9da3683260b83885", x"73549c9ee96279bb", x"71718dbd2e9ab76c", x"02e60daa7c4dc8ff");
            when 28291852 => data <= (x"00a4d266826ddd7f", x"6ad42b413a492745", x"a6af22fe0b9576b3", x"443dbba25bb0d2e9", x"2e11531db1856b61", x"2a3ccf73330208e5", x"9b315f32a904d68e", x"d265356837978f4c");
            when 26023216 => data <= (x"59f5f6f258700d58", x"059a26311c45d4dd", x"c97384b4d9f8e07b", x"de7f1fec8ed204cb", x"78c0616d658e26a9", x"2abe8a573c2211ab", x"be3fa5a06fdca5ec", x"a3cf630e7ee16156");
            when 4075272 => data <= (x"d28c1c85dc108d28", x"b8cbea7b1b0bf030", x"d853f5404c41fa96", x"4f7db0da600f22f6", x"2baca3f7cabe51e2", x"b0f37d095ad484a7", x"c0d2ef6937f454e0", x"36cea2c053bda1f9");
            when 27055801 => data <= (x"7d00ac3a91015e8c", x"a12d5cc025e9621e", x"499a5a9cd3de7bb2", x"b20d195e91083aee", x"24b6522c034e97fc", x"6f3ab61a8d9810b6", x"0549b98800589fe7", x"20bf0aef0b0b00f5");
            when 12384843 => data <= (x"11b6141e880d0c06", x"3d1689b7cb495948", x"4233dfec0f909540", x"b3b67ad1dff5eeb4", x"7c64fe84036374b4", x"d590a0c902bc4779", x"3ba157e1575df28b", x"9e9b2a53ed1f32fc");
            when 31546804 => data <= (x"a3f7102c400e9def", x"8616ce937dce4150", x"45d68244a6451e1f", x"9d4f35af9a6269a1", x"b7cfceb78b30b9a7", x"383a79a1b45a1e3e", x"48e135598d5f570a", x"93aa2fa896742505");
            when 10823980 => data <= (x"b820153b5b5a882a", x"5d2a9e32bd2806c3", x"eebe9cba5e8c498c", x"641908481fd1626e", x"a7eb27947fe064b9", x"f016be542a3df0c4", x"4d2f19fdf70706a0", x"04b1806118e7c3b9");
            when 2044535 => data <= (x"02649e66e0ad37e8", x"6bdfca4afa7c7948", x"30b810a786aef6d4", x"f1b15b6abf4ae00d", x"db54f13d0cc20782", x"ebd7a27734d4707d", x"349b3e4b6b0527d1", x"8117ce38df3d0102");
            when 11911110 => data <= (x"7842ec67988a6ff9", x"f68a6ca28fe9cb62", x"fb9fb8868d1f6b5a", x"e6426ed10bc87b3f", x"65664606d7859935", x"14d9b76fe67b2316", x"fc1f511df57e92ee", x"1b41ee958393c52b");
            when 29378200 => data <= (x"1a3c338c805313e9", x"cf4a2c6c5b485bca", x"4597d9668ed9bafd", x"4548344ea1598645", x"12c46b1a36797b09", x"6d545913a53bc6c1", x"ab48f796265870c0", x"0fa087312d66d121");
            when 22204984 => data <= (x"1b2fa56c9a566074", x"a38eeaa9f61c0259", x"6a4e9be5f5959090", x"fe77a79edf98456e", x"ab7777529cfc0bd3", x"4dbfa7390796dc15", x"c9208b2b1c07d236", x"ad4f8169eb8f1669");
            when 24523405 => data <= (x"c543dcf67012d536", x"e9cbaaf2f7627941", x"dfff5d4266aebbd5", x"fbcae5225df83c91", x"b05d489fa5b8424a", x"876f6d35769801e1", x"2a8c8730a202ebaa", x"eb32410687a313f6");
            when 30009689 => data <= (x"9beb7dc248e75ec3", x"87d2665af7f71dc4", x"4a0cf48c31e755a9", x"1aa62e83f678334b", x"50710523238e4685", x"f07f70d97d1a0dad", x"034ef9fc3a14e7a8", x"1fff1250b35ee7da");
            when 20176816 => data <= (x"832e453bb373990a", x"d98b260367e615dd", x"2818332d4dd8a650", x"bafa065985fb5130", x"3c1a7b11472693b3", x"d75fe8631cc5468a", x"6d476fd1863cd520", x"122fe8a5570ff6ae");
            when 12951425 => data <= (x"b4dc5b058df94745", x"5fdf539a310d6785", x"ae37706919b699e1", x"b4d721d3d8a99800", x"3f1e3d94aa90ad75", x"56b244eea7b15a1f", x"07e5ea97273c1a4f", x"3ce6903ba5aaa0cb");
            when 4032781 => data <= (x"8449cde4526d1e9d", x"504c5a50d2b22627", x"b341539ac34f6d97", x"8aff0cb71cbbff86", x"7fbd2234c0b03866", x"d0e662ac1ca5e62e", x"03f437e904137094", x"d3007a918d3787ba");
            when 8220472 => data <= (x"c140bcafab80cce6", x"d85ed37dda9a72bf", x"cbff6a900309603e", x"a6f3ac145e0f1595", x"fc1915f6ca6134db", x"cae02f0023e30a71", x"669abfde0d9baad1", x"1e94c6a002ec9bff");
            when 2361684 => data <= (x"83ec894cc44b9ae5", x"103f8afad691cf21", x"1d53c53408c81f4b", x"e6236d7271f6f116", x"9eab7564233a4c29", x"d7640705d1fc5cf2", x"d3a8d8e30ce05e38", x"7473376fbc3d06f4");
            when 16134193 => data <= (x"9910d753b040582d", x"04992adcc97e5aa5", x"0f7be54e73581b17", x"dfedea5868d7d4a4", x"e6f896a3567d7e89", x"feaf38ee1b0ff6db", x"07e896ace13a15c6", x"cedc139ee97b26a8");
            when 27942765 => data <= (x"c28c4af57a484e41", x"e35ef2d5e1fd0330", x"6982569bf6f270d6", x"818843ef234282ab", x"efdaa2be2609b5e4", x"4fe91a821fb3344f", x"8b43e60fee0f0b3e", x"b90cca6c13ee2400");
            when 10814998 => data <= (x"8215fb30af60631d", x"42f63b8620352049", x"d9d31b40fae5a8b6", x"6bc32809b39f0aea", x"a77cbfd98233ab2c", x"68957730a79c5b8a", x"cae4f7988e826106", x"542e74104d92461c");
            when 21766259 => data <= (x"2084de7b065120be", x"3673ce12463a1e27", x"e29a9fb07ad5692e", x"591408366087c31c", x"7b45782b226aab60", x"d54470ebb9e21a05", x"78be3adf30a5ec62", x"0daee4f81b8bd186");
            when 33523173 => data <= (x"e19eca6fcae123a0", x"39508a8ddffff31b", x"39572e99f61818b3", x"87990bd77954b386", x"c3a1406c4bd502ef", x"c346b700522d1ccd", x"33a12ecfec2f5448", x"cc6e4dabea2fd8fc");
            when 13375234 => data <= (x"91bc67d23c741938", x"eeb8f127364929cd", x"3b0a62eb295df8e6", x"cba217676c74db6c", x"1e5d3a2739310980", x"29236a73e1b8165b", x"575783a28db87c73", x"1272af3d9cc0b175");
            when 17300920 => data <= (x"63b61ed5a7a1dee7", x"44feb605da4d0fe6", x"6dc37c892a446be2", x"73f7f6df6f24606c", x"9cee686b2974cc9a", x"061c87f5c933574b", x"5ab80f864045fe58", x"69cfc1d47fa3c11b");
            when 5844401 => data <= (x"d5755be070c4ec61", x"d8854f21d4b3117c", x"8e0aa36d83535613", x"ce4f7ed48f7a1a68", x"fb5ce4ab51413753", x"e68ccc6898b2dc03", x"8a52320f0c00a71d", x"3646ace353df7883");
            when 6034683 => data <= (x"7c336c82bf603d15", x"c5d46eb724e5fe65", x"f8b09edda4ac8298", x"af61eedae162960f", x"8275012c09ee038f", x"1d7c09ad861b3353", x"3a27db8d20efd54e", x"bd76dbe62345be8a");
            when 4688476 => data <= (x"205b4c99bc333f22", x"a4c63b65b077ebd2", x"32bb731493dacd7f", x"ba408c838b17c1f7", x"f1937820f6522032", x"ea9bf157d520454f", x"29f21d28338a46cf", x"0f8690a817920772");
            when 8000164 => data <= (x"6536c8b2cc861bce", x"e9cd0970b4d4d412", x"d98747d07de65de2", x"3470a2653e2c57ab", x"c99514316fb9bf25", x"e5a545a6180ba131", x"fbad09f39982b0a0", x"83fe70637b2de773");
            when 4873752 => data <= (x"50a00c78ccbe6952", x"ef456f6c5ad0bd4e", x"0f07f61c9d21d08c", x"4a1d758a07865283", x"f5ca2a1dd3282a21", x"36c6089ea71b04d4", x"04a01b766b9c9ab7", x"1d9257731b9f4986");
            when 15905497 => data <= (x"a8aa4040b20ff2ae", x"e6e589d3a1268005", x"17763fd66c7474b8", x"b5941f87cb854651", x"6734623df1320f74", x"a5755402f1e9276d", x"42dd3fc29d7a65da", x"f652f4ec9029a0b7");
            when 27333716 => data <= (x"c30151a6a2587243", x"5534a204eb0701b5", x"e338fd10cb41ec5a", x"643fac9f16d4d7af", x"edc9e901cadd5f2e", x"74762a002aa55b3e", x"56565d70c84b03ec", x"178c0e21b24e0076");
            when 19228921 => data <= (x"a9e0089ed44e1237", x"bc922b92703e6d66", x"e1616d5bc89695c6", x"a2071fd4ffdab041", x"f85dd65b231745b1", x"df867f29d2d69b7a", x"e741bc29410ec82e", x"4a12130166d5b3e5");
            when 25535632 => data <= (x"00436c8cc906525e", x"27dec9ae4d5dae20", x"8bfbc8cca787e37b", x"3eb088bbf5492466", x"7e7fb6e330ef97f7", x"6a3b13f72bb062a0", x"2899e6462fd9bde1", x"1caa9c45e74e5d77");
            when 4541256 => data <= (x"ae82aad04b54e27e", x"c912a7aad13ca487", x"5e48535813b36f07", x"f21b6ec1225b68eb", x"4a0d095eb195051c", x"41c133b09ddb985d", x"38042dc253aff2b8", x"5013b99fd78afe71");
            when 12342771 => data <= (x"154fa26d48b2be56", x"9b818abd499f6b5e", x"7f574ff2ecca04ca", x"20391970bd34b3aa", x"99d3a29ed7f43e8c", x"acadf227a8b04dd0", x"6f99e08a2c977297", x"d305b550d2cc4e26");
            when 6285237 => data <= (x"2e0220f85e694d9b", x"e224a631f4fa023c", x"cdaa16ca6d1f7a66", x"f60f3a11f18cd29e", x"e9b6afdc57cb77b2", x"568ea0b9c575aefb", x"bccd9771616885e1", x"6a18262ab5250dbc");
            when 24453926 => data <= (x"c14eeb5a3f815f5e", x"501dd05a510c5cfd", x"a84dfc1eee461df9", x"3eac100b385527c7", x"8ddce5225290e8d6", x"450f049640d6a4e1", x"2828c72b5d82d173", x"975442659498d812");
            when 22530005 => data <= (x"baa5221422fa19de", x"d8999e2b34a03ac1", x"1a8e1e64f921f145", x"1a129012b5c68cc8", x"fc4ab328e53bb1e8", x"87066d4283049a8c", x"b3ff2b8e32494c64", x"22f1f45e1463dcee");
            when 30201913 => data <= (x"ee8f5254e574b660", x"e35bb948ee30f16a", x"34576e40d4a04ad4", x"6a0abb98bc33c83a", x"a167b856a091d125", x"1210010004164101", x"deee31c39be63fcf", x"475a7d371da79cb7");
            when 12380242 => data <= (x"3a30387303738ce0", x"e0149e87fad452a0", x"74dffc8539592dcd", x"80ec87cc28da108c", x"017c2d8555dd1282", x"c0f6ddcd65f8799c", x"e8ad01161f2c7e5a", x"7b5c8168f514a632");
            when 14407191 => data <= (x"a7e53f993c16cebf", x"b4792f58771d0ae7", x"5bd17479ea380217", x"f05f1589934078d9", x"a68ad01ce41a54c3", x"579ed553c07a549a", x"9664525c99df4e53", x"92b8b81bdc57d2b4");
            when 1367526 => data <= (x"0ffb1979a5759b52", x"6cd95c1512ac7b66", x"698e732a4d197933", x"118635c3d7a40a2e", x"2cd23470f6fb18c6", x"aea67d2115be61b1", x"e3270010b8a8505d", x"c5fff7ac13177d70");
            when 33087112 => data <= (x"522079a62a257216", x"a3c64f312e81b98b", x"b1e2d102b48a2fd6", x"8ae01e9182cfc582", x"7515cbef73b86e15", x"a9417ecfacb3fe45", x"894678ef2ebf7739", x"f0fb66594cd36751");
            when 23692472 => data <= (x"748a9aa871032d76", x"791ba84873f38488", x"0db0cd2cf2853142", x"b0aa3f9bf4d71d90", x"0017a744c5f6d321", x"f814d3c8bc429ec4", x"3d0ad4060f74ad94", x"2939f08d7c370157");
            when 28686296 => data <= (x"9b085c65172c51ca", x"f545920f14cf1f3c", x"eecbe36f20fa738d", x"cb83f42adcfef4ab", x"34fdfb118a12cd6b", x"594ad1a43d36cdcc", x"a51c92c5773be7bb", x"0f93530160b3b80e");
            when 7633128 => data <= (x"5be82f368d38900b", x"03962049bb4c1914", x"68655f8f4b493840", x"c5d4b986d6c73cb8", x"380a3cf640d23d1d", x"9b3b8a4f9eaa3456", x"1b69d17670f6f6c7", x"a73861fca742e088");
            when 18803464 => data <= (x"4a3b5cada01aad0c", x"7fa2fe51ab3cb0fe", x"3638a20c9336ea71", x"ecc833a7cfc477b8", x"38f5a171edc4219c", x"13e2d386f2b3caab", x"d89204c334742a04", x"e5b6d9c559126bfb");
            when 4868579 => data <= (x"911f0c4b6d1991fb", x"00b614a3f0cee6d9", x"35b31e6760bf0324", x"921a8cc568ac7c18", x"58fd3af0ee87b26d", x"ef8831f7258f3ef6", x"1581b191b3e774ee", x"a3c55152bd0662a8");
            when 25136813 => data <= (x"45d7e896e4f95bb5", x"39c1468e28a62ec3", x"b89c66134a201658", x"2fb285b98dbb8d0e", x"a5bbb9698ed6e979", x"79ed1a51f0f595b1", x"d2500b19d7d2095c", x"4ff7759a542df5e8");
            when 15616093 => data <= (x"2a48d5a460d3e8f7", x"a59c31680e465d5b", x"287b54db305f77b9", x"9863087771f5a917", x"15b103b5b0a4a01d", x"2ff00bc54fa8ad98", x"4c48a62009c90c39", x"49ce36629a3041da");
            when 18456234 => data <= (x"3d64252892101feb", x"5aff5cba01f763fe", x"86e6d3b33135c9e1", x"9a40356100961675", x"5943016d0d048450", x"b246903922961a8f", x"fc678c943d78f6fb", x"f26936cd67b1d6f2");
            when 18021193 => data <= (x"74145b46ca16df9b", x"8bcae4ebbbc93300", x"d14e96c1feef7ad3", x"2d837fe448827102", x"a3db47c65e6b410c", x"2fc85bcbe49f9182", x"1d6be1c062a40297", x"1d1e5458e2a61402");
            when 1960046 => data <= (x"70b95140f626cca3", x"fbafc59ef44330a6", x"fe7ab9142db8a8c7", x"3025373d365ac964", x"31d4a41161d3f30d", x"d536bfea81c299aa", x"c32cb5f07d0379f1", x"aa585f9f33dba14b");
            when 16200993 => data <= (x"46cd1259764d74b5", x"8295c4706f708659", x"294ef248070de6ab", x"fa1e2ae004f7ab3d", x"44076ee7b34f8c29", x"b329926d4e932005", x"76e8f0476ca42178", x"4879281498f91824");
            when 16420742 => data <= (x"ad70224939d93ca1", x"dbe89295a677dbcd", x"34f73ffe5cd925b0", x"1ddc7d3f3681b39d", x"6356d68cc4250cef", x"be5ce63b5c02cd5b", x"4a8c57649578547a", x"0c43731753594597");
            when 28138966 => data <= (x"a7962e2771d3916d", x"863e6a3a78e35dab", x"e696b2e3af8feb96", x"bf3b621d49d9918e", x"a947b07a9aacf034", x"86a9970ca888d1d3", x"97aa44e3b6dbb3d2", x"87a9c26bb297c14c");
            when 4829492 => data <= (x"1f61bad98b77b3a0", x"0324f0b7040a071f", x"7bc814718f1c3664", x"43c62fce931a72cc", x"9591f3bfc7f16cf9", x"73644b9db77d5487", x"5324d751689e35d2", x"28eb2652dcbdd79d");
            when 16617787 => data <= (x"5f0e430713cc5501", x"f499e3046d7962ac", x"5aef382215290817", x"5db1ca2ea0e32702", x"8e2ee0956fea1368", x"29bfacfc6b84d3a5", x"3eebd75403e1915e", x"afb88096b8d8ff1b");
            when 25413973 => data <= (x"89c33992cf5ef460", x"be39ff7d7833bde0", x"deb8e0bb71cb1874", x"810388992cb7210c", x"3fedfc9ef432dced", x"9048f9cc07e959ab", x"68cd12b47492d63c", x"6e62e85d4d0552f4");
            when 7320404 => data <= (x"cf6f54c8ee40d8d4", x"7c093ff9cb7e925c", x"fbabcc19423197d6", x"ca07f4531c0fee65", x"e64e4a1ca9e2e524", x"f8d3afbd13f9dd55", x"9805c35b78b48cfc", x"7d83197ee3cf144a");
            when 22069254 => data <= (x"34d753e5d3ac923d", x"9ce296b1f192879a", x"4bc980d571cf33b3", x"815baa1fc8abb52a", x"a375345aa6c191a2", x"4e5b105a661766a3", x"c857560ede454948", x"f273398dc841e175");
            when 13244215 => data <= (x"ec1a2a98f1d2955d", x"9bd0e19b61193696", x"d82110d23efe74b7", x"ff8b81711868b9dd", x"565541a0ea08d97b", x"53868a75c6b0bbdf", x"b64b2677d5cf39e7", x"f1d909444afd2f3c");
            when 14907782 => data <= (x"ff3ccc5dc83ba696", x"d715f3d220cf4624", x"942a0a19fa1808ce", x"bef55c1bc36b1e7b", x"634a0c3c4f654275", x"919cff943a953b16", x"178368ec3deee482", x"0aa1878cd194e0b5");
            when 30694832 => data <= (x"7deeab1500e28819", x"ee55f909d78bc722", x"753507a595d5a872", x"27e8240cc4a8f512", x"1d1edd3ca24c9889", x"07af75d3a88c0bd7", x"f249aa9537ee9ae5", x"183a6acd74fd20e0");
            when 18306709 => data <= (x"bcd6c5440e599803", x"0e6763abd7f09083", x"296488882c055688", x"fdc18c23e50350d0", x"fe4b7d5156be6079", x"f1f1d0e01a1190fb", x"395b90150bae8ebc", x"3e85d1527778d2f5");
            when 22554607 => data <= (x"8b9ca8b67f89edba", x"4a82f9d42786e648", x"cca45fce60c84afa", x"8bae8b2e35d3450a", x"50a6c3160cc8b42e", x"8b6b79abee92ee21", x"09a6496edb12775e", x"f4cae4efdaf27531");
            when 1266604 => data <= (x"ba6462ea2d393727", x"90168a06891545ff", x"18b97df25b9dad68", x"c9c54d124853a499", x"001a3dfaf89ce581", x"59ea03b6c1f075b6", x"fb30eec3422a61fd", x"a313626cceb0c9a1");
            when 4086523 => data <= (x"dd9bfb7795e57462", x"c9b3489357c6a794", x"a61fad8af7edbef9", x"9c746bd2c5e6473c", x"034abc2141ae0b13", x"1c29ccbcd4ad5619", x"fe4c24514bb5512a", x"e3b723d93bffc696");
            when 15475328 => data <= (x"effdaf4f27a12c05", x"fddcb110bac36364", x"fafffa306b69883e", x"edd73ca0c85b7f2d", x"e9c2c2eb9f46fb01", x"28c581a67a792b68", x"ecc981d91aacf672", x"564f94aba33682ab");
            when 9135058 => data <= (x"d24b173a4a517499", x"2519dd12ac4e6adc", x"95562627a34798bf", x"af5db8e31f795933", x"20b23bace743b5a5", x"722d7ba7fd015493", x"e38f45c4ab63af15", x"8e456acb5b97fbc1");
            when 10255027 => data <= (x"3a0a67707c725857", x"594c765ef89ea0cc", x"6a9aedea87733d18", x"07b410f599629abf", x"cc863a2730ecd531", x"c184834bf4689b0f", x"5f01244d40c4b50f", x"f7f6035222b38fb3");
            when 18613748 => data <= (x"810f9e5b9df93972", x"2d63a9ce32429a98", x"d507f067e328ec2c", x"d32fdcfb539a77f8", x"f11b48c440dbfb3e", x"bf6103bb68979dae", x"36b1a0b26a2ab073", x"a091ed9bc6174486");
            when 15361580 => data <= (x"59a29b4ce2768c4b", x"4f45cea256ef8f1e", x"8a2e0715ada88739", x"a3024d4c743651e1", x"c455fb3169a43afb", x"3bc95d601d6ac001", x"f6edf925a0e45afa", x"213c8e67092f2970");
            when 1370566 => data <= (x"479a5614eb65bb02", x"6e38ef5617e59a0d", x"c24a50440ce1a5ee", x"2fdc0a7a26b47eb5", x"d95019c062b45e65", x"c13a60f5bf31264b", x"ab4cee47c05581d8", x"2545d39e42f750e1");
            when 22396862 => data <= (x"2f2d4a733abf656d", x"bc47a36dbdf0c54c", x"adb1a9a46d228851", x"ac33e81b2d705bc0", x"2a3750a9c9163647", x"6ed386ecab35c4d2", x"bed8298788cb5eb1", x"861360988b5cbcc2");
            when 15952891 => data <= (x"1fdc231ad7fa169a", x"f5804406dccb1ce6", x"d252381861b304fb", x"140817e9e4e08425", x"7728d2018df8c2d1", x"b60d5791e36497f5", x"8069e363fbe920f0", x"85e890edfda6d9d4");
            when 30206187 => data <= (x"37cf65d0411d5d75", x"c9aa7b550fd53961", x"c6423dd759414100", x"dbfca7e7c42142c5", x"661beb3ead7a4d8d", x"09c1a68373842362", x"9a7fbd2900b731fd", x"fdf586d66b2bab87");
            when 5995478 => data <= (x"c0ed0180de931da9", x"0ac6e3b0f44c5120", x"7cfc73efb805917b", x"e6a7ed6a0c3c3d15", x"24cd4c9b7c092494", x"ecb42862dd728736", x"68204878113de966", x"6743a5c4375726e8");
            when 15052034 => data <= (x"473df791a97394da", x"0682eb760e4240aa", x"c39f1655fdbd9d58", x"efbe5a42c16ac09b", x"afded90dcdbb6c59", x"8a6d51352724a4c3", x"32fe19ebf1e9f890", x"f537a1bf74e62c5f");
            when 28782914 => data <= (x"4b8440d30d0966fc", x"ea3254bf01f479b9", x"91c5931a0b472e87", x"b441fc1c470c919c", x"6b6a58645c8aeafa", x"2e7de6ccd0002118", x"1cf601c12ddf1a3a", x"550512c455c9af58");
            when 30037105 => data <= (x"0e3dd5db49ca6cc6", x"59d4ef9b0c8580c7", x"72b4f4bda23fde48", x"6f3568166a743829", x"93dd9ee67e5722fe", x"8497aa34dc3b91b4", x"479f82dcc4392eac", x"1a44d851e8f165da");
            when 19342480 => data <= (x"c2e3d059078ba814", x"c828dd70da9bc3fd", x"aeba41a5e158e864", x"d539b6669fc840cd", x"9052570f2cc2a3f1", x"b1bff5fb8148c3cc", x"156d4cbdcacb7857", x"d40252fcc50a7bae");
            when 12696265 => data <= (x"bf5a480fbbfdf1df", x"b5eaefd232d306e8", x"7bd3b3d6cba7d429", x"f80ecabd73f2aa08", x"c83d9df62dc92a94", x"c7116261f16c2413", x"aafb59a0fc960939", x"dafbf66c204c5982");
            when 24959653 => data <= (x"22df39775f44f962", x"04625fc6f7e302d5", x"a1f1728d41f42cd0", x"f4fa1733f63d0815", x"d300da54fd65d579", x"036214092add37da", x"1abf171089ae0e95", x"9b9a267ffdd26922");
            when 8134673 => data <= (x"e0e17dfea1c36fd1", x"4d4fdf7dc65672bb", x"2149e5e6b3b3cd96", x"843183332423d25d", x"e83a0fc720d80706", x"896b37b548ad53f3", x"982b23f1353b0f3f", x"d1748ef2698727e0");
            when 21433942 => data <= (x"0f8194e317626316", x"b2044cc2512da31e", x"9121a04d1c3243d7", x"1b09fb81ef893217", x"10f51234f3e97006", x"9ae9d24ea7b7859f", x"954aa4e2ac5924e0", x"5d5ad09b749a2248");
            when 19314455 => data <= (x"b7f0c430a2745ee0", x"a2eb4e5963b3642d", x"38494b7c948f99f8", x"8754394bce760ace", x"980332eb1f7ce26d", x"f7c65bbb309b8b62", x"ab9d20e4de45974b", x"d6b6c6430d548c38");
            when 14234911 => data <= (x"04fea7c771ab986a", x"ea75efa338b64bd8", x"126d07c0381c4225", x"c5b04734c56fe366", x"7c195a5b491b4a19", x"4d5f6f06e39fb186", x"54ced07e648aedbb", x"8e8bb2fde5b92316");
            when 3279266 => data <= (x"98c9223524afea26", x"172638cfafde5925", x"ac3eb6cec8365254", x"e8f777487dfa36e0", x"dc1419977890fbaf", x"c5ae7efc87683d20", x"c0b876c21367ab40", x"bc31e7356ae4cbd0");
            when 11323180 => data <= (x"14c338df270e8307", x"c19176f678a9c189", x"48a63300156e2a85", x"52998ba20d109f92", x"2e8851ba8a02c13a", x"85a6063feecc1692", x"6527702c0da6d7e4", x"35aaa4dbb168655c");
            when 14042549 => data <= (x"fd80fd324fe0ce76", x"d41b35396da16bac", x"6a4fad500d49387b", x"d2f9430f57eed0fc", x"2951823a32b3d19c", x"f098921c03a5b523", x"9ff87f3453b5c219", x"f40af55e4b78252d");
            when 1742704 => data <= (x"8e43ef30d0c9ddb1", x"ead8d2a415a6c7b0", x"2a68741e2ee29406", x"dedc0b56227cb53c", x"fedbc9ab097579ae", x"0c9c5b6837f12e46", x"e5ef2bcece75a3ac", x"cba9090a7555e1a3");
            when 14303282 => data <= (x"3cef1bfd8ab834d7", x"ab3f7e69b7030f8e", x"5476aa29a96ac994", x"3ab6aaaaff2f56e6", x"ab9dd8a6e6580e1a", x"ce692b46d309bf24", x"5b53e30aba36156f", x"17cda596738a2492");
            when 9217873 => data <= (x"e932ddb86d80b566", x"2cf06eb1c2ee3921", x"506f2e20165b784f", x"7bcd8b43666d8a72", x"1884d4283494e27d", x"138af7cadde8fac9", x"dee7968380eee8e1", x"96c38939cc8ec947");
            when 7663037 => data <= (x"ee3082f00abf0272", x"9aa81ddaced59150", x"e5bbece21db7c9dc", x"0434800885042263", x"06020becdef788ae", x"b5e066b242ab141a", x"af490f9f37f4f50b", x"09a118fe2e4324f7");
            when 23470537 => data <= (x"98892b1b9abd422c", x"9ec02eaf7dade3fd", x"3bb9077d83ba731b", x"67d59f78d33336c6", x"f4bae10fefb09c9d", x"16dd62c4b0c0e0d4", x"5927666c45d77b0e", x"b654e061bdd6abdd");
            when 8825039 => data <= (x"0bc810aee60ee3da", x"f3c7e9ea40873af1", x"b1931157491fa01b", x"247b980823157e68", x"32adc27eb8017907", x"9e599ef5e360a394", x"675ecc32d381f077", x"5ef6cd087683c6f8");
            when 31745202 => data <= (x"121a60cfcd2debfe", x"eb12997bdb1b9a4b", x"7574d3f691f21fad", x"10385fc3cd47502d", x"9ad37a0fc54c1adc", x"84290ca3a31dc6ac", x"924bb25d5633a0f8", x"383b62b6761a0866");
            when 12953849 => data <= (x"e1f0f15029cc07d3", x"013024e0b171ff72", x"ff93111b7cc5591c", x"c6630c9a0960776e", x"2f0748291e6c36b1", x"c632146a98e03325", x"aa92ea369acf6c67", x"7fd8356599d1e712");
            when 33220527 => data <= (x"4e6edeb1c8355cc2", x"9b4909073fa3c825", x"48bb8755fce6b59f", x"5f8e2c7d116c857c", x"165b4de0622d90ab", x"c68a0b7ec649456a", x"cc7313dcde284050", x"45e6d864b6975f11");
            when 13265375 => data <= (x"728d16adaaf09d51", x"10ea42c8f4b749cc", x"996568498e410205", x"939fdfee7f3b7b00", x"505015458ef192b8", x"5b331f360f1bce3a", x"a15adbb9d8a5aa03", x"e72e0f7a9077a185");
            when 29754290 => data <= (x"d7c1b8153b8e5e4a", x"53fc312bbd284b5b", x"3dcc40b08db73621", x"3acce20eaf2579fd", x"4f549629b8c06412", x"29e7353ebea2d37c", x"b5f15b4abdd2dde5", x"027a22346939d1d9");
            when 12607183 => data <= (x"4ab014b050baf384", x"b6a4775ef4a86db5", x"1a359583333650e9", x"e8cb43a6cc88f6eb", x"c7ccdea846f91a7e", x"bf98a55b217496ed", x"8e40810c6185fd72", x"9645f53e9da393a7");
            when 31024859 => data <= (x"31da354a1b5b5aa3", x"17b9ccf92ba01d9a", x"7e15f9116c12bfac", x"6a4b702e189bfbd7", x"999951fff29cc613", x"b999edb6fafe0938", x"10df2fc7781a1f21", x"92b378658490be6a");
            when 19349939 => data <= (x"b431e7e83c8edafb", x"239ab88e361ad4a6", x"7ce35949a2f8143c", x"42b017634060f08c", x"6b204658fc8952f7", x"bde16a659a4231e2", x"be2ba0d07db3cfb9", x"83a9e5b9d7cabc9f");
            when 32386809 => data <= (x"a838ba2219491ed6", x"86f13e606454b482", x"1e107930c77de0eb", x"900071797f0a8289", x"8bd93cf85cae3bc7", x"983f27c1696e6410", x"b1daf33fef6e1599", x"60f80b7e8fe2070a");
            when 16475571 => data <= (x"b763d19ca2576445", x"29b7d69b13e81ff5", x"1a76cd9ace49676f", x"8164fb255539a3bd", x"c3f3c8560e453bd5", x"bece04396e067941", x"96b48fcf5f10b714", x"ae57612c0bc82ba6");
            when 33226652 => data <= (x"ea2a50e9db1b2438", x"0293020bec2a2c37", x"1750fd5c52f31053", x"610b06fd976df597", x"ac1059e35fe4429f", x"1cd19f4566185ded", x"832194e6e0f22700", x"218009287626d740");
            when 5287328 => data <= (x"a7cf8a9d99eb1896", x"620753ce4decebce", x"e8cb02316503893b", x"058cd2c1513d339f", x"9f6131a4de23a8f8", x"a6b9af61364eef2e", x"922f40eff979e3c4", x"3e5e65ff831a1717");
            when 22712706 => data <= (x"61b5a92cdb80dfe8", x"de55157fbe3ec996", x"5625030ea0fa0d3a", x"0d29abd6f79c5d3b", x"2dc05df0637bcb97", x"d77536d39b826a0d", x"693a4b07e3bc5483", x"f6f7b1a66182eea9");
            when 10147692 => data <= (x"9b9e140d4c114646", x"38418cdf57b2571e", x"0eca33be26320482", x"980a54c0c7782ea9", x"a5e96304fcfbb71b", x"56e5a37b5a1c14c5", x"7f14324efb66bc9b", x"161f42ef7f7294a0");
            when 4915498 => data <= (x"045a5893f3daae2e", x"0d6975e986eef931", x"ed0a369ac63fd17d", x"61be49c997ea08f1", x"337960554008e1f5", x"6d5e1e5febdfe694", x"3dabcb6f899ecc61", x"6399339e72efa434");
            when 23493412 => data <= (x"61475f9e4a534b75", x"cc0fff6ec36faaba", x"39739a309673b790", x"4c47b12a9b15dd5c", x"24264b375bce244d", x"1a2ad260adc13a37", x"ad7bc13871c5525a", x"b1e18d0c3a61f08d");
            when 11905102 => data <= (x"da12ad8e25870f5e", x"f11ae18afab8afa3", x"610ee0f5c8dcfd8d", x"e756f0de5a716d28", x"d4354b04eba21cbb", x"3a5726b070873963", x"09027a52dffaae94", x"328e117b8c7ad61d");
            when 21531299 => data <= (x"8c73b00a588ea7d9", x"1c9274ead0716cc5", x"e018e5f820002fce", x"1efd506c021c807a", x"af5fc291f88eef01", x"5b3242ad18849eb3", x"1b29e60889c91cc2", x"ea95c71856922433");
            when 15864130 => data <= (x"0da9932d6b82ab97", x"f9e0b67939e65e1a", x"49cf7de5b4197e3c", x"c6799818c8219bd5", x"f006ae9e48fb749c", x"10e4f16c5ec15ea2", x"e877ed322671589c", x"63849e5ba1a33f91");
            when 10093809 => data <= (x"7111711201ba05cd", x"81fa4471aebfb820", x"fab495441f39dd9a", x"9e1e03f9b13d512d", x"77097a3d8ba9bf8e", x"5d1494cf9fac27cf", x"082062670bdd76ee", x"6a48759feb619e2a");
            when 29344305 => data <= (x"b3e6db65bbd0c0a3", x"a46f1cd8e3cc769b", x"2dcc2d91833d3ae2", x"98651f55a80cf6e0", x"6467105eae7688d0", x"1f3f2e44ee9080b1", x"0cb628e904c33dba", x"c0a3d8d39a6e9a90");
            when 28859974 => data <= (x"940b0586ff0102ca", x"184ceacfbb0df8f2", x"fb98fc28d16047cc", x"30bdf4736a541b4b", x"2a31fd691444db62", x"fab16418dc3ad777", x"ee8ca1374aab2c28", x"d0f61e076898ed19");
            when 16555646 => data <= (x"c34e5b436123bdb6", x"0d0933f4d18a7564", x"4275242454be7064", x"dea12787bbbdbe5f", x"5864f08104880846", x"b57c77402d2ac139", x"f5e898678dcac368", x"3b5cec38148f1891");
            when 15644700 => data <= (x"890ffc3ef9d5482a", x"795d34c9612787a1", x"994d095929750574", x"0fd02a6bd1d97344", x"86f3b19cef88449b", x"e3784749cc87607f", x"08396660c4787401", x"858e486b6de92c7f");
            when 8963058 => data <= (x"fd6baca64c0f84f1", x"fba39686c762d32a", x"3414646ea476cd21", x"f00b483576a2d7f3", x"9df4fe57b7c9cc5c", x"89b5ee251a2f20f0", x"4c6443ee96294cfe", x"f998b9d6ead694d1");
            when 20539376 => data <= (x"9e9f4a665035e49b", x"0eaad18206786dd7", x"3584ff6c5e71d15c", x"272f506e2cee1bfd", x"9d2f44e3da58d819", x"fbf5e30ac0add48a", x"573e0436cc805631", x"18e51f778f648959");
            when 22524546 => data <= (x"b5e2c5811c6af943", x"67b2ec5493df9799", x"e7cea997fd6d76c1", x"50f0047238333991", x"2aca3d3388e43b9a", x"03ad4e5e91169bd2", x"01c5802215b3d963", x"9326cbf5389220a4");
            when 32380097 => data <= (x"8f633e92fb448859", x"a19f394c5a707e4c", x"16a5c942bae7422e", x"2fdae1aba7ce087b", x"0f65e02f5f4c4358", x"cd1341725b8acae3", x"87ffd1577a40cac4", x"b0a4610e64e0b1ff");
            when 32423894 => data <= (x"75ec2f1bdf3179ab", x"045a8b4d2714268a", x"c5cdba4a4fc76241", x"77bb5a0bf971b735", x"3bb4c735511f8706", x"ade19440007074e8", x"48464ff140de9827", x"c86396241ea3543f");
            when 21557471 => data <= (x"54231d67f30b6cf9", x"25ba69d5fd5f0134", x"ae9dfc8df6bf7b9a", x"6bb66af72625d2ec", x"0f6c17b48cc1423d", x"c1a3fd09a1590000", x"e055320fbb442b73", x"54ab989f138166a7");
            when 10673305 => data <= (x"107a3195b1b80f60", x"9eb79bab077d898b", x"b861b4f7b6c70437", x"236a0296dfb8448c", x"f0d8180ded294237", x"600f7c8dace51201", x"1b00140fce06742e", x"781a76421d680e69");
            when 26478158 => data <= (x"b074e92fa8d885d2", x"a87f949f7564e629", x"207aec69af3609ec", x"47ea4d5999a4100f", x"3246c85bb40cd828", x"9a73101dca992700", x"3fc4ffff5104d7c6", x"61c561e82f32432e");
            when 20043303 => data <= (x"8383cdd665f6fb3e", x"d8d643d9d1fd602f", x"05e720e758b25f12", x"19760f598e6d0b3d", x"97759c90e9967adc", x"016ab02ce16916f5", x"cd95a685f31b7340", x"31eaf81c1b048a0c");
            when 13478001 => data <= (x"c3c697678642b0e0", x"fca31e17786cec8b", x"9644b84b4e8b7cf9", x"22111e3c36a72952", x"89e4bde9d868125e", x"df642d5619b6d1a6", x"f210adb55340d87b", x"1c3c0fca05025f6f");
            when 11623459 => data <= (x"9b42f79f03c9a543", x"27550864d22fad41", x"45732b19720454a9", x"77e775b8f23780ee", x"ecc2bc1172491b87", x"7789b6de60f8a1eb", x"a11c7ec2c35d621c", x"72805456a1889e4b");
            when 26245833 => data <= (x"4f26a2d762296d2a", x"d46e0c8440629fb7", x"2a889994fd9a8f52", x"b4ead9a1d08d6787", x"709c9ac7dcc9f1cf", x"3a379a844c0db7b2", x"8a929b6f4f67794c", x"1b470f4c8748c4fb");
            when 12080708 => data <= (x"e1570251e24e6d0c", x"8a376f263e9b1d63", x"9136fcbf4428a8f0", x"a4f4aee127e89030", x"6414ff8f81325583", x"0ba92aca225fac61", x"3e117de78cdce11a", x"1e5f63cb21143ae8");
            when 31926159 => data <= (x"85c036f14d2c2653", x"f25fe71d8e1edb81", x"a4eff9ca5a05b3dd", x"c4ee94e4dc94e1d0", x"f7d91da1ce140daf", x"7e30d89d38a05d45", x"afd6d8ee3ce7293b", x"b42995d0dbc19136");
            when 11374868 => data <= (x"ae77dd3cb10d1746", x"a32755a2c4a97436", x"b867093b24008147", x"ef71f99ac752b480", x"edbbc3e3ec31473a", x"f94a357ab8f0a6f0", x"d62b7f4105b15e44", x"d5eae2320d1389ae");
            when 22569683 => data <= (x"448bf3fdfaac6932", x"43017b2c9e1d1550", x"36348158b4d833a6", x"f2900a2d1056122d", x"ad00bb6ddbfeac7e", x"b3717e7273a68eff", x"cf4259d7965a3bf8", x"8731f40a5e34dd03");
            when 2217226 => data <= (x"439bb71ee005f152", x"041f96b97880ad29", x"8547e1136e65101e", x"11950f712a536cff", x"e15c738e1460d83b", x"5e0637dedda69a64", x"ea53d084fdde4c2d", x"89729a6fdd577ba5");
            when 8502972 => data <= (x"aef2b9cc48ed663a", x"398667c58eb15001", x"c189c403848c3bd8", x"36a570d0d6fa92e5", x"3c79fe92779009cf", x"576b51ca9749edd5", x"f99d7e6eabf3a86b", x"e5aa9dcea461c0cc");
            when 15784031 => data <= (x"4a0933fc01efea70", x"81a1b04a6af8f899", x"6bdd9a31e40ecab3", x"7f75dd7c74018c0c", x"bcd5853721df95c0", x"4d1843be42bf6b4b", x"ac03cc62f6842b94", x"030ae726dc2aab6f");
            when 2456320 => data <= (x"03e1e2227ab9c314", x"bb3eda6e39d59c48", x"eca6713af4596058", x"fdddfe2de2b985b9", x"83401bb523e109c5", x"388df903af80f7d9", x"d2bdf8299decc7af", x"dccac51529a1b22a");
            when 30796308 => data <= (x"a114bbf62867a96f", x"1089c1292ae934ed", x"13a3f597186c855b", x"20b753771db6de87", x"1168662483e14f04", x"3ae110499897db59", x"ff8ea8eeabb9d71e", x"809d0047a59e9437");
            when 18578741 => data <= (x"171af0475915d958", x"66e723a9294a531f", x"12c39d7b5f73c15f", x"ec5411dbda7e9446", x"30c24dbd14e429c5", x"95bac9d07bf4e3e3", x"046eeecf4d213bc2", x"e9833e02a55ec62b");
            when 17109642 => data <= (x"2d84a25c76578449", x"9f3a40cd671f7872", x"3cd0dc10c3e8cb64", x"c7102b540e2da057", x"0a64c7ef8065cbff", x"9ac0ffa89a55ed1b", x"ac78e4fca2fbc7ba", x"b016241c7dd26646");
            when 34015496 => data <= (x"b562e6fa5b140015", x"74ce6019c8cfd6c2", x"961311d2540a53ca", x"7513d11da03cfd34", x"3a6ea0de411ecdc6", x"c536d034cfd7a373", x"00c3a911f20597ad", x"8bc689c6454d7405");
            when 24892686 => data <= (x"c5f0ce573f25bf09", x"ec00cdb7b4da1d28", x"31421d804e4ddab4", x"77d30ea2dc49a9ec", x"1f36d8357a8358ef", x"6ac65341c1a65781", x"aa26beba66b7ab0b", x"79be0b1d6a5519bb");
            when 6112286 => data <= (x"97f1684165d1daff", x"7d643d29482f6598", x"ca0d81e33e6edec4", x"c158f374967444fd", x"e3631ba319a3a32a", x"642fde8b2f8c2cef", x"7fa0d66cd77d6b71", x"114744e8af3102a6");
            when 17391362 => data <= (x"9a0685407482a305", x"e5b5d06167caf37c", x"665b5fdbaba46c90", x"c9c13dfb7fb4ce72", x"bba7b5f752d4448d", x"d6dce1654f406e34", x"e8a8867bf17c4602", x"0ff93db4ed498e58");
            when 20680187 => data <= (x"1847d1869a9b4051", x"b74a3cbd83dbdacf", x"bd6de6d067594680", x"9a68e3af3edf0f5c", x"2d2afb0f8cb31135", x"fa8258f85668833a", x"afb48cf364ca035f", x"36cb1187ab58806b");
            when 14310872 => data <= (x"9deef7535a905da9", x"2af1cba147f467c0", x"9cbf992f534b8229", x"b9305c4e3ccedb30", x"278d2e7b2e85719e", x"561a5456d85d7783", x"c2b5f49a461753ab", x"0eb893770f8c3d42");
            when 26634104 => data <= (x"be2c9e6f6aadd5cb", x"f68d7014d004be80", x"a0760cd0acd8ed9b", x"eca85fbb310aba25", x"05370b8cd6e67361", x"ecf6822977f5cc80", x"bd1d8e73ca2ac1ec", x"b5796ca492d9315f");
            when 28272998 => data <= (x"68a3d39385d53279", x"6b855d56f59c9430", x"03f35b2afe2cf531", x"67f0ca713cba9aa2", x"978d6e7439c18df2", x"d5efab6038605ef0", x"d7169e506bb3baef", x"f2d84e64d36c7e79");
            when 31534651 => data <= (x"48322156794431d4", x"5222b1b0a8216a42", x"8cb09ae49b2fbd9b", x"36400014f00a890e", x"f90363546fcac6ac", x"fa71952ed37e7788", x"c64243079b1a9a1e", x"e82f60e806264e5f");
            when 4273855 => data <= (x"bb392e53b355ff03", x"071ef646adae8d70", x"32fc66b640386150", x"0f02322c7bb50186", x"6bbf4889d722821d", x"e7ab2fda3072bcee", x"429e809e6a5b04b2", x"1fa9514e69e42b8f");
            when 5437113 => data <= (x"3eac18fd3b71742d", x"feee127ed19c4849", x"5350348488f6c2d4", x"545072b55878bd8a", x"2d9a784492d5e46c", x"2adfd3611afcab41", x"f56f8c914a62c873", x"63e2a5e6b937762b");
            when 16586181 => data <= (x"7ac8d32104f60be3", x"7d8456cc50f0a312", x"d742d49dc00963a2", x"790768a22ee256e4", x"da4ad7f00dbcb16a", x"0791ad6ac0cb2fd3", x"b8a5691bdbcf322b", x"e09845ca7137e491");
            when 18403267 => data <= (x"6d26d9ba46fecdf5", x"a774b9f969cda726", x"3f24387bad59f7c3", x"7906fb66a4888723", x"94184fe7203c1d02", x"117c8e7a64279681", x"89511d6a43c1bf19", x"97dfcb214eea159b");
            when 7122426 => data <= (x"8161bc2a940b1da5", x"dda7826402115f90", x"976f97786c669cc8", x"54c3f154fc5c737b", x"1f8683828c19fe0b", x"f3e712548abcf15a", x"b996c0be9e2ed151", x"7f481613d457fe42");
            when 32085201 => data <= (x"1de28165a8395693", x"6b6d63714fbd6214", x"f51dbc3cd7f5176c", x"b6160d67e1054378", x"7336f594a31c07f5", x"76048211964e5b5c", x"236862349a12ea74", x"882eef0b717f4be5");
            when 18813022 => data <= (x"99befd41ae44c505", x"fdc19eff85e3f2d3", x"76317a24d492df12", x"553b02bc2ba9ca15", x"11559bc40b76deaa", x"3b0eb898cf1131a8", x"238033d4e3520a65", x"440f802234de8d07");
            when 33481102 => data <= (x"ac03378856a2a8a9", x"37ac6d1b5d17c270", x"f42a06ee1c04c78d", x"cc81e33e15d6f688", x"c6d27ae8abd925ec", x"10e203548b49cd64", x"91be6c55d89f5d0d", x"a3a2d2d7f699c57a");
            when 23622560 => data <= (x"47acb72cfcc79880", x"ed3e496993d789a0", x"c1fe13e898598a3a", x"c91d54a4e433bcad", x"3bf4d2ae3f04a05f", x"aa2911b280ffdba8", x"264b6bca75c685df", x"7d5b04dc1645041f");
            when 15009814 => data <= (x"b5ec7461f4387bcc", x"0ed53b9f0ab5aa3a", x"7df7b7c16a5413d3", x"c25186a199505abf", x"6adb44ca0e1e93bc", x"bee8bd8faeca1da1", x"d54b274806f65aa8", x"df58fcc6126ff2d7");
            when 7416750 => data <= (x"71c66fac8bec885f", x"5d0a61e929de55e1", x"763ebbc8edf451de", x"fffef186b40d7a4b", x"895334202a88b614", x"a52c69525bfdb3d3", x"088e7e4ef227db4b", x"0656ba0b719c4234");
            when 18828239 => data <= (x"f5fb02c403ffdd7c", x"b2cb80d89aa8974c", x"9572c22675fc632a", x"17f843bca372305e", x"e9200ecc4a57869f", x"e76ebf77b964477b", x"405efec0db15c7b6", x"9583a8b8446536a2");
            when 4218977 => data <= (x"647188c8bb7be6e0", x"f5aa114fe9b74bcc", x"28998eba9fe52584", x"edb855a9e6cfa4e6", x"8ce347e869549e0f", x"acb381ee401b446d", x"581f7d528aa5f7a3", x"72e5ea19a533d783");
            when 2596144 => data <= (x"6bf9d176feb026cb", x"89857394f97136e0", x"9fd95f8145c91170", x"6546f21758f7707b", x"a73beaaf065417bd", x"ff6daca30cedf99f", x"57acdd994600ddcb", x"6f116e3ef6d24b9b");
            when 19839633 => data <= (x"77d7c7be28277cc6", x"33ccefda8152fc98", x"d9e9a1caa789f172", x"b60eee94809ff0d4", x"473cac33c7f75b87", x"f71996cedb7ea4de", x"6f59cde7d1643bdc", x"ed6d7d88320394ed");
            when 12099406 => data <= (x"ed3ec9eaa755d5e9", x"8d0e8a1bb95da90b", x"402063efcde5ab31", x"a01897766bce9ba2", x"af865fb69f9386b8", x"f97f357c42d614aa", x"a3d06c1c622477a9", x"d48c4479d07a3911");
            when 5797983 => data <= (x"2dd739cbe3d481b4", x"c59c340ed12bcbbd", x"f417ec15e79590ad", x"dd4d94347634a0b6", x"7d7d5d7523911501", x"a0c507b63396ae36", x"9a5352cd0c297e41", x"d3665b3a7f30d944");
            when 6619176 => data <= (x"a0f124906c74de87", x"489285c67cfc9b50", x"b3fa00135896d51f", x"1062d6daa4555dd0", x"5336f32082c075ae", x"aa12731c9f9ef015", x"5d760adcdb0c3af2", x"d41fde8ba916cf1a");
            when 20876140 => data <= (x"1d00f3335b65b614", x"26897d71c8787318", x"2e28355625eca6a9", x"abb186286fdd6413", x"2e7aa16e72fd30a7", x"a78af2560a9a4cf5", x"5e60ecad75daf76a", x"29c4f6c6e001ce21");
            when 10341066 => data <= (x"ea4f62de434e0fad", x"b9bd697c5294e151", x"645e26d458ee2238", x"78ca7d1d612413d4", x"3746050fb1895d58", x"c741f9a000d0deda", x"c745f426ec7c1586", x"930a8d1daa956f6a");
            when 29119387 => data <= (x"cce1e7ec2d32774f", x"4a0f9419116128a7", x"ece6134c3e2dcdc0", x"1c70fbcc61b8201d", x"cedefcde328cd052", x"65754db3549eec50", x"3f3b6e140859e365", x"2629a1d3189edc1d");
            when 29060265 => data <= (x"2d46df6e53b7c483", x"1b8907d7c70ea712", x"2b8d5503430c6329", x"a5f827ed3ff7bca4", x"67c6b9e35b5acba0", x"30b78a7cb710aae1", x"bcbb3cf67581a668", x"e5f91c9f3df2f3f3");
            when 29704235 => data <= (x"b0f4e13e12653b15", x"aee632c943447398", x"b14f5d44e839988e", x"3abc6242b700c3d4", x"75f0d61f8da1d8b1", x"b6fdd85915e54a54", x"df49dd2519fb949f", x"7581f0ea90f83caa");
            when 14411655 => data <= (x"b9393d7372915574", x"86757b222ac326c1", x"14e21011cd9b9b50", x"9baadb65f243d8e2", x"e36545bf6b168f38", x"cbaa36b2df019526", x"3316fe5800b5803b", x"cc1166f62cceb231");
            when 30276512 => data <= (x"7c961f1106a0452c", x"1db5d46d91869f1d", x"3cff2bffa9a0cf78", x"210f473b673e496e", x"95cffeb8cde9830c", x"2828915280c29524", x"a82bc72bd8a324b8", x"48284c77a0e24fc0");
            when 23012151 => data <= (x"2b14995a228762a5", x"49f150cc70699771", x"79e8d1b4193db3c7", x"6a8d5d1e3c6f0a38", x"5b272a3687db4e12", x"ba40f57f9bf4e6ac", x"17fcb9215c745724", x"42751437f5970f43");
            when 20169500 => data <= (x"f60b1f483a76ca9b", x"9799540654297ce4", x"290a50f5672d0b0e", x"e35fcc49dc1b1ff0", x"d9810e06d1411ad2", x"3ca66a8123fbca6c", x"9b8370d7fe64952d", x"3f6902b8e2a9a5db");
            when 16267734 => data <= (x"ad15cce25c676b2a", x"d1bcf0bbea5d3bd3", x"c23c2eef0a7b7eeb", x"8e3865b5766827dd", x"2e73e3a3fbdfc78f", x"ffb550e53d5949c4", x"0e4f277497d8e929", x"5bf7a5127cef9fe1");
            when 22957789 => data <= (x"a8939afa97681275", x"5f8889068aa5d319", x"4904aa9dafe5e585", x"5172efb01b5307d7", x"23797ed2ae8f170c", x"caec9b5f45397a35", x"82bd8ed40d385250", x"9fff25138427ca12");
            when 3091731 => data <= (x"e361b5ac23f89279", x"db8c64cb4d4549e8", x"b184a3ced5ad9aad", x"3d9dc8750d7389a5", x"ac8131080b14b432", x"d2193ce0fb025b62", x"0eac8a31d2ee37a1", x"24e2c8d01a230c0d");
            when 8063226 => data <= (x"9d9c3722e191226b", x"08391c6f3fc98668", x"19b0c929ca7f0e44", x"065b1f135962a396", x"f460c4a8858680f8", x"564ad3058cff4405", x"4678cf38072bd16d", x"3c99080421e3ca05");
            when 33103176 => data <= (x"7366df53fe531e7a", x"d732036e1ecae40c", x"d850cddfe2f6b258", x"e8b31a1ef2629da9", x"d6e2929913ec7444", x"436fedf6d2b76d31", x"0a7aba54b4895125", x"2c14b607dddb3d99");
            when 9704821 => data <= (x"b5201ba774e63ef1", x"df4f18c260f4cd0c", x"461df3dda8922890", x"5ecc595c0986cdde", x"cb1d8aff5e6a6afc", x"39e2b62bf0f8b214", x"c7fe08ff61d81d79", x"dd2e7ee4c57228c9");
            when 9837268 => data <= (x"960bfc70fdba8b66", x"ae8a6acbd6326a87", x"7c1bf604fb2d9ddf", x"b9a1d9d273384a3d", x"1e86febc5e7edf3e", x"0983089871a06651", x"bab1c6c83edbed45", x"d092434019bcc762");
            when 29516030 => data <= (x"750b85ddc9ef04d5", x"932d35443977d3b7", x"aa73c1952e9456aa", x"ad77cfc5548bd4a9", x"b255496ebe7a5f36", x"72a1f6518f9cf05d", x"4a2632384282ed07", x"e2562a4b0cf4f1d1");
            when 14403653 => data <= (x"b62ff36b09a5cd8b", x"ed777a06de6ea16e", x"98f27d2f9745880e", x"2656c82a34f111d6", x"52a6c86bb5a23e92", x"a444347ba282f43a", x"8f7ecc5a19ee96ec", x"a9c54e4c2dd8b5c7");
            when 16744670 => data <= (x"a251c9e3ab4acd30", x"1509eaebc0b8f22b", x"a4c4d90602506854", x"8890c23a73b2cd20", x"19c695caaf68af29", x"7250de465bb801f7", x"5ff8fb81ea0d1eb2", x"a4c36416cf26a598");
            when 32453475 => data <= (x"c97853e2211de5d2", x"2f0e411d3efdc4d3", x"6e1c73f1c7c4bf01", x"8cf47fe370f80a1b", x"a756080a036173b0", x"c25138e9020b6410", x"019e6427e70b2309", x"a249e2866581ae03");
            when 13410983 => data <= (x"e00caf2d10f3baa3", x"73003256a0b6ec7d", x"3645fa27818ee792", x"9c0cbed80b084be6", x"02b38a33cabb2b8e", x"3b19bb1b002d491c", x"4c68778d3d2423fc", x"ff0366b81b9b85d0");
            when 16451736 => data <= (x"d8f1a6bd7ed0730b", x"f798d462db85d452", x"8de70a05192e4c25", x"29bdbe755a8d7dde", x"d865d0f6a9a2c378", x"d54e3068595ae36d", x"a5138ad58e9fff6d", x"4d8121188d0ff9d5");
            when 29216319 => data <= (x"95a2a5049f398d95", x"b0f378aae3053361", x"308b676c8b3c1b99", x"c1e81ef9b102e1e8", x"eb25f01b06f2c2ef", x"0a840f8b3be0573d", x"a21b2bfcadf457e4", x"226e099a0f1f231c");
            when 7255455 => data <= (x"36efa419ef967207", x"0ffd956d62a6a92a", x"9fa5db65b000c24a", x"d7ab3151ac0b912c", x"bc2c0e7006f74589", x"a22b05170950acf2", x"4e7183868b0c0cc1", x"ec1c78d52de44c38");
            when 11320115 => data <= (x"d69379ac1cc38b55", x"a4f3e684e85e417d", x"bece514c0620ea18", x"3dff82cf048d96bf", x"2efdbd944561d6b8", x"b9391527db4284c4", x"8ed673f7870e9566", x"a808fc4976d21e34");
            when 21939980 => data <= (x"826268350d40f38b", x"f7285823f9f29cfe", x"066d473c262bc382", x"25c012a2f18b4468", x"0cf610bf4b59aa4a", x"96ca3cadb5a1b71a", x"01d5f9b5bbe2b0af", x"14fde4fbe21c946b");
            when 7274202 => data <= (x"b948045689fee63e", x"7726a821f4072ad5", x"cb20ef5d921370c1", x"32495da372f51ea1", x"a7dd414c6f1ae360", x"395795a95d3e76b6", x"af6a86f2b21cb6e8", x"4e9d434267e3cb07");
            when 20448740 => data <= (x"b5ebb9f21210e818", x"d920189aa1e8bbd9", x"427cd6cbd33055a7", x"1e7838c4b65757a7", x"7374ff3d6cc1849a", x"77641f7a0c54964b", x"c14f6ef06a49d290", x"38aeff0c1e370bb2");
            when 13400491 => data <= (x"3398b747b591ff09", x"6777d0ab077958e7", x"b51dd05bd8936ca7", x"cc440d2476335bff", x"5cec313fc842ddc5", x"f75089448b24a4e6", x"f9e3845fbf582a14", x"85e951538834bf22");
            when 9884172 => data <= (x"ec782ef09cdf24bc", x"f4e62134249e7456", x"a3bbdf8a3cbf16b3", x"f4a79c8796d6436f", x"70d1c4edc266e25f", x"71a39e43f68def71", x"ecf22e1a5857d81d", x"df4a021eef16f3b5");
            when 26602142 => data <= (x"6f09db449897a932", x"d1ce294c21966f1a", x"9412028ead1dbf6f", x"cda4f18ec358b9ec", x"f5a561f94fb63057", x"fc3c735f83c92ad7", x"5bc697951e7aa33e", x"3f16874a57549455");
            when 14803717 => data <= (x"2d00b3de923c59b5", x"e77bb482c0ac36f4", x"405d337f8449c624", x"1f73af7684c119db", x"a7acf9f14877d927", x"84f304de03be33a3", x"cca38d48f0caa9ff", x"8d91c903c7c5567a");
            when 31599967 => data <= (x"6ee59a64a29e4cf0", x"51a7afcd2b0aed92", x"ec70960b3f8bfc7e", x"3548d2af4a5b972a", x"d385a6dd09a6a294", x"f3b1aaeac6422ea5", x"6de2e4639c4625a4", x"f4b54ad53b4c17ae");
            when 18822842 => data <= (x"d04883b83bcc9693", x"6cfcb7059ed00728", x"e72887a3be9806a6", x"c89495aa147a3ee2", x"6ca28169c4bda075", x"d4c4eed714445b15", x"e039414b39244cd8", x"d98978ece103e162");
            when 22168418 => data <= (x"3d0744c29bed6d0d", x"7f49933a3fce7d8c", x"64033c5691a51627", x"142d8bd4b555ec0d", x"ff67a5f0bf5fc3f1", x"d77730b9b69eae1d", x"ca26663af4524fcc", x"1a2f4efe253738f1");
            when 17653743 => data <= (x"d335cd98cd0a78b3", x"134099259d4bedf6", x"5b562b30c3d93096", x"a00082c96b0f6881", x"ee38f71dc0d793e7", x"7f5f6d8b580d9de7", x"192c1924a582f16f", x"6f1b1ad6718dd441");
            when 9957579 => data <= (x"12881463c1aef7ee", x"be7da4b2d0d354a5", x"f757403be22079f3", x"5b1b715abc291704", x"76032f861136fd5d", x"7562e9e07d67b2bd", x"a1b267c98719265f", x"1be87d3e2b129815");
            when 13159614 => data <= (x"b55ccb0b6eb87eec", x"f8e803ad8e8c2bf9", x"80d9835500ef871f", x"66de245f2e079996", x"0f455d0a08ab40e8", x"4200ef7c138012f4", x"4bcc7f5c26200269", x"1faee13485e4b028");
            when 16082902 => data <= (x"053ecc851e497ccd", x"09bfee4c10ee8ff6", x"11a7b98f26c1a7bb", x"297bc2ecd4e93c05", x"521921a97d40935f", x"db4ce6b66036eda5", x"25130b59f5f3ad60", x"376bae0981b9398b");
            when 12421838 => data <= (x"070fee6438897f73", x"14b11dabdea9855d", x"1d908da5ac4d9c6c", x"d2090c9d9bcb031f", x"6feaf315808a4d43", x"f54e20c0fe0886f8", x"92f5d77d50f84f5e", x"beb5029d26f37b12");
            when 7686587 => data <= (x"4824fedf985910db", x"f52cbeb5e67623d7", x"a7633d36ffb1a5f8", x"2f9824cee3fc3bb8", x"a0ae897233b8e666", x"519a95b84c240239", x"7f1a8c16b3218bcf", x"67394f0f6fb4b89f");
            when 27154190 => data <= (x"15b0a80ff9fe0312", x"f9671356000acc9b", x"6ffa9e06db1abef2", x"c749d251bde59e49", x"dba77ce111d6ba5f", x"7dee468aca705d5c", x"805b0363ef8c892d", x"1a6cd1ac93b461bf");
            when 7037615 => data <= (x"3e82b6ea97cb1d24", x"d1d660c51e9bce7a", x"a9441f818123b983", x"7cd4498db40821df", x"9cbecd0325b2f895", x"a0babee29ed1fa90", x"228d1e79952d2a63", x"032f703cee43d1a3");
            when 31126678 => data <= (x"400983c583fe7e73", x"3a9102554d7d3a9d", x"babe780ca7d79a98", x"f4a13c26c95e3b62", x"18c185ea8e8a5f43", x"85018648419b4c32", x"dc7b3106d185bf06", x"d946a92a4ddb96c0");
            when 20762371 => data <= (x"a6747426d5eaccd2", x"e59b4bf040ea523e", x"107749c746d3971f", x"417fbed34925892b", x"a0d3f8e324a522ec", x"a9953091496e9da9", x"e693a517333316f4", x"49f40607bfa4fcb9");
            when 30107206 => data <= (x"2a9036bbfbd9408e", x"74d3d4644345646b", x"3ae907bbdd9091b6", x"1a72c5458dc1847f", x"8c2d3224084786e0", x"5f7c5361c1c9270d", x"a848c533044c4f2b", x"7f6f5680cf2d4d71");
            when 11157005 => data <= (x"48357732fbf6931c", x"ebc91070eb6c0bc4", x"d32aae8bfc5972f4", x"0c524113cf2b0843", x"8a8b41b5db717755", x"3a343562b675ecae", x"d48de364b73e7f3a", x"3ab02f52d69f06f6");
            when 33662125 => data <= (x"fbecfb6a7fbb8942", x"af524f11ec77892d", x"c93ec0a441cfc644", x"2358fba9e6c04e84", x"297ec2ddd9c1e9f3", x"666a2f69390fd806", x"9341082847e16453", x"0bbc63877e525b42");
            when 14684127 => data <= (x"f3df96f8fa1c5dde", x"9a6bfe9cefd062d2", x"40e001e30e0afad7", x"b311c4554e16292e", x"58632b4c4d3e3db2", x"d2aa638dcc48d69c", x"e81bfe1dfcde101f", x"0e533ca2d2a27f21");
            when 6918086 => data <= (x"0db3f9773d5a339f", x"0c0de8848ffbbaf1", x"4fbe717bae938d0d", x"41be6c713d87c396", x"c15ed80e5667169f", x"a4ac6033cada3f1e", x"9d22e6f4b0591bfa", x"6325f92af32d4b59");
            when 15131279 => data <= (x"67f3b1b1d53f7c4c", x"bcf6a457e84190f9", x"ed250f6eb268b2f4", x"a63092ccdf661618", x"2c0a533df9cc38de", x"e76ffaecf0379926", x"5fc50485e6058b85", x"62b56f94e390349c");
            when 28993884 => data <= (x"5723c58fb86c1a82", x"277421bef345c6b7", x"5da7cb93e22063c4", x"5a1923b131cc7c39", x"dc3d50ff6cb5f0df", x"1aace9822316bc91", x"827ab4e5b6287d29", x"fa3231a2bc8f90db");
            when 12129448 => data <= (x"4b6ebfdc1680b6be", x"aa571c5b4d7acb40", x"ecda24c6fdf28746", x"49ccd0ca563261da", x"8a4d56e5d5cfcb1a", x"86421d19c8d7ae21", x"9706d056d21df4db", x"85b373baa5bd4e1b");
            when 26959919 => data <= (x"b00181c316fce830", x"9e309740c18bb104", x"72fa31e6f66dfada", x"389c38e106feddc4", x"b8a7a41e01f4659b", x"699e3ea7f4bed9c6", x"7e3d7cd0cc0b41d4", x"37bce24459309050");
            when 6533447 => data <= (x"27fb6e2794d003e4", x"e47278d3e9dcf196", x"67931b0609d7c332", x"ad8495d2c18cf139", x"e6e250dd622c0cc1", x"890378026e50720f", x"195c7407ebc6cf3f", x"254cdd28e318e317");
            when 16289696 => data <= (x"23367bf33c1bd342", x"b2965fbfc70d2536", x"006806abe6268f89", x"59ebdf409b754059", x"20178d6195f45acd", x"8543a8631f789237", x"a1e70d951396cd1c", x"184a92b456941def");
            when 14974086 => data <= (x"fa9ad29dfbd4b233", x"965041c43e08f4b5", x"d23fad1aff29fec0", x"1576f0b87d22ec33", x"bba97545505dca7d", x"fba3b40b77dd7839", x"a8d4e289a7054e9b", x"4981e1a7f8333eae");
            when 11284909 => data <= (x"924a34c67af10fa3", x"f9ccd9fb416e245a", x"c58debb14bbdb18c", x"7c4a777b80353a40", x"2ca64f180cac855c", x"51b297b1a8268e33", x"e811827787b99328", x"30b24dec4f435389");
            when 3285706 => data <= (x"c1defb606b4c69d2", x"df126a6a3fe70cea", x"564a3024648cbfb9", x"6114369ec096d2d1", x"95d223d145ab9c34", x"dd203c0c809ad61a", x"b4361e9c4299a40d", x"65d07483aca8243f");
            when 22367484 => data <= (x"f37c2940df3a75f9", x"b9f8a62ff7208f8c", x"76c8ecfc088efef6", x"bbd0672e54daaa79", x"f040290bb57af13a", x"8ff2f58494007dc3", x"f0b86cd9f17516b7", x"866ad52daeb9fc6a");
            when 4190934 => data <= (x"db5e3566327c5a75", x"4dbc1a878a8da994", x"fb0268a16fb17598", x"d8116dfd6f93fe74", x"0f30f8d037d896dd", x"e355607c4f4e6922", x"06f87cd2b8e59513", x"b5dc7f4074cbfaef");
            when 21560086 => data <= (x"eefc18b74227ab27", x"66270a5af74fed98", x"3e3ee7a79bb5d0a1", x"bd3cf82e37245e71", x"138e31bdd8eb8a5f", x"da5f622c5926bde7", x"c29948c7d8486e79", x"4e33b54e9442fb2b");
            when 11787818 => data <= (x"11f74af0a8423974", x"9a94fe1a4509b46c", x"a06c5d2da30ee8eb", x"8aa89d410039f3cf", x"25a95f6ef937fd93", x"fa7b15713f430a09", x"11e1838e38a1387f", x"8b4dd51e7daa6b77");
            when 28951859 => data <= (x"4c53bf360d6d9f8b", x"ff87e23c708469e9", x"ee96389cb9591ce9", x"aba930a0d86b2d8c", x"e979b3c0396a29f4", x"af212b5a8bffe09a", x"c3007445fedd73f8", x"c7fa6e388e28a2c3");
            when 32077096 => data <= (x"c7e41da1d4852a77", x"66286a8d085431b8", x"0c074480a7aecb1f", x"4d8d9674bcb42bf6", x"618f8e1054e540c8", x"58b3bf05ceab75b2", x"97cfd69b98b975cc", x"8ae233f22714582c");
            when 14243233 => data <= (x"060360e0b622f576", x"4ca5b7e8e1e68f21", x"74035eec58455948", x"22dc779ce804ba28", x"b7f81be8e2b9ce32", x"20bae282702c30b2", x"58ccc92d8ecfb711", x"32d93c9d73ae8dc0");
            when 11667348 => data <= (x"190f929e54d49ee4", x"8cf64094970bc726", x"28f5899e5d8fe146", x"8c251754c7a40152", x"eea65d0c46c35667", x"6b420b706ddb5acf", x"c8cdbb5b837fd43b", x"e3704900ba2de68e");
            when 3011716 => data <= (x"fb7ed73fee66a2fc", x"1fb1972c364b909e", x"05ee70cdd135d5b9", x"cc5b8e118225ad94", x"e0346e88c92c63cc", x"c75c70ceb41708f4", x"4a0bba89250a357b", x"e1b0c1f4eb1ea273");
            when 33734919 => data <= (x"72634f04b4332b8c", x"31acca2711a13d42", x"c776a9c9d855c34f", x"ffac930e8ded60d9", x"aca6aecebf3ace07", x"b50f0b357766acad", x"185dae47f472a054", x"2c692c985d5637c6");
            when 1769249 => data <= (x"b9bfff6f0830184c", x"6e1e10505e1a9f09", x"ba0e0ed7fa21a9f2", x"58f1f565635517ef", x"4ed9860d05fb4ca0", x"681f37af817fb7b0", x"a3226185e8b31bea", x"6004b9940f674724");
            when 22429514 => data <= (x"65707aa8213a6701", x"c7e7b7a922c1c1e8", x"e5a7901ef9838f3c", x"d3b146189283b7d1", x"dce4204060886d12", x"95fe2d68e33c425e", x"6c3718b7beb1449c", x"d63b4d6dab4bcf41");
            when 24471194 => data <= (x"1ba713ece2227e73", x"d04d64ab0ce7ca29", x"fc925f2fe911e377", x"00b9972a11480896", x"f9f0f527b92408d5", x"f4872cad1613695a", x"d408fd5a3117591c", x"1168bad989cd8ff8");
            when 20978151 => data <= (x"ab9937b25d7182ce", x"fec27e33674f45cc", x"fc9bbb801226fe4a", x"4f1352d94686876a", x"e6275b2fdd4e4f5a", x"1e3d43cd2bf3456a", x"b5ade6b4951049e5", x"a3e014f1fd041f83");
            when 23873086 => data <= (x"d6f4f5658b858e08", x"d7906d6141bfe112", x"fc63ae7bd84edfc7", x"5181bb91b6c29e2a", x"2cbb0fa456c2100b", x"e548a0e771467d3a", x"8828563ad45edf86", x"19985094dc32345a");
            when 2887720 => data <= (x"5083bcbfb21a5f22", x"299f891dadc48f59", x"f5cf3275a96242b2", x"34e843d6ef0e059a", x"f92509fc91aec853", x"62b0b8d78649a869", x"8d8fe62ff4f29730", x"69a4dcf33087a833");
            when 5521362 => data <= (x"dfebd7b8546e9983", x"c2e78a497ce66b43", x"ff23f33286992f03", x"3cd9c434ccaa75d9", x"9303b1aad3e15252", x"badc7c414eb3b362", x"9eb006d2cc06d9f0", x"f4a146a8b74c26a8");
            when 12637673 => data <= (x"b720e0c3c422fd13", x"7ec71b683b3985bf", x"dd22d7e0eef6dc1c", x"71f69658e144f36f", x"7fe3148c6311233f", x"492c60a3c1c6fe37", x"53c449e635dde7a7", x"6f3ae2dc52c8e76b");
            when 10710562 => data <= (x"80ef2ce63e20cf7f", x"eda6ecefbbd1481e", x"2aa5fbac99a74536", x"786db1b2d1f8e48c", x"4f75d334ecfba145", x"54c2ea171566d95e", x"3184d8f3b91d1e87", x"c80fe73f5897b968");
            when 29285986 => data <= (x"d3f0dd7544270dc1", x"5374fef54c677a98", x"2441781950520ba7", x"af65a1a27dc20559", x"3d81f5dc3c409b4d", x"889104d193125860", x"0833cd12b6beb98b", x"141853eda527eea6");
            when 28527790 => data <= (x"e19d736e3edd2575", x"b2af5404f6e52e3a", x"e18aabefb7be9b04", x"b1b1726e089a67e6", x"27b599f0e2e18265", x"742f39b9414294da", x"c3b2427995945ab3", x"852b517a2bdc5373");
            when 13640795 => data <= (x"db4b06bba82475b5", x"4920496b7ad46f46", x"cacbad6998fbf7e0", x"c2fba8515dd7387f", x"669906b89526f383", x"112a3d6f9a69f726", x"c684cd9f7ab3ab80", x"d46e95502d6c4a5b");
            when 31431576 => data <= (x"55d8279875d4958e", x"e4d20269d1626d73", x"6533c0e465d2b517", x"244c859381de30da", x"314c41397a4687a8", x"79a6849aec165c8c", x"ed6f528e25651488", x"efdb1c62ddd0dcba");
            when 5430728 => data <= (x"2980df01bf4ceff1", x"e3221d7dbe08bca5", x"0c8772700223366b", x"50305bbb6ab06352", x"73832973581976ce", x"728c4dfb9c205b85", x"5c1c27cb6b11df4c", x"92e13b45f00fec60");
            when 2244084 => data <= (x"890ceccb5e0bbc70", x"ca7381eaf625bfe5", x"ea61bef610bcef09", x"dede001390b8267c", x"6cb490b20d07fb69", x"a6ae5bfc9baef311", x"b5a34df4f9ec1347", x"c8ede6a9b1adccdb");
            when 979589 => data <= (x"c147ca3a20a0b194", x"9dca38c586d19dee", x"b72778db9c30fd0a", x"b783308b0a2aa57d", x"a7eccf2fc1171c76", x"75c5919e9d141439", x"2e873728ffc19941", x"1daac5915b7001ed");
            when 18400075 => data <= (x"5f33aedde9b8efde", x"932a5dee5d977a4d", x"82ced05e2d1a45e4", x"90e4068e0b16232c", x"de6b0ef22c887217", x"6aaec18d65ae389d", x"ffc55d747e7a813f", x"5f685629e3ff9557");
            when 7813747 => data <= (x"296c336562cd829e", x"e9ea53176e30f4cf", x"fbfa611d81be9941", x"4aa26d91a0bb611d", x"da94280073ee5de9", x"9c1486db3b4f0361", x"0750d8b1e38d8910", x"5adceb15c2c985d7");
            when 13449633 => data <= (x"e6d5cb4d663e165f", x"1b44138db52382ed", x"87be35bc1559fd1a", x"174742586f425273", x"a7edb49933af0862", x"99dd7622104cc840", x"c1fa6e79e7b2b686", x"db22f02ed714d1c4");
            when 4851759 => data <= (x"ae88ebeb75ee6720", x"3ae4371cfbbb0a4b", x"c5742ce4a022a67e", x"7f556590e5db55bc", x"a0cea270ac7615c5", x"d4be1c0410f50904", x"81454572204f8818", x"edaba04de0611c16");
            when 10143095 => data <= (x"0581054ccb624f15", x"d9f621bdfb72d8c3", x"795bd9a3bc37fc7b", x"5e8f3dedb4ae88f0", x"6523df72e5305578", x"b8eed0a84774fcaf", x"7fcd23bb943eef3d", x"c5b3303e96768ddc");
            when 4924375 => data <= (x"2a7b5f9864aa47a2", x"6dc05326078fb7f1", x"701832dfd669777e", x"b9d33ef76ff1960d", x"795de130aa5a3520", x"9f6772b9db2f8628", x"daaa5589a021526d", x"b7719d7c39039fee");
            when 7169044 => data <= (x"a5e787c615afa439", x"72779991469f3c0d", x"fd0190ff9bcf160e", x"5020d3496d8f4939", x"98864de29b82b00a", x"1a6411d2e2cdf4bf", x"bc8efbe9507ce1e9", x"ce4111f995972193");
            when 25218268 => data <= (x"09823afe3dd1e853", x"e2234ae96c224bb4", x"ebaa7df6099cd426", x"c24a805765f7fe99", x"8717bc87e11ad617", x"f5fd25de2a3ea619", x"d293c8132961fc2a", x"4679fa92e09bfa15");
            when 740528 => data <= (x"48f25cf7ccd64d54", x"ca601e98bed3190e", x"f86519606c926e90", x"9d395ef08c666d53", x"34b7efff895a38e4", x"021bc83866e08915", x"b1838d6197fa226d", x"d390402c5bd5ed68");
            when 15896678 => data <= (x"b4d35f480c360527", x"f4cdb9845fa69b80", x"dff9dcd6b79f0096", x"b42e25a8d5fc7ddf", x"d4e1850e8d9076d9", x"a6aa51941236e4a9", x"4a54d2e05c531379", x"d66b2a3a47ded7aa");
            when 16367958 => data <= (x"a2e870fe6251967a", x"20e3a423e97eec69", x"8f21c9a47572b6f9", x"68ed2b58ac3cc4b3", x"124b11700debbce8", x"6234b3e179206031", x"fc78fffbd3485c7e", x"e436f4d30760f07a");
            when 25999733 => data <= (x"bd17516cd54c80f1", x"30ceb6b3bbee7ccc", x"0f02d52f479c6d31", x"92728d42037910bd", x"600fcda20c2cc7c1", x"3b64c5bce5d3415a", x"b35f251581a5d4e9", x"f1dbad9597b6b800");
            when 3958973 => data <= (x"1f79b8432a2ee39a", x"fbfc9cc1c895164f", x"4fab3717222b8c62", x"58a39ffd97d65ca8", x"99daf81726403a98", x"89ce9105f996eabc", x"2773a4794e939fb2", x"b402be5432a464a0");
            when 21312605 => data <= (x"82ba537bcb9d1173", x"be2afec6ed688b34", x"6ed6dee4cb51df2c", x"82c0eced6e25b320", x"8ae9ca6aedac6ba7", x"08e34bf7b6ca625a", x"b983a95ff0151e0c", x"1ac95eb9799671ea");
            when 23697530 => data <= (x"d398cc23f8682834", x"5e3e4c0f3b93fd78", x"de320d02f737b057", x"8f5ace5c8056aedc", x"21b401c3c0f1f9d6", x"573c987956ef00bd", x"9ce0f2dd9480f478", x"3de92c3f4032e621");
            when 13127019 => data <= (x"37d4bf62b4008cb1", x"25f4cd39c80cd9a2", x"db33e16935b583a9", x"cdeef913225e9bbf", x"6758840362fa091e", x"f5654e9b9cb14758", x"e1b666697f0da17e", x"7636b9508fd3d382");
            when 29576971 => data <= (x"3d276ad1e11bba3d", x"6a853bb38874cb45", x"baa9d40b2745b449", x"a44e9525a8fbae01", x"84e44fa7d6b2fbca", x"810f14f8d44b9b3d", x"bbb1151342e2a01b", x"15cf6a33b2c3fa7b");
            when 29285903 => data <= (x"b472ca444eefe66f", x"3f1998dd2200ac5f", x"339956460a250d5e", x"ce62e76e8024f6de", x"3f1b0b91dc274a0c", x"f20d694ee67d1261", x"77a1172ed5c07240", x"6c2af4d49aee7fe6");
            when 8499017 => data <= (x"9d8fe0084e713fd6", x"84ddcbbb30e63947", x"97be896e2a5db3af", x"bd7efe918f4a26b5", x"49f16115aa8faec2", x"8f3ba1d068c4c99a", x"b0096e5a1eb77ff2", x"11e362076a8fcbe6");
            when 11091617 => data <= (x"30fcc8dfc7e8966e", x"f37702ea4126fd7a", x"0587f4606e2a4ecc", x"cddccbb6b8af0a49", x"4ff5ee600bcf9150", x"4f7e1a60675c694c", x"84c285c9b4ad8a4b", x"2a4c07904dc11cbe");
            when 7712050 => data <= (x"dee57c723af48ab8", x"19f6fba1c58dba42", x"60f279f35292d874", x"269f4342e28b2531", x"55eba7cad91d3aa8", x"dd0f6558be9050c8", x"58faae493b3a1db4", x"ec03fab09ff4aa9b");
            when 7013847 => data <= (x"042f1baa35b90ab4", x"98ddf8c22f9ff825", x"f86e2cf2efa5c88d", x"89ca451c864c4aea", x"904a1327432fdeb5", x"1e3d10da21eccf97", x"1d79e195fb5a96c0", x"cfef412f004da1f0");
            when 10149160 => data <= (x"e5b0f259d8e358c4", x"bf69fe7a1919b4a0", x"9178429d5e9b49f3", x"6843c135c422ccca", x"9fe3a9afe7cd46b0", x"bd9db6a4d5abd83f", x"66cc03d992f320f6", x"e43c321452192eb4");
            when 22035462 => data <= (x"e53ccbb132b6921d", x"7901e13185577681", x"f536dba446bf8cd0", x"b1a6ad9b200cc50c", x"a32ebb3457f6c563", x"85e3488133c57b6b", x"2b40f02445cd02bd", x"ed655554a1818fbb");
            when 9319664 => data <= (x"58f36c691962e74e", x"b054b77b1158cc83", x"4503b24108d7b034", x"6ffcebc5764f691d", x"8e6b6db0179171ea", x"c1a71f60c59ed40e", x"3d9bf0825fc23c3a", x"cfcd761721f2b5c0");
            when 2855247 => data <= (x"541a916938c4fa87", x"2de0cdba29ee0133", x"1dc90faba8950cb6", x"bc62d7ada98d448f", x"7fb473e8ed388ade", x"5ae06ac92afed25e", x"2d5b2ddb1bd289e1", x"dd617a7ea6e2b859");
            when 23267745 => data <= (x"4caf8149ec8162e4", x"8cd68f090fd2134d", x"ceb63bf2eaa59090", x"4e03ef5092937be8", x"3ba3671f6df7ab62", x"2d4a3be6e141574b", x"6b1d8ca194ac9362", x"d18d110bd600b6cc");
            when 20518449 => data <= (x"96a3ac240e0093a0", x"ecdf1dfa7cc73b57", x"a120e4125fcb7fd0", x"60e899a102a11430", x"7be2771f4257d28d", x"41bd4e96af67b7e5", x"aa2ef424731d5a3e", x"d9e1c4d28d4f893d");
            when 4825066 => data <= (x"4ad33b47dacceb91", x"75d86f7a52dff2cb", x"be5189b7583f1d5d", x"afc18aa6a71d8453", x"1380d4506de167ba", x"158ad9974c5b584a", x"4b7db3e501d25435", x"1bb9b1eee32ad9a8");
            when 31505276 => data <= (x"9564a6c2bdc37ff2", x"2612b84f57817889", x"3aa1a5a3619a29e6", x"126550108b1b6e4f", x"4162f5a8a13a3109", x"d0126edd1bf89671", x"93d24c63d20a5158", x"9cca6524ea0657fb");
            when 1840282 => data <= (x"16e1a33725c56f2c", x"a943341190d6534a", x"cda6c3f776da6899", x"75b61762c27c55b2", x"0415f2eeb6c81fae", x"0441fcf3c797f8d2", x"ca0035a4e243156c", x"b1455365e35a68ba");
            when 31514576 => data <= (x"bf5152acb0a1da0a", x"fa3eaf26dedcbb71", x"0c90a3889f9232ed", x"81c132e526c677b3", x"ee440c3580aec0dc", x"bf64085042760db4", x"2de9abc4e3dc21b0", x"f337f9b4e2568843");
            when 9857182 => data <= (x"e9a643cd5f9888bd", x"87ffdf958f638744", x"d7a5e340b1bbade4", x"cd26de260cc804da", x"b9401b43c1c86657", x"2ec9880a0eab28ac", x"81826df52587e7dc", x"ecb99e906851456c");
            when 2349977 => data <= (x"a8488ea336efdf7b", x"23296d8c9b4ba8fa", x"6dd4df652e7989af", x"579e3fb74c2a4ff5", x"4b74514b8e7a56a3", x"a12243afdb2f007d", x"9459f651c2246b5a", x"594982f3a3c7d90d");
            when 6073964 => data <= (x"69d04aa2956467db", x"5b3e023e7e94d8ee", x"123d53ee01dc2866", x"4db3015d1f2d55b1", x"2c7a012ec8f1a46c", x"e5812c19f6d4ed1c", x"957be39f3b7cad42", x"11d515df4431f19d");
            when 32492204 => data <= (x"5f6e73c04617cdee", x"5caca102fe700a12", x"c2ff92fdc3f67292", x"268f9aabfe77e722", x"b3ea37175cc80c21", x"11c20a7bb5897c07", x"161918eb272adf0d", x"bc48cdb950622329");
            when 32127119 => data <= (x"5001b40a886b2e9c", x"6b2262cb864885f5", x"aa499f33dd45feb1", x"7a923a014f5eadda", x"b468271cb2518cc2", x"81c895d24de3cf5a", x"9228a3adbb5d207a", x"1364bc7e055e96c6");
            when 19580806 => data <= (x"9b38b04e9f1fe706", x"c248fbc331162276", x"46586a85636f996d", x"f085b98efdcac72b", x"d1f6bb4a0644fa49", x"fd7f6abb2e942f5c", x"5d4bfb57e4ef6a57", x"30c24fb90a5c7c70");
            when 9513681 => data <= (x"ae75d951c5cf47e4", x"78725a29c8ca9ecb", x"d14bf6502f628492", x"43a7824a8b521258", x"2d37a923133950fd", x"3aa761cefe55e8d4", x"f725e7d6646983b2", x"7662800bb3426943");
            when 28480073 => data <= (x"c04fe708ed629533", x"10d94346ae13c0aa", x"0246107fd8673ad5", x"4cda0c3d5d6dd42d", x"25d4a9d338f98adc", x"ddad44962a21c4bc", x"f4acfb958ac8fccf", x"6e978835be8d30d6");
            when 22005533 => data <= (x"a097efc1c69ee6ae", x"717580cdb32a1434", x"4d26b06f037e4767", x"9d0fdd27f9ad4b5e", x"942430ed17b6810c", x"a5e317e14c7825f7", x"db5436a4c04c06ff", x"73b85e290c0bc747");
            when 29850628 => data <= (x"7b8c8d239fe25eed", x"3383e8bde505ff36", x"75db634525eba948", x"98290dd24faddf51", x"413d04ed3d74dd83", x"714e885bada9f4e8", x"8d46426383b85435", x"1ed6f8786b145f00");
            when 8876261 => data <= (x"a7e7eb2ec152e637", x"40870f074ae52c81", x"86789f5a95df20b1", x"27b90caf3d8299b0", x"494a26de0368a0cf", x"5a47d2b1da7a654c", x"eaeb05e81280739f", x"807405c0b966add0");
            when 16985486 => data <= (x"51ace3334ed35265", x"85df9bd6012d26e6", x"3e7b3c61b98b79c6", x"465ae4d1f103cb26", x"d344ab9b2b7ee91b", x"459383fd6035cce6", x"f62719f988bce53a", x"178f131d8826aa54");
            when 28469022 => data <= (x"d486a33c6e2bd447", x"e29d44c73193ad2a", x"2f90c54802647465", x"71c23134f286f52a", x"a87a549ae1d581b6", x"225f865ec57d29b6", x"fcb420cc9711e8f3", x"8b17959943159311");
            when 21111056 => data <= (x"a9432a24a5c458f5", x"1a331fe49d23ded7", x"d2cc0f133b53ce9a", x"0345cc645cf28443", x"e644a372001c1e8e", x"c8d79fd6214653fd", x"68c923718daa350b", x"67a3e2a79f6533f4");
            when 3847300 => data <= (x"5ddbbea3ede0baf4", x"c1f328d7d565bcf8", x"3b408d038d2b98e0", x"461e545c52ffc3b2", x"bd13067751a13c61", x"318127fd48e2e290", x"34048f2103435b8b", x"0de52f35e5280b80");
            when 23480585 => data <= (x"ef47f0bec9545ec4", x"6b0f6d07466c9394", x"8335e3d6102c4cf2", x"583b80a103269df7", x"ca2909c99321c901", x"e2d792191e028908", x"0e05a0646d0c17b6", x"f197e3aee6d51a62");
            when 7588133 => data <= (x"ad62a91597ec5afe", x"c03e382577691248", x"e82ac9155ad7009a", x"2cd91dded4e195bf", x"1200899a03ec55a9", x"49913de3ae850a2f", x"76ee4bb6f4d403f5", x"537694cb2a5db9ed");
            when 25117457 => data <= (x"b03af6d442723f62", x"aea9c673b62a257c", x"999d2860e4f8d063", x"af3237915aaf7855", x"8f209ed51fc2ca4d", x"058976a4a004beef", x"47124e7c19aa6226", x"2abd64eb8d53f3e7");
            when 20059016 => data <= (x"a1c30a4f652823f6", x"c41a4c9890b7a708", x"2650d6e786141478", x"dfa6fc1952c0ac97", x"bc2735557cddabd9", x"9b8ed7ec2411eee2", x"6bf191eef362ab75", x"4277584fb872ceb8");
            when 28807013 => data <= (x"2cc84658a408b913", x"b349a58aa4d0885d", x"a6916bf76d52081f", x"cfd75edcd291bc88", x"8859283e85dd600e", x"86d1a5433f6bb287", x"ede1c71a371580ac", x"b4c1145ba3d7e0e1");
            when 31355360 => data <= (x"2a3b3802d58ebb7b", x"9c968993e7de749d", x"4f303e3bc8fc7159", x"4dd9ed98e9809e5d", x"fd3ba0802b6818a1", x"49e0311eb750a9af", x"035ae3af2e8cdfff", x"352dd0cb27f5c558");
            when 19002190 => data <= (x"03071d854687c0dc", x"8fa7e04d7b7639e5", x"e15ec79f93031fdb", x"c795fdcbd6e838ba", x"c7c4d23149c25b86", x"143a19ad1785bd88", x"a6f51bec3f45123a", x"3e826f3aeaea2ba7");
            when 23950315 => data <= (x"c003ef4896fc10c5", x"d915926081efb30d", x"942766b490d75b99", x"54d7ee4ba8ceb301", x"466bd8a0ab317be3", x"2959a35ea27fba38", x"900a961bf1be4b6b", x"b815855a625b9698");
            when 32902233 => data <= (x"af6492c792b2316d", x"9e81e16bfd2ba03c", x"a91155501d9aaa62", x"dff79dfa9e1903f9", x"18c4eb98a74a04c5", x"c812ad2040ef2274", x"b428a2b409e5052c", x"78b7a44207439b36");
            when 10350121 => data <= (x"65729b8d2be88a89", x"37f804b90006c390", x"5557e2bea15eeea8", x"f84640382c9a82f3", x"e9ef288f9667407c", x"0d356ae82c9ea04d", x"ca045c105c78255b", x"29150e2c2c809e51");
            when 18870746 => data <= (x"ad3f8940bd8e7787", x"872a807b578bcaf1", x"e68d2472053f0557", x"864ff4eda2204795", x"7d9e96eb70afe6ba", x"a5cdbe8b3948bf09", x"34d6feae0b187b1d", x"34095f2381535d7d");
            when 4708015 => data <= (x"98b0fd6649ac2039", x"89de50aa8a07d3ba", x"f03451d553977b5c", x"fdfcd077bed35533", x"c35259eb25206c05", x"1bc72470c4f1917b", x"cde053da2e969dc2", x"112f786a4f93bc8d");
            when 15799817 => data <= (x"5dbcdc8f7b46bf93", x"9ac9d04fcf08bdc9", x"915d80b3a8b37594", x"5da40e2d8d60a7f4", x"07ff173d98118113", x"1bd825dc0a369838", x"1537ba588f468697", x"f78915ce040326ce");
            when 19155462 => data <= (x"8f6eda8c3a6e2d9d", x"c27a57399f64321b", x"0b13312e34e1eacb", x"0ecf509a344180c0", x"dd2e5c582ce65ce8", x"c1a9cac153b565ed", x"e7c5ab864039775b", x"17d96b7999ef1532");
            when 14669200 => data <= (x"a7b4238ec97471aa", x"068d6252c9d3cb7e", x"bd090dfd5bedb5d7", x"97c38ac6ddddacdd", x"97abe946f2b00fdd", x"8d18f8acc9881c37", x"86ef6c5e7e33989e", x"154f1b7b5050ed37");
            when 24768911 => data <= (x"54f38d25c5d6b3ad", x"011c1ea0fe92c2a4", x"6b99916c23cc5b24", x"bbc58f66885cca77", x"dc3800329c487f33", x"714bb081b395dd59", x"a1091d1357a55a0c", x"0da6d6c1ce423b01");
            when 20729274 => data <= (x"03fdceed5b3cceaa", x"4c5776be550d92e1", x"121368bf42aa8179", x"615c7e3b5946f21f", x"a1747848dd33235f", x"5bcb440cd8d55658", x"1a5f7cd91c819c7b", x"f7d0625dd6fa340f");
            when 33145523 => data <= (x"27416a8a8d3c46f1", x"731919870dfa703e", x"95dfd54365953492", x"fba28fc5cca02dac", x"536bf92495be8375", x"0cc454e9ea2255d0", x"a82892f2bffc79dd", x"234374c2a87e7754");
            when 22058273 => data <= (x"c9c0e6b3118a9fce", x"517618aa10431f7a", x"c009b11109c7f54e", x"837bb6d8d2ebc276", x"be8dc8a8c1d158e4", x"c68d7d2af7331b1b", x"7fa81039c32bf4ab", x"454980cd0f65188b");
            when 3937737 => data <= (x"f7467467152ed138", x"8d888e6ec6305176", x"7122a54109864c49", x"3c6e0d3fba8445fb", x"e6b6ab0d6f3c2aae", x"7297d8a31741ec83", x"349a7cb68d4d052a", x"5e1b683a12caac7b");
            when 33221252 => data <= (x"274eb4a44135bd05", x"98e92b7316731ae8", x"d25db23542295017", x"a84b8ca7a948407d", x"12f871873234537e", x"fecd611a246bd9c6", x"b88526e0fd21e09f", x"ebe8f5672fa9a63f");
            when 851388 => data <= (x"e734466399f199e0", x"b10ff78c4cb9ddaa", x"6c47f963bf7fbc8c", x"900cd80ad956e899", x"c040cd2331b1720b", x"0af5a8d49a2051f0", x"b4fcb6fa4dc890f9", x"48c9008549073010");
            when 32944897 => data <= (x"af913fe627f4d02e", x"4782fec068acacf7", x"97119a1619344931", x"b33cd45ad60c0040", x"db194e663e134fe2", x"2956cfe8c18824a0", x"4ed99bb765065e72", x"0fe2fd7741639ddd");
            when 20000561 => data <= (x"f1ef35bfbd052853", x"4fa6fe633a9d2be2", x"4a5b7d30d533e4c7", x"93175ef20877450f", x"0902a4f95bd5f4ab", x"23166538b1becb04", x"9f60f033ac6c9a1c", x"3f49e52128d3557e");
            when 15573498 => data <= (x"d5bc0daecb9c7d5e", x"cea93f6a810005e4", x"7a041671b429ce2a", x"f3fd7adc35abdadf", x"2a20c0a956c35b48", x"af65621d0b7166e2", x"ecc9bc093b4ed799", x"86ef563ceb127f8b");
            when 1943290 => data <= (x"07cd9c62f891cdfa", x"02943d99ca420436", x"2288808ff01c66a0", x"bc9f44ed8227072d", x"391fc27c6a3a02cc", x"37924c2ab405dfcc", x"4d092ddbe01e68c2", x"83394ae7eb435cdd");
            when 5883303 => data <= (x"12c6de3ded3c7c97", x"87d8df07935b458c", x"e1ac3293e5162ac0", x"97638877b0d83a9f", x"c00ed56de7ac5253", x"6b8df3f2ff2ec55a", x"db2531ecf4190350", x"c8f1344c59d05c0b");
            when 17736410 => data <= (x"53ef53e557fcab20", x"b62f9c202bbe528d", x"a80d051f9944e289", x"a9e4123d5850f1fd", x"c56a9222c564912b", x"866b2dd761779727", x"d90ee54cb1b60aa8", x"d80df53e263ed792");
            when 11787849 => data <= (x"3499ab4217cec774", x"0dd3084c01aeb81f", x"4aeb190a43f9fa59", x"a07c1a0ce6e4b1ce", x"a5c9519c7e28c19b", x"717ec647186ffa31", x"68298f93ccdb8c14", x"1ebe93f7ff190a8f");
            when 11156532 => data <= (x"ccce907c54e5ef36", x"22cbada49a8a47e0", x"d47b9ac0a2a0942b", x"e151c0bcd786243e", x"29a292e401a41628", x"3f032e2939f72d3e", x"90524016095cb57e", x"48d9ab702654e18d");
            when 18062819 => data <= (x"283c39f0dc0f5bf7", x"53e1b12669241ed5", x"f1cb08f2b21bc00f", x"40e5d0d84f38c387", x"bac471ab76b4f2e8", x"9eac6f18dc4b3510", x"6f0046e45fabdc19", x"f1a1ca74ee72fef3");
            when 30964807 => data <= (x"95691e64c49ba87e", x"b27fe9890ccca07f", x"8e2d828fa8c56168", x"b481fb7b311fcdb3", x"3aa7f05368e7b458", x"e67384348e648729", x"56cf6fce1183b4f2", x"299d352f2f6ef096");
            when 30855557 => data <= (x"7feb0bbe9e8aad33", x"b80613667009e387", x"983d482a8699c48a", x"370a48ef2444899a", x"f658b7d31472d262", x"9e1337b08245e429", x"3313ebc51beb4580", x"26475b9363afff02");
            when 3191967 => data <= (x"73fa0dde497e580e", x"30ab8dc5337948ee", x"539926975fa8cf58", x"b25563a2e6c4d30d", x"948f2791e14302e0", x"1cd3991d00c674c0", x"594b29826fce841b", x"a12d516f8a1d28d9");
            when 30998827 => data <= (x"6524f511162c4edf", x"2f87fb88c0928f49", x"2f0ac8084318b9a4", x"77f66df92f5cf0dd", x"307f4d5b4493bd7e", x"ecbb956dc560c6d0", x"ec790b74bc688b57", x"e2eb21867b61540d");
            when 26080193 => data <= (x"22216d2bd5329f20", x"4e72cf93986ddd3d", x"2cd659c6679c1cb6", x"d46af1acde46247f", x"edd8d5ee1e938b38", x"ee4730418f7cadb5", x"0abc38bf3022f251", x"fa2400c4b2a5eafd");
            when 5852997 => data <= (x"6aba45aa9c61e295", x"6af130d80d000c21", x"55ca20d7a7a0f8f4", x"679ae1c8a4def2e8", x"74bedae9536e602c", x"edc86b91ff3a45ee", x"80b37c24d73342b7", x"1fe97d3ffd69868b");
            when 27022856 => data <= (x"beb845cf64a5c5ef", x"0a76b9e07bcf1001", x"8a1cfea1fbd0bdfd", x"a9751b2ec6245b62", x"dc4e7d57d1447b42", x"9870f726e8c2b806", x"8af4ff7742cbe491", x"36fce2b8c9b43d44");
            when 32487387 => data <= (x"aa3b283e7dd8f867", x"fa22d2cbb4446210", x"bb0e05d1f5e69107", x"e58baca5c188dce9", x"df6f4b8ad942f0da", x"2d61807f91e77ff8", x"a1d369afffd223db", x"de110d2fdaa2598d");
            when 15872984 => data <= (x"d86c3ae63eb7045d", x"ad510b11c67b474c", x"6b79744bbe70d152", x"0e8750ea17d1fa99", x"94be311d5cb0de48", x"1df1eed93a95dac8", x"93f52a29383bb9fb", x"9fbe6f0f771fd7d9");
            when 18909860 => data <= (x"418ee3ee3c33e2ba", x"5f24f2fdc46a84e8", x"7a5e9e4376157d72", x"791cc1334e3c85c5", x"0026b731671ea71f", x"ca09dec34566ea8a", x"596120a85d972eac", x"b72864fb1e3f7bef");
            when 15416495 => data <= (x"ba4b36e249c79d70", x"c71b22b9e6022a54", x"60ac0e10a539c17b", x"adea9f168d66d2cf", x"24db330c51f87502", x"71846a8400c92ba3", x"2752d0b7fa2c4d40", x"5fcec47352f1573e");
            when 22530058 => data <= (x"b020efbfd503e907", x"57ac8f3dc04f6354", x"3d6a6c4b992f10ca", x"0dc8b9d704751880", x"88a91df6b5480fc3", x"1d5e5386e66c5eac", x"44ef7f7388349e34", x"f3d6d4ff180f47d3");
            when 28304890 => data <= (x"deef75fa6c638722", x"e2361edd04ec8675", x"7957654bc2398e66", x"c55018ede66ea34f", x"c0de88b125baa787", x"5405fbe80ad9a80f", x"dd4242a38a36ab5f", x"9332c841350c80b5");
            when 4014952 => data <= (x"093a82576b10d249", x"46fa753061d2b256", x"6c86739f3fe16ebc", x"5935c6fe51d08aab", x"0e52b6fd14e66ce5", x"c49a1e80066c3f24", x"157330c082e0bf00", x"56d9da11ec0e5f5f");
            when 5111362 => data <= (x"d9fe3ba67b874e95", x"7a29702c5d0b2835", x"dd926d2d876bc965", x"efcf6ed352ab6a95", x"a7c5b23d7ba47d63", x"e43d8279a327dd23", x"6b266dabbb3f0e22", x"cb500cb2bfbe6043");
            when 5264696 => data <= (x"b28aeca07d575ab0", x"6883bcbf1007c49e", x"f8401b4404788db9", x"a2d7de103161161e", x"741ada7fd8cb5cd9", x"72429349bcb978af", x"35638166cbc45f1e", x"2e45532702a818fe");
            when 22803138 => data <= (x"05af032dd92f6606", x"b2c52e4dd85661e6", x"d1025ba684d64273", x"c53002e430f65126", x"44f3c67635316c62", x"62ca3a6e2a7323c2", x"9f70e4a9379a4c1c", x"7a427ce44e29b828");
            when 33308408 => data <= (x"672ecd3e7b8c699d", x"fd82a2e6c23193a4", x"4420fd2a3b23bd8f", x"7e89b6e27094b12d", x"cfbf759206f891fc", x"6ef3233a8e771209", x"f69021d39b930f0c", x"875a266f98c27876");
            when 8266994 => data <= (x"2a221dc79c0d95c8", x"0329ae35922a6dd4", x"59804e79a832eed0", x"01ea08470bdccb25", x"bf6b58349c6107ac", x"b0ec0b217dea7a77", x"a36a25e3126f8567", x"cf1996ce00cfe4e8");
            when 13349905 => data <= (x"768b270e8bc634bb", x"94c68199c263cf5a", x"51c58f3ae9e990c6", x"6fc9f2b792d86e1b", x"29968c8d8e2b3960", x"529b01bf1e6f0ef1", x"f62f755d170ab48a", x"a4398dfced4896b4");
            when 12419678 => data <= (x"7cbb6f7e8f975d9e", x"fccb62e9f1bacc4b", x"63f7e0453f9c32ff", x"e083c26c9f4f7e51", x"4634ae9f9333c6c0", x"78e26ff7478de749", x"ccfc4714a39f81b2", x"991388d9ac8723a7");
            when 15993039 => data <= (x"a043a4a63b227dc2", x"ed4b04d62b5cf80d", x"cecfa3f40d3952b3", x"1633f6618f7079c2", x"1d4be04fe4db44b7", x"bccbbe632d03d9b5", x"299c02168abd72c2", x"5ed5ef48b72087be");
            when 6841564 => data <= (x"eb8d907646fb8a42", x"13409bc8c8280226", x"cb36dfca14269a41", x"a5caa836e5085cfc", x"89845cd87330bc55", x"5b42ab01e311985d", x"356774e5aa5dfe81", x"2ddd427e2c9af549");
            when 22848924 => data <= (x"02b9acd840a9a916", x"fa816629ba44bc5e", x"5179c1d323388054", x"ed4475a3a24b3e46", x"95894ae150fe521a", x"19af183b54e6b195", x"5b5704766818350f", x"48a47a52af19727c");
            when 16585219 => data <= (x"8d51111a7ae3dd71", x"1c74db1e4d5dd59c", x"2f374b118fa30091", x"0d1a7b72eb389123", x"b2ec2ca9745235aa", x"7f67517f200b52b0", x"9d6e3ac1531b0aaa", x"8726355374d16f6f");
            when 15289404 => data <= (x"4380e9c0be39e263", x"6aaae2a6f06e22e4", x"8e68a827a717e9fa", x"b7673d526982236c", x"4b552b2d1178124e", x"ac57ca655f9d2c1b", x"080647770133366f", x"6f995884c2dda550");
            when 13655197 => data <= (x"0a95ffca6760abfe", x"a26758eeedde5e93", x"0473891476cf4bc7", x"16c6fca8efcb575f", x"aa4a7f1a57fd69b5", x"44391365ef30d73c", x"ecb79fc53600f306", x"c7c098de1864f934");
            when 30613746 => data <= (x"50e49cbb6ba47d48", x"8fdadd00763d1ddf", x"45d06348456645c0", x"dabcceee0931ef09", x"1aa29c3d2907e2f2", x"d053a23f45898058", x"26cba2a65f04c813", x"256f08a723c98b7a");
            when 12616077 => data <= (x"33c6925ed5e0c5ce", x"d0fb2c89e60026c9", x"39c47b3683e66cbb", x"4ceb05b27ec46043", x"aad32a2c67e258fb", x"d679b10c64617765", x"28256ab11f9c29da", x"c3aaa676a28963b5");
            when 12846767 => data <= (x"5f095d59cf18c701", x"e61fc9c817f1b319", x"65dc32f7470da9a6", x"a8c6b7b2038b9f1e", x"8f9e42d21de389bf", x"d714800624997afa", x"e5cade452ce995cd", x"7d4d30cb50c1d3b1");
            when 17021564 => data <= (x"7b5654dc4b316514", x"0417ec16a9c5e207", x"595a8a3de598e594", x"6742e6ec5da7c451", x"821f1cb7b7fe57c9", x"6f24761549d33e14", x"bf1ece0560d302df", x"788ce65749ec612b");
            when 24717943 => data <= (x"68fdd67f0020f119", x"fe017c85aee53997", x"016893618e7965ac", x"b770cae09955eef6", x"146a0537c93b2076", x"216b1e7f138b1541", x"ed492cb078722ea3", x"e78bd062e1f9ff94");
            when 32855996 => data <= (x"e71e381334da2c23", x"f1dc8689a5393ee2", x"63733eb437f9abee", x"bdcece7600d5653a", x"15a6c9f492999079", x"8d9c8afc139df763", x"514d4e7a0c3f55d5", x"10b6d302b74a4fd9");
            when 9933692 => data <= (x"d95843d3d3d21028", x"c52ba530f75d3246", x"1ccce60f10ff2426", x"03b5ddcb89d8b9df", x"357af8907fda47b5", x"b0f73b30935e38ba", x"5d09b09d87ab7f06", x"861f84692d39ff50");
            when 13080776 => data <= (x"d2a1faeec2e23d55", x"824a425352b2b5de", x"d81c9bbc8ca4d59b", x"e44e72c0f8157951", x"c2fc71bfff5d40f3", x"06204700fb8653a6", x"287e48df89d93858", x"9cd1c53b33a25d7b");
            when 14013778 => data <= (x"c4851d4f447cecb2", x"dc67fb9e7c7e32e9", x"49e0bad2b82bfaa8", x"81883af45352dfa8", x"65fdd50e5c0963d9", x"ba899d9e916a3759", x"8d68a7fa1c795d2f", x"b3352b7301b20506");
            when 21726657 => data <= (x"458bbe77f9e74a0d", x"c163871f94b68f3c", x"86de69003148edbb", x"150fa8882b5be70d", x"59851b70631e133a", x"e3daa564817aad67", x"21aaa583a2a20394", x"1c040da2e60750f5");
            when 29432957 => data <= (x"fa3f2eb145a64527", x"ea2be87e09f73cab", x"0170b3d4a8f74284", x"c04eeb44499e3684", x"f963cd1368fea75f", x"68e2e9bdbd811343", x"d1500d6f33976f7d", x"594bf1ebbb419770");
            when 17860669 => data <= (x"ac708094626f475c", x"9a84cf0d46f8bbf6", x"88e1eca8c57f3bc0", x"4360d520d919e035", x"9f5d63960ee912e9", x"5500f15a6c899e17", x"ccfba27f548215e4", x"0c3d2d0127db8a3b");
            when 10912611 => data <= (x"fe8a5d46916d5cf1", x"889158fb0cb517fc", x"999cfbdbf6ec6d56", x"2a3c763fae8b924e", x"33e32d202930b892", x"de2d907fad353cb9", x"d29bc0c6ef155a2c", x"3b09642ae5c8d43b");
            when 5280942 => data <= (x"4434803ee1f9cb80", x"a27feb91ccea610a", x"c3aacc3072c66e4b", x"6e5cbc9f188e6464", x"dd41f796e7d4ef75", x"8aaa7677f50a7a30", x"48825b7fba363279", x"168180b20716a1cd");
            when 10316887 => data <= (x"d4d8834997eee169", x"b1c581386a36eb20", x"387182b65138cfae", x"447386ebf8ae1ebe", x"7cc638d5a3f7faba", x"1936f135b30af254", x"a5db7afbde76bb1f", x"5846c5e1f4d78d51");
            when 13069124 => data <= (x"2896e49723c6087b", x"8f1ee337193224fc", x"3b3da1ca610fd629", x"d294a2ce28a3b1a1", x"63b63fe202e3d577", x"9805027ba6be83f2", x"9a5adf03d02d0067", x"86f1628e8541a7c5");
            when 15072788 => data <= (x"91f1645c97ea538c", x"71335f66fab0dca5", x"fba1b475f2facacf", x"cd0ab9fe1e6fb997", x"33e77649a7045f93", x"8384d3591905ed23", x"32579ef8f2af2543", x"d111f41f165af0f2");
            when 24656425 => data <= (x"5b47c27c00431a2b", x"3bf952a222aa282d", x"2c76f342fb7f3fbc", x"8f14e3940881c5df", x"877c627c62a4b66f", x"9a4f81da4fb1f624", x"8da842f3ab5d0a5f", x"664e4b84e49ccf1f");
            when 17427866 => data <= (x"8b71529cd5be3b40", x"ab82a4166519ed6f", x"31ffcc5dc2e21b0f", x"78740e87fb07b41f", x"823b23612b087404", x"155ae4b8fd3c23bd", x"43e45a8ac45fc9cc", x"3ed90f4e608482b4");
            when 33947927 => data <= (x"53c0fdec3aed983f", x"ca9454c1b6efd2d1", x"18fbdd049f416095", x"647f4542a215aa9d", x"0f600a926d6126d6", x"27e425b3e9477724", x"80b530bc5852e4d6", x"a670c04153e549e7");
            when 20146111 => data <= (x"e314da99d8e73adc", x"3a5feee951990de8", x"1fd9e369c5cf53e4", x"fabb37ed7f808006", x"85b9b1de5a8423fa", x"ecdeabba228d7b06", x"ffa92188d6c547a1", x"578dde5428a98f52");
            when 10682777 => data <= (x"0747304cebec4a4e", x"774b4b0b5e91db0e", x"b8f7632fec664cda", x"8ebb96dd2e8b7192", x"99a62730183476e2", x"576fd7399b903fc5", x"e5fa7bb6f9b90fd1", x"237b45801db39a88");
            when 23469256 => data <= (x"521d9362d72ed132", x"3a2b7014b3a066ef", x"9d013103613da041", x"e5fec3eeaf29eef0", x"95a40f2ba6c24ce8", x"9b25a98965ae86ef", x"32bd64b10d9c229e", x"8a9b7a4639995a62");
            when 28552828 => data <= (x"1c863a96a26ec203", x"08610bee63b54fc0", x"f52ac9623edde276", x"fb4afa8785d93374", x"b144888779fbb9c4", x"772fded549303939", x"dfc9568006b8054f", x"f7b0cd4cfa87b179");
            when 31458648 => data <= (x"0674db9400a1e0fa", x"296dab67ad6c8b90", x"7b7335375a067e20", x"d8c691244c2f41a8", x"89ebcf77b38abbaf", x"34b7684453cf9c8b", x"93beeff07aee374c", x"c5e90433e86336f6");
            when 15189132 => data <= (x"b258d8b78e9d6aa4", x"40b793d8e060ca0e", x"fab38ff2d284911e", x"89c7bfa7bef8bd43", x"0c4326dad783cd4c", x"d989a4440db88d2e", x"cd5d7b6c0c9d432e", x"bca236b196488e86");
            when 22639536 => data <= (x"7d78b391d6bfd003", x"0129df18b5034d5f", x"d505bfc28c4734a5", x"a9b6b3374169ad2e", x"bb47cccd89310256", x"fb107fde89ee07ac", x"28fda228e97461ec", x"ca1a1d61b339ea27");
            when 30782675 => data <= (x"0a549a5d02eee751", x"a503df752d908282", x"604ab188c8b41dae", x"140b6dbc7046d193", x"1da89665f2dd43d2", x"ac7b823ce1f75ed6", x"4fa3621363da931e", x"c58972d856faf2dc");
            when 12962474 => data <= (x"9a673dd9538195df", x"6ed0d87bfe45a9da", x"68eb08c08d9e6ff6", x"b9e7b1a9040ecc4f", x"57edc5ff798292a2", x"437c1b1d788f3292", x"f386c1bc480a1f7b", x"16f3aee93ab185e2");
            when 5084622 => data <= (x"dd92a0dbbacd0dee", x"327d0fe239e01a22", x"3757de7f14412243", x"f28c777afc71efbb", x"8877bb93feb9cd0b", x"d700a985a31b6856", x"168ca122205bfcf8", x"611f1c284e0cc142");
            when 18631203 => data <= (x"98e8204a1eab5874", x"4877e8477c98a12c", x"0e0cea09826f75c5", x"cc6c206a0d03e37c", x"714b29282c4275e1", x"cb49f368bbf17a45", x"063dc46c69f057a0", x"50a4f57c80880c5c");
            when 19601086 => data <= (x"f418dc171c6b116e", x"01568a607c0f62e6", x"b6ba363e923ce724", x"f29bd72cc42e48fb", x"30eaf96b39787c3f", x"634d54c00c1d6228", x"954183097d0a563e", x"f15996663e96f302");
            when 32359559 => data <= (x"43f0e45b663ce9d7", x"a2352f3ed7bacf47", x"2c1c5f3d69a3e345", x"c2335e3bfb036c30", x"daee6eaec6c9b6d5", x"d627b1b1e6a8124a", x"3d1c95cfaf141154", x"a64165741faf48f9");
            when 8231682 => data <= (x"c55ed35a7f2779ac", x"000e0d346f369c54", x"9a69b931e08f7976", x"b7d7164dbee26136", x"ef4dd1ec6b07b886", x"6b5e77f3815fc89c", x"03fedca207608590", x"9e2b2123bd994126");
            when 14882299 => data <= (x"02ec3175a3db9cc3", x"06431076b5efa8a3", x"ca46c8327336cb5f", x"8ca1a19fa720d7c8", x"d3c0a9789aa2e410", x"db2b2a2a46b55eab", x"ec3b82ec60d757e3", x"4fadcc77f06a8ce3");
            when 1329372 => data <= (x"935b7282f62786d6", x"973a3d68127f3444", x"f8244e763bd9459d", x"875913f7b632db64", x"e9796b44a78c025f", x"6acaadd5d599cb36", x"447bf9af3ff97252", x"7e3995e214c75750");
            when 18177298 => data <= (x"07f87137ba7a6fc2", x"468dc8b80ed68b1a", x"ecf392d9534fec9c", x"b753269d8d8d3966", x"80d1e87fe2c44aba", x"c202f877ed9e6fa8", x"abf76feb7cb0cb7e", x"c65761a57d298055");
            when 18648742 => data <= (x"1d06aef8db7ee821", x"354498566a57bc63", x"23b224d0c9745c16", x"29aaf6d569956427", x"05be95eee9493d26", x"c2ae52afd8ea7516", x"a0edbe11c4771c48", x"c5591e8843a2b444");
            when 30311722 => data <= (x"db44d29c42b78272", x"7ec3d249ef6bd128", x"5c9ed2dfadeb73ac", x"eb12abc9587258b9", x"c9d7695261d855b2", x"ece2ff57f6c5e0fe", x"1253a4347da16cbe", x"1125cd084ac31c52");
            when 21480946 => data <= (x"dc35a2aa3870bff6", x"1730b159be03b042", x"7bf469d3d26eec31", x"bc80e7525d50ded0", x"0f5455ddc08b0379", x"79dfa1080be466bf", x"6ddd681256e88a11", x"be7b5be752d2aeb5");
            when 10923644 => data <= (x"f0648ac6f38c92d0", x"045aac4ab4f4f923", x"1ab9eeb0ec05bc3b", x"4ffee43db0850496", x"e053e2b3f42fa9b1", x"67ed41822adeef2a", x"7c6a9c792f4898ae", x"aa1cdedd9cff76fb");
            when 33566704 => data <= (x"7e50db4d61bc3715", x"b3341ad712199e7c", x"bca568a46ceb2271", x"c0bdafa927ae87f2", x"35a41f57d6d7f02c", x"cf6cadce89e6ddcf", x"8e6d287dfd5be801", x"8a927da4e0bf4b45");
            when 20155681 => data <= (x"5ca73e6ff1913c34", x"47c2adb5cdfff0ed", x"1b5aeda9037a7a5b", x"73496a0305a2c5ca", x"797642a6e7c25493", x"d21db688193972fa", x"6c66ed6ee3f1b443", x"ebe970804c332c40");
            when 31963829 => data <= (x"7cb00ec0906bd221", x"b536f11567d48ff8", x"945e1c9e541dffe5", x"a1bbf07fe066660f", x"eb9de343570b76e0", x"adbc51dfe062e0b0", x"f882be18f5a4b937", x"55ff4bbdb2875f54");
            when 21319252 => data <= (x"b924ae4baf4768da", x"ba6839ec5c6df4e0", x"e605fe24f8b03c38", x"dec4c53bb7458637", x"5292b0abdf4684a7", x"924c5c6ce87cc4e5", x"41752e91a8572257", x"1dc1dca18308db47");
            when 27969834 => data <= (x"b2860f0b1c0c26d1", x"8efac1098e0edbbd", x"c0fa304ab281bed6", x"fa7b33a3c9680652", x"2e52ea8478e28d08", x"93caf588fdc7520a", x"345cea871d424a75", x"971bc9a371c257b4");
            when 23569363 => data <= (x"ecf6f1a73f43e919", x"a534e1429d51a2a8", x"a0d4bc811c9e0781", x"b7101ee03dfb5ffa", x"23f4c40c3ecde4d4", x"6b3a99f0182d69b2", x"dc2f07235a0cc1c2", x"11e956e5ca19d67f");
            when 18722742 => data <= (x"2cf6d04149d0d7c5", x"548c218c63acb3e7", x"b6f20d3a6e6de0b6", x"266df357eaf63309", x"6978d82739cff210", x"5eb4d035d6154afc", x"42809f288ca65967", x"830120c5b9f656bf");
            when 22944070 => data <= (x"715815432e565fc6", x"704eb89a3fbc9c37", x"41d8db9f8fe957a0", x"6266758cc83dad80", x"a59c68248fe4ae06", x"4883821e98c20760", x"42173f6a403d2c43", x"2920979c502cc292");
            when 15629998 => data <= (x"6f207ed109e82c34", x"c8d08d224d2a0204", x"6ef95550e7a79f16", x"186fd97b259742e7", x"123f60169ba26913", x"72c07c09318b779c", x"596e180dbf550158", x"3529115d9ae28670");
            when 33752253 => data <= (x"df6468a8671cb7ad", x"c3ddbf7ab4f357b7", x"dd2bf8a6833a94fd", x"2bd05f89a8feb704", x"11d9e4302f60bea6", x"52458ab5d2dbebe8", x"c213b57a7a30b96d", x"e2b76a10ae042569");
            when 10993435 => data <= (x"bb4465bd8b95c1e2", x"9ca3ce5c244e9062", x"fc6020ba7627efc2", x"a6c948a84160def4", x"97f6ee703a687912", x"24a3a3d453248605", x"33c72a675f4de4a5", x"242277815c797cc5");
            when 8821284 => data <= (x"bbf5e2f57ac4dfd8", x"d7b9169c3e6fac3f", x"251dd49848d07709", x"728be8ffafd6aa07", x"c6c0f61b8232c5b8", x"800450c7f57cfa7b", x"adce5d161a731205", x"f74cb097c51d915e");
            when 33018684 => data <= (x"e9902d8d6c1b802a", x"8821f72f6bd1b9a2", x"b215a70aab89e11a", x"4de5e22dfb7525b0", x"adcde104c46344e8", x"298479254435fb4d", x"aa19cba3b1b29ed1", x"b9426a1945e48cb0");
            when 17615149 => data <= (x"b3eadce83cdabb15", x"f5338cc280bc6852", x"173490367c48f0fa", x"2974a83f4acd5384", x"e9e444ea137cd4e1", x"602333764e623899", x"35755ffb589073ac", x"7c07604f75f5cedf");
            when 22594623 => data <= (x"6757d84f5eea214d", x"3bf89a747fd4122e", x"513960a27aa4a2c8", x"1ea6467055eb78f3", x"726e5a36e644b6fb", x"8713212b5c449ec0", x"9464c748ee41df61", x"ecc7bfcf1f21adeb");
            when 21531302 => data <= (x"b1b91ee452393dee", x"80dddbdd6c952a4c", x"99cd5e466fc45131", x"c086aff61a371992", x"279669ac658acb79", x"ee6126f3aff673b5", x"c9d7167304db74d0", x"e58862fd76a5f551");
            when 13959026 => data <= (x"fd2c0286c44fb675", x"e0578e159d717090", x"430f012d23b50f29", x"8b53e1aeec0d91c1", x"12da917a77d106a2", x"7634404a8581d217", x"9452fc35fee6352f", x"2fa20bab63ee92dd");
            when 4619753 => data <= (x"a7d02446e6218913", x"9be9d9f08b7d2ac8", x"54f3b50c1ef7ddd5", x"b0849a21a2e0efdc", x"10f53121599f2f3b", x"930622aa1101f0ae", x"5be109f40756ca89", x"35583076fa2dac9b");
            when 22686438 => data <= (x"5b5d02bd03d0c2e3", x"66882ffcd411b5bc", x"7f368620d5e9fc5d", x"ab40a47606e3bcb7", x"f88062ac7ee3ad0b", x"2bfc36c00bb38d2c", x"2d0f7c93d7109798", x"acef6de03fa69cd0");
            when 33791849 => data <= (x"637412b91491dd2e", x"fcc652293562f358", x"e678559028074253", x"c807f00ee3c6fed8", x"232a45291e07468e", x"498b9eed1bd9fc37", x"d433ebb9cc745d90", x"3ecd97403130552f");
            when 13896521 => data <= (x"0540e51786ae05ea", x"565f74b0e1e1b212", x"eaba1a997dd10945", x"5e6e9ee3e27f25a1", x"c5f7418c922c06d5", x"4e517e00218b9af0", x"0cd2da4116e107c9", x"9480f04df274b750");
            when 23793395 => data <= (x"969314bc31b23ac2", x"6ce8472efc3271c4", x"673bcdc768e47a38", x"3ac5222c410ad261", x"b8e3f975717687e6", x"e569f16b522a102e", x"b36531d25786daeb", x"eadc83ddf6b4bf33");
            when 22707860 => data <= (x"92de227a8fdd5236", x"f7839cca75dd1c2e", x"1d19502b9751dde0", x"a9858cf94924ff65", x"0be8d30f987e6980", x"b71e8e12b0820a18", x"de35d8df9ec4ca9a", x"fa0b53df0eba8a1c");
            when 19078400 => data <= (x"80fb5893ef19cbfb", x"0806863595be2028", x"189b3cc4d34ca2e5", x"1254298961c75a15", x"72907c28890e019d", x"c057376cd95a8364", x"0def6bd02419fb5f", x"f4a33685d0282f6f");
            when 28773423 => data <= (x"fefc6e1e3799d7d1", x"7ebf8232fe1420c6", x"15469894c3a3836c", x"e55b7f4972b02545", x"9a82f280802908b7", x"6eddc30c12d5d27b", x"77a7c9e257012bf4", x"79a65b12a865aaec");
            when 8151477 => data <= (x"7708bc352079c217", x"e37ebe51da9b5f9b", x"d7764a6d2cdff01a", x"8082a377523ece7d", x"3039827bcf417d3c", x"c27ea2b9ae3a664b", x"a1f98647a063afa5", x"3a43d74140ad7319");
            when 22268487 => data <= (x"a33f5e1a4194ecf7", x"6a12e6bb1eab01a9", x"636ede554a16eb1f", x"b0949736003ff47e", x"9b20c91c4fea9d1e", x"6f1707dbb42b5058", x"83756e9918aeda5c", x"2998fc7f996a8674");
            when 25878461 => data <= (x"283f0f6a19f87749", x"384bda16d9ddba44", x"ee77595f2576b014", x"0fd5ac1a20dd1672", x"15d152a23478b95d", x"0db980477d8fedad", x"8f5b60082cb7b403", x"a41b8388d5993d4a");
            when 7747015 => data <= (x"51a7723adb04d2f1", x"a656ab6b3a024861", x"386924901f1cffad", x"e0cd47c7016bb3c1", x"06144a04a0f35a8e", x"351c3695c4e1dae0", x"a20a69767d4e4d4c", x"2a673ba9de99b00c");
            when 25361786 => data <= (x"a8857f3c32bbf64e", x"501a084e87e7a0f6", x"825b20cd7a41dd29", x"8ba2815a3beb7cbd", x"6b8fc813152e6e31", x"707e458c337440cc", x"102288bd58799141", x"0f785f5bf503d0d2");
            when 17091388 => data <= (x"d1f52056e7710148", x"b435c570d2a109b0", x"900f5d1bee1f9100", x"f41567827446e7b5", x"dbdb7bcee73247c7", x"1e997fb7c2832a05", x"e1fc179edb39e912", x"10e59af12b6af64f");
            when 24055053 => data <= (x"da59d5966684d756", x"a569c43cffb3244c", x"a51f88e551d2ea7d", x"b5f76dde7362a117", x"bcaddee8778a9d57", x"78942bdfda2c4343", x"9be6614a87260f40", x"50b90ef27f695640");
            when 7177128 => data <= (x"6cb92ab8c5eaf54d", x"b483a3a66f6dfb91", x"d06e64864653823c", x"6e3390fb85e73b7c", x"ba58a4afcc69dee0", x"e30c0dcabcb4afc0", x"0ccfe5f069bb83df", x"58f7d77620238751");
            when 17383223 => data <= (x"91ac908cc553fce7", x"7336e5badc4040b1", x"7a630fc7eefa541d", x"6623331d0dbb5d94", x"8734179f6878f42a", x"c206992f8fd1004f", x"46d71b0d8040fccf", x"b4276293209929b3");
            when 8785579 => data <= (x"009770059068636a", x"45e552a48ecbf622", x"03bd07c5d2003514", x"f702c3270f7bef2b", x"863c4cf308b8ec22", x"d7a25071ec0ff77e", x"83676240cf4c2772", x"108ae345b2f807de");
            when 4541816 => data <= (x"0777a88e2a82a0cc", x"7f48927132932982", x"5731116bb722892e", x"34abbcb095e93e20", x"e446d2a79c36c885", x"61b666601d93b959", x"6f64ab21f4d8d251", x"43333fec2851fbee");
            when 5475605 => data <= (x"343bd8b4112b4b80", x"6a99b406ffa098ac", x"d5e0c34a93e8d466", x"136c3ea348249425", x"bf704e7ae40365c9", x"e473b5517b7f7565", x"98bb22b7b178d1c5", x"8cc46183508c2bf5");
            when 15308281 => data <= (x"e06a69eecb0c770a", x"e0e2af8011a1cb76", x"5fc9aea3b9fed801", x"a5db7a59d72b002a", x"8504e2df6e6b66ab", x"a88f60977555a982", x"47363f763fd18489", x"df90b8b9ef528a89");
            when 11013142 => data <= (x"f8b5ee767e486d52", x"5bbac0697f44caa9", x"bbaabe99849a6973", x"8ed2a90e3475fe50", x"e303fb20e04befb2", x"5cbe90895f48283a", x"caa9364309f1ca79", x"5557bd8bfaa48e5b");
            when 32702697 => data <= (x"d09776fee9338245", x"8958154cf0bb7e3a", x"8113ee6bb72a39f7", x"d988390ddec99100", x"890e3762b16405fb", x"4ff726207dd12de2", x"79fc7cf20bea5827", x"6d32996b2eb5505b");
            when 6970384 => data <= (x"a72f3c0f26981727", x"c891f50c9b73b402", x"70e3f906ac111f94", x"7098521cd4b87560", x"4db0a8647ded0567", x"6cdc4f52defb7c4a", x"8b6f8aeddc5c2c79", x"ba9e51e8f8d80e1b");
            when 2528628 => data <= (x"7eb970f5686cf478", x"af477db3546dd7e9", x"bb56e2c3e8fc7c5a", x"2c3e29944a27b435", x"bc2a78cd4e56189f", x"b74a64c27f73a399", x"2c64bb7f48e88cb3", x"1bc3258b387e2377");
            when 16861048 => data <= (x"e2590e92660f7081", x"122a8f938060f0df", x"ea860bc0d764bd30", x"fee6e20c5e55a10b", x"733ac2fd2e4c6ed0", x"8489b5924e48a984", x"016e6f867f14d482", x"96cc5afc96fa9f9d");
            when 15694698 => data <= (x"ea28700a9eb130fc", x"6c4246730da0abf3", x"fa5815ee8d111957", x"39104e903db2f820", x"fea0d3aebe25a966", x"24498eed9fd6941b", x"ab1356e333c17f81", x"235414fe4d8bb765");
            when 28616048 => data <= (x"a721e6090dea4130", x"9c0259b369e482bd", x"8fe72f69121b062f", x"9213bf0cc0ad2296", x"7e154f201baf6fba", x"bfa806326970ceab", x"f7507c0907f17d9e", x"51753b05c262d62f");
            when 15501246 => data <= (x"561d5739119c307e", x"3194c5647c22f78b", x"2f9ebda5271af632", x"8e3d884bbe341a1d", x"09cc80795225371b", x"3c587ee01fd38a02", x"e13d0a888016b43b", x"d6a26992573ec5bf");
            when 1151327 => data <= (x"eb42093ce800361f", x"8523c10df5db6610", x"6f24a604597e609c", x"c34047ada6748a1b", x"2f58fa8c42ef96b8", x"5f1b35a9cb8fcef3", x"5d838b0aad2ea136", x"fcb36d0add87b549");
            when 16162173 => data <= (x"d37223668649d7cc", x"ec618a3e42686f2d", x"ea3a6762047e500b", x"0da5b84a63dcc57b", x"0a224b7dd3e4df7d", x"40db7dc82d9416a1", x"abfb3c5d1be45973", x"d4df71c05aaac184");
            when 24126861 => data <= (x"8ce2ab5716921605", x"eed5cb3f7df74436", x"d2c5d10b04132e9c", x"170d0e968d2c08a1", x"2276012250a98b65", x"f1c36326dca14bf9", x"99bd30d80fa140c5", x"acc02a61532999b9");
            when 31979573 => data <= (x"f1bc783cb62fc29f", x"524ebb6142330875", x"e9032dbdd149af55", x"1d85c4a28205ac5a", x"4426ba270bce91bf", x"6408a873bf93ca1a", x"c9086bdc1d89e0a7", x"fa991500a3ce4951");
            when 23984777 => data <= (x"11affb1f6a4d79ae", x"9ae84e3271451ed7", x"0390bccbf2b8ce90", x"00fae25cd77ed83b", x"e2e8d72f6c1f88c1", x"62986cb02a5dde8c", x"37f968c9d943cb4a", x"f36d1be0c82abf29");
            when 14062591 => data <= (x"ed3003b1abd28382", x"7d1257d0991a4e3d", x"0d960b1b2b363f1b", x"8a384e7345e62121", x"c36fb218c0f86311", x"696a3aad28e3e022", x"d582a3758b086bb3", x"8a89d7286a9d7a1c");
            when 14810146 => data <= (x"bfa489065ef1b7ed", x"9a49afc8800f5b65", x"170f0a5702b6d3c2", x"a6206493b611f25e", x"88fb49e08ff5baf4", x"b269416b40e21ac4", x"4b63a4add0284ba7", x"84f8e1b7bcf8d12b");
            when 33933096 => data <= (x"be180cb6df076113", x"02e4c1fda6f8c82b", x"1dbfa9c02e980133", x"cd4d1bf39f08bb2a", x"8225bba7bf2e8255", x"84c7b6d736b07bc8", x"bb2323b4b86ceb52", x"0300645191d134d3");
            when 26215489 => data <= (x"30aeefe2c67fa76c", x"cb8f3fa0ee6cb694", x"403b56a2c0c4e7ad", x"7fe974b059ed935e", x"ce35bbb262f2ecd9", x"314c3522b7fbd259", x"de7bbcaa9dbb9c53", x"b5e69b48068ad10d");
            when 20292328 => data <= (x"62522b5dbee341c8", x"36c4c041be932685", x"4d73904929cd8564", x"74b2c8944c818d2b", x"6f955fcc824b8e05", x"262560221235fdf6", x"224439e058c9ebac", x"7ae16052053a809a");
            when 15085713 => data <= (x"88d86ce3a7782afc", x"a36f237b003228ef", x"126ca38198616dbb", x"03d251dd8023447b", x"d5e9f65a5902d3e2", x"7370f3c607b4fb5a", x"d2cc0e5f1553e74a", x"e6f9375df9ca7fec");
            when 27284464 => data <= (x"779393aae0cda5d7", x"2a08b2473bf3aa0a", x"2be0f273171a8fd8", x"2bdea476421c2e42", x"637cb142c4b9a2ff", x"1ddfbb39a85dc208", x"78069d06fd41974c", x"d09bcb48046c5fab");
            when 29913292 => data <= (x"9aa446b806a3a216", x"ecc540999e40ed72", x"f113d098663a67d1", x"10467dbbd73dfafb", x"c061c8da460fe74d", x"bfdeeba833a0aba8", x"4c4fdca6565ade6b", x"b51167a5d9c8d2c1");
            when 8284977 => data <= (x"05a81c40f615d8ef", x"8780e65d94e9fb0e", x"d5e844f344cc485e", x"ddd1fad626affc64", x"8dccdd1b7884e1fa", x"8275ae9472e4a81a", x"0d745d57976f685e", x"877689e94440a0b8");
            when 27237399 => data <= (x"f23be2b248ae4d75", x"6ea3c13550c1aa3e", x"702c160229d94330", x"0efb545e88d1ce9e", x"40c812361ea5d1f8", x"a52e5474bef5b58a", x"9f5565e5bdea5aad", x"7f3b0cbd2d414f8e");
            when 528785 => data <= (x"a2db7fe2969ebf3a", x"b3b6286cb2641efb", x"8f9645e9cfb1e568", x"af6cbfd259f23e72", x"24fb7a775cadc696", x"55b151ec1ac8f862", x"0570d590f7ca2603", x"b145529bcb74f846");
            when 12236918 => data <= (x"e4f4f2d6722e45fe", x"9f387cdd977b25ee", x"51bce1d05d4b5afa", x"0ffe2723d1b73f6a", x"c3baeb4eef97af08", x"8489e2261bb5eb23", x"81e7e017e8488a70", x"cb8546968ff72b5d");
            when 26725321 => data <= (x"721779a0585c8509", x"54880af6a86a68c8", x"fb284334006d76e3", x"874befda7a356551", x"70135caf2e62ccf6", x"644a61f4d3fe3a8e", x"19d79970320931df", x"fe43d495a115e211");
            when 17389044 => data <= (x"85fd472c4da48235", x"e5fc92dde40a0020", x"b813eb6a957225f7", x"a6b0b76f9dc0dbc2", x"c9a8e75dbb7e73f9", x"7c9f47562db79479", x"58465abfba3bdf66", x"8044f396a395df8d");
            when 9008511 => data <= (x"78326860b1c00199", x"eda21c273fecde04", x"414e2c3b87bb1711", x"0d090989ee25c12f", x"ad518bec0239f6f8", x"38c6d6b8c510fda8", x"26e13f1f9f9e8724", x"a0f77e369b3dece2");
            when 12289228 => data <= (x"4ba73b2cf2c60ee8", x"c48856e10774bee9", x"a751192b97b8b839", x"12ac93f4c51183d3", x"0f20d2478bbc9200", x"aecb3432686b8712", x"308e21f38b5869d0", x"8d9ae46b5a0587eb");
            when 30346980 => data <= (x"6d051740b60ff913", x"34a409de012cf23d", x"6112f8a22e3cad9b", x"0bba409d694e08b3", x"bd0b7a2e92bc563d", x"148cc2853c871349", x"164f6cb7e26ade72", x"5b7aa8e3d6bd0b37");
            when 26603116 => data <= (x"eff6687da99d7ad6", x"c69e444772ce002b", x"967186100d49feb5", x"c52f08f0b05d6485", x"fbd36e3e95e83e81", x"e007becbaa362f51", x"80e26e8d143e715c", x"b8d544ad512778d8");
            when 8528332 => data <= (x"5403ba36329333c1", x"9ff392a68bddebdd", x"a6e4ac2fedfc9ff8", x"17bf784eec0b3bd6", x"76b00aed89bca891", x"268a4b89672438a0", x"314be4fccd00c191", x"d7baae2af9aeba54");
            when 11912385 => data <= (x"4bcb43f1b7c64a63", x"bb9b1679e167330b", x"f3c5cb5ee1b1a8c2", x"9bd39d1076d97c31", x"32812139febd3861", x"6d43b0a8d6336533", x"e66908ce69b32745", x"8e24bd4419745ce0");
            when 11946112 => data <= (x"6a7e3ef1c3657b8c", x"1dab6925aadbb71b", x"a33ab14b09d2fe41", x"6469d6f1e35b5058", x"87ec8bcc2e40c4fa", x"c72a4191b7cae6d8", x"3a00422a0335a0fc", x"7f98e1a7b341466a");
            when 24691646 => data <= (x"966556240ec7c219", x"701be70596c06592", x"6d570054282d10c1", x"af45f205bb572463", x"c43a41bb227901f1", x"6ce9d5b98574ca36", x"0c68a9ecb6d9c3b1", x"cb18d5bb3e2aa21c");
            when 21681029 => data <= (x"5dd51f1122c6a38d", x"ed4de4e28579ffc2", x"391b8405bc512b87", x"add2c68048d18e92", x"35287f29c75c138f", x"4cd32e2228aa14dd", x"5fbdb50220091a45", x"99084a06007d931c");
            when 18794449 => data <= (x"36548b0eb6ef9b9f", x"43a8f909c0d90bf7", x"915e4b2b1af3b2f5", x"b24ec32afd248138", x"ca2221432c477929", x"44fdacc37a5aafbc", x"f5134affda4b474a", x"bff9151f8c2308f6");
            when 23540611 => data <= (x"74b149c62fe96a02", x"48ccc28b7cee41b9", x"497ae371f4e278c6", x"65e1863f61ad2aba", x"f96cfb5dea4b0bb5", x"b916793e27fcd642", x"dc3da5f9108db149", x"afbbe4a4614c03b2");
            when 26178078 => data <= (x"b8fc6187ba5d8d90", x"b942350b099107e1", x"c10ca51bdbbb921b", x"6ad860c34310d91f", x"2669dc767f62c6a6", x"eec8f6b3980907f6", x"834a2e739aa2d909", x"fd3a90ccce9ca992");
            when 19133573 => data <= (x"f42b5b046794f724", x"13de7708e216b523", x"d75862cddcfe5487", x"4238709a7407d4cc", x"7727226d75bf833e", x"67767b02f3e3ab4f", x"6946b51823517b61", x"8162186e5d6a40d4");
            when 30835064 => data <= (x"6b9ab8d546da1bde", x"5d6e698a50dc421d", x"deec86b757b0e53c", x"961716506b76510a", x"503432cbf0b6b185", x"a27fc619b42c982d", x"3137fdc149b26118", x"cbf056efe3b96594");
            when 20560945 => data <= (x"c87dc67e9a2e825e", x"ad7627a42cf04690", x"10ab139b04b879a0", x"e6241dffa5ee1bd3", x"058b02c7af5bb61b", x"347d64fdf6aad86b", x"669bf392d51b35cb", x"90d61565019480d3");
            when 31082433 => data <= (x"73156023b3f12b81", x"daa8bba39893c07e", x"24aab6ca4619d89b", x"58d90dd3b19682c1", x"adcd3720eb14bc44", x"bdc08fd8d09155df", x"add27b56ef0d54e7", x"7396e518a4606fff");
            when 10337808 => data <= (x"bf742f7be1a08527", x"d585ead2a2261c8d", x"66b753d4d6e6527e", x"8d068d1cc72ec4fc", x"7c3f1a6f1c1e0611", x"495d5eecd21e951d", x"7110e6819c05715d", x"313f5528f14e9e6c");
            when 11672434 => data <= (x"24018f98526069cf", x"ffaa78de2f3acedf", x"f3dd70d03cc8a549", x"31d8e0821e2f9444", x"51b34c4092ca05f7", x"57f9fcd5805e9f77", x"d578668659154524", x"943dc14f1f831234");
            when 27932788 => data <= (x"231ca9e2994a299d", x"376a189fc7b770a0", x"b659a1473da64155", x"88fa7c2738cf0fdc", x"78f3ce23afdf9da1", x"b535c1b6afb4af44", x"6e4eb54e615d4eae", x"db91eff5a2d7a0d6");
            when 7553738 => data <= (x"3fa255ca0ec25970", x"bc9d9bd5d060a5be", x"3554f90c39a17ac9", x"6945cf92c23660de", x"f4cfd10239145197", x"5a67660b57460daf", x"9ffd5285c01d5f8b", x"6fa265185ab5f478");
            when 4819194 => data <= (x"7310ff4a4df20ec5", x"ea5ad0c1c9fd9b4b", x"04f02c1caaeada11", x"72b7f3500aba444f", x"783103677bde5fcb", x"9e0e55aafca0ce5d", x"c35014c4f9b8f6de", x"de42bc9aa787cd95");
            when 14124825 => data <= (x"2a7ad81bd2c714e2", x"f0fab0384c9afb84", x"e607aebcfc933cae", x"bb9ddd64a26482a1", x"142303ec85ecefee", x"012ec87ee3640661", x"2368cd8150a904a3", x"2aa3ddc35d44074b");
            when 3151750 => data <= (x"46cb2e4bac52aa08", x"c285400a3c2f9ad4", x"4ce3f1a505dce901", x"a9b4051e31372b4f", x"d81991ef6781d4fb", x"fd398c68dee6ef40", x"e4c44ae4600bbfd0", x"9cc37eab5427bb46");
            when 8133577 => data <= (x"085b9c2cad07abc9", x"f0a56898617c4f59", x"1c58042deb3f5e8b", x"cde1f7a2363322b2", x"2396f81f13e201bd", x"b9f34c1c43cce4bb", x"2cfbed2bddb1e3f9", x"2a566a6ca07f2ab1");
            when 20216843 => data <= (x"6a52fbb62acee6dd", x"712ff249b8ac4526", x"205d0148fb575f85", x"9731b26d8ebca800", x"a84b5ba69de1519d", x"a673ccdeea37dd90", x"23bebcb54e38dd93", x"752928f649b005c1");
            when 14390561 => data <= (x"1822eec197197a57", x"0802cc0c8018408e", x"4083c5f4b8976fac", x"ac4774b9812c5a50", x"bd3ab98a83951682", x"75cfeeacb178c32e", x"958f439f365945ea", x"e82d26b21d74cf44");
            when 2729003 => data <= (x"98e3f803eda16b09", x"71b4af5192772935", x"ff15fc0ed69729e6", x"5a8eed99ff637a0d", x"7d4d04ee04b77375", x"78bbaf6865e779ff", x"c4d0124a39bff7f5", x"8b481a8710e26bc3");
            when 14716066 => data <= (x"ef491b1dcf4861c2", x"09ebc46bdf3e22b8", x"4bc915ad7811641e", x"cded78302b58402c", x"79ef658a9a2e6a20", x"052318a4f9e7805f", x"65bad287fdb0bbc6", x"dba9e2cb21f5b079");
            when 3145942 => data <= (x"e6bb2fa9658cf422", x"f3947a763dd6f284", x"9ae6fb91dbda7497", x"2cef6e2bc146f517", x"0f919224d72227ff", x"2c4b331a36717811", x"fdb747dac089733a", x"121676f4d1f5dc14");
            when 1266214 => data <= (x"f30fa11d4a818dd6", x"c22dab42c45f4c0f", x"90dd1b56d130c465", x"8bebac94f505b00a", x"c204651b0df4344b", x"7188cc3d25837712", x"1bfb2439b36392c5", x"f5a652d21e81ef33");
            when 27453341 => data <= (x"c12e0db6e0fee9f2", x"1106d28122163a62", x"05db0f4f99cf9caf", x"33d49687891e7340", x"85b9b1a25dfc3831", x"70436ffb1adb17e8", x"621c41cd81f0a7bf", x"df7dd55d683577c6");
            when 15026717 => data <= (x"36bfd9cb9eed780b", x"19b2c6a537d87141", x"a2811afbf9698616", x"c20c387e88b1b290", x"cefc754c72bca414", x"7aabc0e0d47b5c4c", x"727ed2b95f5f6e0f", x"c6378919033f5285");
            when 1073861 => data <= (x"d2e181943bdb8aab", x"3f7964564d8bdef6", x"416e73db06e7388c", x"3a5cba00e4b5eb50", x"ba4371bd35b730d2", x"cd25fa04cb664637", x"ba18aa826f2e826e", x"351f50a43c0d3f86");
            when 28563748 => data <= (x"73f0a523c6a1bfbd", x"e59b41f2aeb7d3ca", x"1c5b1508a93a005f", x"f496b12969d5af89", x"5035b6685a62daa1", x"e0f790ee2ac3260b", x"b831879ee67cb858", x"1f479b63a378f1ed");
            when 19678038 => data <= (x"61a8d6551c2aa3bf", x"ed438e99a4f142c4", x"dfb0527ef9c622bf", x"c2538334982d31f3", x"803a3134a0f5e2a1", x"d8bb953217defa4f", x"87c888d1c4b1302a", x"07bd8a7b1712b092");
            when 10815172 => data <= (x"b274c7cd92744e52", x"3d000a16f0df263a", x"2ff36d92834134a8", x"8ed73cc93f83f0ec", x"4d710b64c652c6c6", x"0e7edf487cd5a1df", x"8ee33a8c6fde9d32", x"6995d8aff3305c59");
            when 776426 => data <= (x"f71b41b892e99757", x"a4d7ee0cf3213cac", x"f232ba7a0a9a8054", x"75b4ec9585994525", x"f51226840ba7a435", x"fbc97fe022f95180", x"8dcbd5482d8770c3", x"b36ef2db76db9151");
            when 6798664 => data <= (x"b58aa2e127a51050", x"f5e3a469c60a7a1a", x"3e8431b826981a37", x"035d19e3c68294d1", x"f16d39510d493ecc", x"418909cc51e7cfc4", x"cdb04f23d3c058be", x"72728f60a7bf62fd");
            when 2910703 => data <= (x"75bec310143431c1", x"dafc2d7710913b01", x"5e2383a97bead9af", x"9e348437f94fcdec", x"261c58d820af03af", x"3ba20ed552f11df5", x"3272581382fc895e", x"f77eee3a27896e92");
            when 28300733 => data <= (x"841a5fb859adc8aa", x"93e5c5e0d232d686", x"51f3611981701f4e", x"be49ebfaf04a2606", x"af0d094a61fe37f2", x"f1cf9147cc0d39e3", x"b7f3178b8d31a195", x"444b892b5407c44e");
            when 5175753 => data <= (x"bc3e13a02df009ce", x"1f0859a8e67ba66c", x"c421c04b9c99bcc3", x"edefb817cf67a83b", x"dd4448f8d0a92ef9", x"c5cbb8c62954d4e5", x"40e0b5890d6385ec", x"46a49cba97205271");
            when 12568115 => data <= (x"889284a3d9a0bd80", x"5f9016810adc58c6", x"4506e9fb045f0552", x"2b312e8a1224701f", x"a3b2ba971054f5b2", x"1421d2761b52f140", x"1a21909d7df00e87", x"83b3943a04ca8999");
            when 22839408 => data <= (x"465e1f04038fa730", x"52ffd3a8c49b29cc", x"eac3821350885c8b", x"6c8c2141245f8a8a", x"285dafef8df8459f", x"ffd927931d877b1d", x"24a87fc82921636c", x"41a3d7f595a52b02");
            when 32321942 => data <= (x"6d6c339b76d1a67c", x"56e35b685da9504b", x"07e9381e4b361923", x"5fb459a228bfe3bf", x"7f2b51ad71c30f03", x"5851408884044d6d", x"8297b3a78d08b913", x"dc6112f22249614d");
            when 13611191 => data <= (x"c926655a88463cfe", x"af8dc23dc0f690a6", x"e978045a8d02db47", x"52044ce3534e832a", x"1db7adf4485a3ba7", x"5a5729f4998949ed", x"b46652fa13c66e91", x"0e3b1ad1ca39401d");
            when 17008598 => data <= (x"baa2bacb1cb71db3", x"0231da76278dcfa5", x"263a310d7f4b0082", x"84a2d3d62f60150e", x"a87144de43518865", x"f43ff5eb41c21a20", x"8d3160f6e10cfef3", x"7a1d3b03f9dfd2cf");
            when 31955198 => data <= (x"ef427eb03f1a0819", x"08a250c087047881", x"9cd509224c8c7b8a", x"349473cb9fd6e6bb", x"d740c99cc0f3e5a7", x"f5394301f5dda5b0", x"1173c2454e3b924e", x"f209a99f36f76e2e");
            when 19591541 => data <= (x"c8a8bddaed6791e4", x"cce887a99bb51201", x"2d50a14445152ed4", x"4c32247b8b472432", x"0a0f0739abce226a", x"943789041d896492", x"5be20acd6cb04565", x"1007dbc12691176d");
            when 9556956 => data <= (x"914e006401cd08de", x"b4416d3bce73515a", x"713471aaf6ca1734", x"abd9a7bb3dabdece", x"107154caed5c67d9", x"6c83827bfc3e5a55", x"4207721ad0e0f85f", x"08b5b54b111412ce");
            when 22599330 => data <= (x"28022c74c17e44b7", x"cc29c74ad93521e8", x"3ac036b03dbac84b", x"8de7817dd2919f30", x"0febea5890795079", x"8aebcb0608ee9f31", x"ca41b2a7e057449c", x"71a5db60d4bfbdf6");
            when 16063017 => data <= (x"7578eb9c80c96cac", x"1d84423c20f0a759", x"c6376086094fdf49", x"f4323a10970d8abc", x"7bbccf8c7c3f5f5c", x"eb859481b0e64b73", x"b34a1f36ab7f6a9b", x"4627a47346dab038");
            when 11042727 => data <= (x"2ffc00d74c9c5222", x"442eed89379618cb", x"169547f95c4a94cd", x"23ac56b750a67f5a", x"3194120ed892bd96", x"5b56ba1b15cf91f4", x"833371a6a21efbab", x"1707291feae23e25");
            when 931061 => data <= (x"a56febd3a5098605", x"d3498cfdf0516b03", x"c9c32340821af48c", x"8b70b6c76c16cda3", x"9430146c9966bbde", x"7bf3a3d61c072dc8", x"5277e618db44d819", x"8734f997db517111");
            when 21988696 => data <= (x"4facf1e1017d9889", x"8156f99a306f173b", x"83bef24b1b6cbb6a", x"1c7b8ba52b6fd0f5", x"4a4896afc812da53", x"220c1fbc5a78f9bd", x"44a2fc97fae5f90d", x"16e1ed5fa8dd5e2f");
            when 27093158 => data <= (x"80e0eb030beb62f7", x"9590b28ca4c41c60", x"ff96444bbe8b09a1", x"a4913de33ebd6cf2", x"2c6bf45fb1ebaf71", x"71ac294c05b51cff", x"318a50442a88480d", x"dc100e7e7ffa651a");
            when 21823149 => data <= (x"fd0186fcd0711723", x"9d4a47f6c22c7ab0", x"1c2f0c959aac5614", x"69a03722e9cc38ec", x"3a4e66efbe3672ff", x"cbc4a1da6ca1c4f9", x"6b150a2d6f13a17f", x"db1a1be5d6e5736f");
            when 17712343 => data <= (x"aa3cb52e7b75ae40", x"3782cb7731076754", x"dc46ff58a7326a24", x"c5ea5033f943a75e", x"5b25801f95377d99", x"b9ff1dbff567b1f7", x"879005c0fb50f7da", x"b3131224e22f2898");
            when 26051535 => data <= (x"1a40b98f968e58d5", x"fa89870f5eba4431", x"658133d0c1480c24", x"888653b1f0f8e40a", x"a3212d060cbbe955", x"6da3e658e5f09e8c", x"f9eb61e3b04d523d", x"f9e8ada9595c4078");
            when 15789679 => data <= (x"73c73947f0e22742", x"6d446a8919d09239", x"513c25285425a100", x"944f6b4d849614dc", x"5c70c266183c0724", x"b129bb39ba0f78c5", x"a9469b03d9089512", x"8d3e6ff4a1a8777f");
            when 28320462 => data <= (x"f49fe295236a37b9", x"0465e5d1c891b14d", x"0ae3bc097af3f9ef", x"19c3ae1fda112361", x"10d41279711f7201", x"edbfa347e14f6ee3", x"48d9ef49c72daf93", x"d9fb5d9f5f3fff0e");
            when 4798444 => data <= (x"90e070f9ef4974c4", x"1902cb572797f5af", x"0863b342945a7759", x"445dc9ac41b8a198", x"7c2469d1256d7790", x"c7148a9c4a499f0e", x"d628ac33b7fdfc12", x"50115259f17f978e");
            when 22732166 => data <= (x"fadc80053485d5b6", x"59d035eb0bed8485", x"d152cb2e1c2e3fd4", x"f4ad17e601f70452", x"bc1cbce840934b60", x"9ba56d36567fddbb", x"9dbeb25cce0dae4e", x"084f553ba6c80d83");
            when 12325674 => data <= (x"3e991b12bc5de9d1", x"905925c6168d7a3f", x"f1bc84985a6d3570", x"4a8f3f1b268712b9", x"4cc2c0e979bb03f3", x"78a9937e80fe85b7", x"76458fe7002a7009", x"d0f8ae4b3d426dcb");
            when 14510741 => data <= (x"f66a4d1e83942c06", x"29d27ce74741f0a4", x"d5066d94e2fcd872", x"7474d03c92e474e5", x"81b93a32c8e0d984", x"829d381bd8b08d27", x"d1a8f5824235e985", x"17f7fee40a3c830a");
            when 3003095 => data <= (x"dd3c594627a6b84a", x"ab6820726c36a79f", x"d59b26ea0404a907", x"db0f5216b6fbf0e7", x"4d920b5097c3e1d9", x"af7721fb21610036", x"eb11fd3e591e6fa6", x"f6a6ac863c77cd45");
            when 29490490 => data <= (x"5d13740df79ba81b", x"b69e0228781f0783", x"65178e3ad9de35c9", x"91b8c97bf34e5fe9", x"2e0e677c001eda41", x"e3ceee06091c75d2", x"f8c423810a31cc38", x"af6a0e449d1ec388");
            when 23219090 => data <= (x"c99e159c66d47727", x"fc4009c4ee43d4ae", x"1741c4730737a242", x"25a5b387910b8597", x"e4c850b6928851d9", x"4aeab295f02e45b7", x"e5d5d7b6cb19b662", x"a9600c0f3492e5ea");
            when 10696833 => data <= (x"a9e5c7c201f74795", x"ac0a6d6c448a72cc", x"960275971439b6e4", x"4bbe657cce6bc7a2", x"24698844cc3967b8", x"8098701d811d86f2", x"8e77ac00895861cd", x"ebf3d71cc9318786");
            when 19994169 => data <= (x"a36339d4f0931f4f", x"83273c8dbee18d08", x"bf5d943e9ae6830f", x"01284a80c29532c1", x"b4649f741f6f8722", x"006be54c50723551", x"f67383d1f83a5c60", x"59c2f33f7420f3cd");
            when 6505204 => data <= (x"26a58ccf4da8c235", x"33f7c59f786bcb98", x"415b327adf7052e1", x"a9744fd265c06673", x"16da8b0011106b8f", x"c37051d00aa665ca", x"a5dabd78ae4ca246", x"c6a4244142150916");
            when 18252488 => data <= (x"73bca212780adc26", x"5a748cee478234c1", x"36d1069aa50c6f7a", x"0af56f8000333aeb", x"e21c59c0db11d2c6", x"0bba4b31e28d79a1", x"20bfd81c80f9cf42", x"b9b0666f76e17faf");
            when 24789056 => data <= (x"0bdac45f98ee76c4", x"1316c41355859c69", x"fc41b1a4a345b1f7", x"412483ecf9145f45", x"cbe53cad4eeed918", x"a874a5f441277f19", x"f21630b8f330555f", x"cdeba4874133b1b2");
            when 3652150 => data <= (x"4e575b399a69adcf", x"c20d3c2029440522", x"9bd0d610a4730e7f", x"a77a26d5552b88c3", x"cc0943ca5f21c8d3", x"e42e80b691022527", x"7f523e3bdd2b18f2", x"0cb84b43dec4631c");
            when 13872846 => data <= (x"46bca12703e9eea9", x"de672a32aa810f63", x"676e3089825d75be", x"278d37bf4b7ae08f", x"3a0e42069dc4e5dd", x"1e187e087c4ccd10", x"bd65b1fe445182a6", x"9c81a921580b098e");
            when 8645090 => data <= (x"0a1eefd83e53e5b9", x"6c54b42d3909180a", x"cef49d270195ac0f", x"cc6a7e8907bac28d", x"776b66b882632905", x"cbdb812f9f566dfc", x"f77f62a34bf246e6", x"19e3dd54f5e59ed6");
            when 23151630 => data <= (x"2d56e6ea15815a96", x"326ecee47df398b5", x"8099f21b8cecc9c3", x"9abb46ab7dbd61ba", x"ca9df800e99a2e67", x"10e5aaf24c39ea22", x"6517d18ea4f69f52", x"ed94e75926340a24");
            when 33212433 => data <= (x"7246adec36f7230b", x"6eb025642982b459", x"1fdeef1e00220b28", x"15b809322497b044", x"5129832f65a259e0", x"3ebd1f9dae852653", x"ec8649a96f2b9d9f", x"e0defca6d1ca0ff7");
            when 28780919 => data <= (x"87464adef515634e", x"333743375816c300", x"afb56eda6a069fb2", x"bc2a396446463960", x"1fbda1a299ad1295", x"aea4a290b60bba3f", x"273eec19f14c7107", x"2f20e8cb53ea5202");
            when 19652710 => data <= (x"f64f9d1344db9ea3", x"b0307bb28899ee01", x"c6e93d9a587cd80d", x"2e7f46eade5e5c1c", x"8bcf4bd3402280a9", x"0e6b33a57e3738f3", x"5cf1831b1216b580", x"9048903a6b3b2a2b");
            when 10740461 => data <= (x"78473a696c69941e", x"3a11534b4ffc2e1c", x"21b8acff39f08ea6", x"b403079fb4c8802d", x"6881ead652d2c22b", x"5bf217d29f64da2c", x"9afeabaae1fd2fdf", x"ead4eb1814d8c8f7");
            when 19233303 => data <= (x"f39191e560deade8", x"3b204d7dfa73a561", x"c66e18d2bd90d416", x"57baaba3e4abb2ca", x"3fc2fb416ac867f5", x"6fc160acbecd8659", x"29d9972126eab751", x"3d2e3a5221586de5");
            when 5507134 => data <= (x"6424c899638dfc8b", x"bb368c5ef1b542f2", x"ce4829680370dc76", x"a2628a0007020f76", x"1e1e1c9adeda6a15", x"a9d7858c461f1f2f", x"f75ea71919fb1e3e", x"cc19bdf99dc05d8d");
            when 18578096 => data <= (x"3be7f827509e0d7d", x"f306b27440e86688", x"d8d1ef18d403b5dc", x"d9e2dec7a2aab9cb", x"4ff5ee5a71c9fd5b", x"3d89e97fe855c737", x"473ed784896d8604", x"8ace16c4cabffb33");
            when 21428504 => data <= (x"9bbbdc6356aec8b0", x"4c9ef9d8627fb99f", x"4850a76516da70d3", x"07a61db7a085b62e", x"7cfe892a26aa6ab6", x"4e2301f0612c3b8e", x"ab429e317c593fa9", x"728fa6e3b5e11f1e");
            when 22467460 => data <= (x"0d956d768cdd5c45", x"9145b01056b7b55e", x"9a2fcc4731305030", x"20940801a45aa5ce", x"4bc1d89ea3516782", x"87ae1c11e9dfd262", x"54c31dc84ea53e08", x"8d6e4f8d83ea3a86");
            when 31763143 => data <= (x"6504323f6b466399", x"3927173f9dfc3a76", x"3dcfdc39b927700b", x"a99955effaf5ca30", x"ce18796b060efb45", x"cfe3f304b5b99b96", x"2a8182c81e5bd055", x"f1ad07f901b18618");
            when 33465809 => data <= (x"1dad32e7bf49561a", x"52a80ef7df4b3e55", x"c4e901a5d1ba9e33", x"0abaa0dbcaf3c942", x"968a376eb05f8786", x"8ee661a4fe86216b", x"21d91bfdb9a4709e", x"48644658efde3271");
            when 12090256 => data <= (x"c3a59288f88adf66", x"3efaf60ea017f05a", x"de635d4b1d4b7e80", x"7970685b32d76217", x"bb8005b3136ca30e", x"10b47b06ab9b14dd", x"9e422f40043fb7b9", x"a715e0199c0e1300");
            when 11381151 => data <= (x"426f61c69cca5406", x"d7b62766f59879bb", x"cd7423f9188740cf", x"56f2f4e986193bf1", x"baf7200b34650fc7", x"23390bba1a192d09", x"fadbd914234940a2", x"a43f6cb02cbdf069");
            when 6278771 => data <= (x"66fe0a2bd0aee814", x"bd1ca0b4d5724d63", x"b2817c0b48350808", x"8ce2689da1dcbd5e", x"1225fefd41e14eef", x"ed6ea77e7cf51928", x"fc6a8ae6365309d2", x"b23a7a75c3a9b656");
            when 5217049 => data <= (x"790a89f98a0672fd", x"ab03d0ad947a087a", x"b9d7aefd98f553ee", x"cd34d902aa4ee684", x"44e141afc85785bc", x"d49047a5218fc83c", x"5e6bd7d18f66d61a", x"c591ac2e04b819c0");
            when 8706815 => data <= (x"1a35b719388bcd61", x"19773780564973ab", x"3245796edb42ffd6", x"d67677e6a3e65343", x"90760e6aabe2df9b", x"6f21af1ebdf7ce70", x"2171bc205dccd12e", x"5a4ba589ae6bf449");
            when 33809055 => data <= (x"e09ad0451d2bd7b4", x"e2144c6a33351f74", x"96cb89fe56d5327a", x"d1c26b0dae40d244", x"efae28d1d26b13c8", x"640b1111bcbb0feb", x"e65f13e2a541c122", x"2a67165408037844");
            when 7523011 => data <= (x"9738a3cedac77e58", x"4e89a22e994f93df", x"66fdf5b72d809307", x"e8b854d6ce7dd8c9", x"4f10aded2b240523", x"20c6c74f545700d3", x"e46b24fe97d8e75a", x"7a36da749d7b1a0c");
            when 18634521 => data <= (x"7c59d55f116513a0", x"15aee5c413f06eae", x"7f9f058413ddd0a2", x"2d490c86494364cb", x"7994d685480c785d", x"117f21313e259c64", x"e4fa07f3f828a039", x"af9a3d169fbf990f");
            when 28077193 => data <= (x"1b6bf2dfe3a5dd90", x"f5d69832de858179", x"9aca05d437d75441", x"25a481e06f557912", x"f545dc0a09ef775f", x"b8f171310ccea2dc", x"2d0ce5589b81852d", x"cb211eea4418a048");
            when 25680552 => data <= (x"ddf47b9d323d4bb1", x"bbe62b50a03e29e0", x"2d76215a3475b4a9", x"8ead291ac58661c3", x"bcda6cdd9cdb63a4", x"c5d9e6f132c392c2", x"4c8c2a72ca80456d", x"9aa002184c321002");
            when 24481152 => data <= (x"84a59bdd84c33e0b", x"0fea33ffd91d9fa8", x"552d9b2d532373bd", x"5756c1abeed710f7", x"a790b5df4c4e8174", x"8d5ffd1d92a53167", x"4b2ce089dcee260c", x"6b6dbb734faa49d8");
            when 29897748 => data <= (x"ea4e38a80b91f9ba", x"89eec9cca2d24efc", x"4a5fc8c10ece03da", x"f93ced1dce4ebaf0", x"6cf8d73ed99d1f0b", x"b84d19d4d3114db4", x"2063efff9429bced", x"ec69824755619da1");
            when 17578068 => data <= (x"36817cabf427bc92", x"bc663d38a7cfafe1", x"d3d0a3b9916e662e", x"ea1a3209b4683265", x"b2b077ecf48688fb", x"954539e2e049066c", x"2e14d6d6960d9df8", x"418635dd3dfc33f7");
            when 19310373 => data <= (x"da107cb933b4656a", x"d188247783a4a51c", x"f16de65724eae8b6", x"5719e2cb8c7466f4", x"ecc6cf6d65d14f91", x"e88e8e4994205ae1", x"314a9b4c0909d475", x"c536d22847b07363");
            when 22645961 => data <= (x"e27bd2167670a7ba", x"4966122d3acf2a0e", x"a2fb1d8fb6d9177f", x"77fcc823589051be", x"998b75aa3bb37559", x"7a28f48bf7f46034", x"c161a1ee150f2056", x"5df8a51c4419175d");
            when 24026838 => data <= (x"0cca940fc865bc0d", x"f1a318b71e8ddc1d", x"acd7870df6e58d5e", x"923fb45df95d7382", x"9b54f886c4ebc223", x"dfd71b08791cae02", x"32ed18232e376275", x"6085cdf62d9a7825");
            when 12120043 => data <= (x"019c917e9f1fa656", x"353d47cbe9c2f382", x"08a9ef220a255d62", x"706c8abc27f9f1a3", x"f11d415f5623eea5", x"d3a70ef52ae87a95", x"945b8f7541a15965", x"3d52696b61a9d3f9");
            when 16278342 => data <= (x"b38e2123f81f647a", x"76a196c1015375d3", x"674d570692312a7d", x"6be0180a3b3b9a6d", x"8252317999fcff41", x"016d181bfc08e304", x"ebfe6d13e938741f", x"265c1bc597a5acbd");
            when 7261426 => data <= (x"5a43680c65fc4fb9", x"1f9c62b90df55da1", x"0a6836ca579faafd", x"fdb77a2ed8022d99", x"8f2676670de1266f", x"119b30ca6f29fc43", x"a661b4c38974a8ed", x"d7d77c1a8c637c17");
            when 25555589 => data <= (x"fa8be4d1e4c4885f", x"17b9f3b4843add18", x"9e8da2d7588cb231", x"c1c4040acc0d2653", x"b49596f1c41e560d", x"c77a86eab1df45e8", x"c8b0376de3c410a9", x"72f2d4fb04a8cd0f");
            when 4316241 => data <= (x"0f3ffc5fea848ec8", x"b3c21d38d8f9053c", x"548c7c9ddeb20fdc", x"05cb63cd5b7bd078", x"6f2aee7f77feca3a", x"e208e274d5db7e51", x"c5a651578dac3213", x"e8f098f70f78f5cb");
            when 31759721 => data <= (x"db292850e85c8abf", x"90de2c3c0f7b7aa9", x"32e181d700e891a8", x"98ddabe4cfa977ff", x"9cfc6a7b3fa991ed", x"47bece941d709f64", x"08cf303392e3c467", x"de49ce8cd244cd55");
            when 30769989 => data <= (x"300cc185b9ec50e1", x"ca36ca482be3666b", x"cf08c22cc2a0beea", x"099b7aaaa39340e5", x"3eccb93b19e5fab3", x"9dd32dc3075ee111", x"19586d7f5d0fbf82", x"434c079894fd66dc");
            when 18239320 => data <= (x"5a46df2e81120fa0", x"e8380fc70e6c3b7d", x"bc154a35d7b235a8", x"c01194bc8493414c", x"e8b3aeb31a240af0", x"3a25d20dfe001c3a", x"d023c39350dfd39e", x"d4e57de2d09aad9e");
            when 21745914 => data <= (x"b647e5615b8982ee", x"3145c9a44ab495c5", x"582c7d833703f393", x"28917706d3431046", x"265c6beb818576e4", x"3d66fe54b38ca863", x"2f27d80593be1a74", x"d62327426fc68327");
            when 24366349 => data <= (x"2e6d69b430ddfefe", x"a99696f869be35ac", x"0f6e35d1232035a4", x"8a764c612e3abd64", x"e099ceff2dc24646", x"927e46c57b12b11a", x"bb3c1e2cb6f89563", x"3d01405b3647b04f");
            when 17551928 => data <= (x"7fa3e3285a909135", x"008e98fb15afd6e1", x"267798d458c3763a", x"07fd34f41035ae3e", x"af1d582a8f57d213", x"98fb3ca85d256322", x"fc5466eb46963134", x"7e90d135a3f60a57");
            when 22288230 => data <= (x"36ca797a3517e5fe", x"54dc58ac84baaabc", x"883446d0ef3c0554", x"6f4a7677b2ff5b68", x"671d31360dae6561", x"5bea4947320a1dc8", x"0dd3476b983216df", x"5ffbfe5b1da8fa83");
            when 14337387 => data <= (x"247b4d494a1b6dfe", x"56eb3ed0116f7f4f", x"8da2f8731eddf8dd", x"caa886721d68c1ec", x"bebd0b6b9fe33620", x"8f949868d7ed78ed", x"f5c486bc3a70ea1c", x"6053466a3da59000");
            when 2221771 => data <= (x"45b334f002a09305", x"63cdd2f2f8271a08", x"dc7fcc15e1538f1c", x"b976ede08f3c103f", x"23095971fb84cb4a", x"321fb29d158029fd", x"22b665d36861ccc8", x"a1ccae775feea3d0");
            when 1925476 => data <= (x"d63d5314f4e75ad5", x"f2c655745924b8a0", x"1b8e6b4822b85402", x"4656e0a47366f0ef", x"8c82edbac20f03f5", x"50b19b8a2f5c28f3", x"9c663a4068b895e6", x"bbd3fdf47a45791e");
            when 24690910 => data <= (x"6439eb08fe1359fc", x"e326bcd6646379e2", x"4fbe6fd133f5784f", x"b2d8d6e59cfd0835", x"0f0cbaf4b9d9f518", x"0694dce66c928cb2", x"ce01ced0a423d7c9", x"2dda1e1cb61bb4b7");
            when 4107760 => data <= (x"a1b0595a952b5e0e", x"85dc81a39c2b74c4", x"ce3034f223747254", x"4296d2723ab1d5b1", x"076e6fc00de1d373", x"258702228e66b8a2", x"ebf9778bd60a22f0", x"94c485078a0c7c23");
            when 8947610 => data <= (x"28749998d61841e0", x"0c8d0e36a9e57626", x"9789c47911eb1573", x"96be2c9293061be2", x"b969af9e58827d78", x"8fc80dce4675dab9", x"c2eb58d3acc945b7", x"da22f055220bdaac");
            when 16000020 => data <= (x"c10a8f4c300af174", x"ebccc8067e20486a", x"cd3f8161d5232618", x"b257787dd1d8b716", x"29ad98c1eca72f9e", x"c658e0befae007a6", x"878913d3042dcb7a", x"7c88b87488aa0c07");
            when 20280145 => data <= (x"5143d59b3daacac1", x"eac3eb5d1df4fdd5", x"04f238007f80eae1", x"f7f2b7734a9ff379", x"ca17ffa6ef8b8ddc", x"2af4f0eb92008aa3", x"2aee1cf80859118a", x"5a6d4036b2cddd56");
            when 33779803 => data <= (x"29c6bcf504179710", x"a2e402b9c1490269", x"b158d0f412cdb287", x"4b643f811f1004de", x"ea18d9f57d9414d6", x"0d74cb3d1d029d85", x"1c6e3ec7e25f199d", x"b0d80d4ecb695c2f");
            when 19065624 => data <= (x"642133c4dc6dc244", x"fe9b17d04b8f4549", x"e98292b1e7d554d9", x"561d8c8df75821ae", x"dd56ff29125763c9", x"57faad2e539a9647", x"369de8339c56d7fd", x"c1e780d35dfcb390");
            when 22796875 => data <= (x"e2455e83a43fa294", x"c55a42945b018cc5", x"02864caff3e31382", x"554cccd445442417", x"6ae1114b54f13af5", x"85a8ac8a401857fa", x"22696ae94eb019c2", x"89c8b74db1d68e08");
            when 18083243 => data <= (x"e96765ef8099fe90", x"0a92ec5a691a1009", x"848b34c60cc3a146", x"c209b45dbe95b858", x"e49bb60373f73fae", x"4b3d7b4eaa97a536", x"f4c12f59ba63164d", x"4a767d43d14d2685");
            when 1604214 => data <= (x"5ed7dbf43b32a35c", x"1b03f400f168718d", x"90dd7d2dd6c4c009", x"0c0e4a5fc36f8b94", x"f64866b1c37b73a7", x"b065a5b909295406", x"d53d495cc9465e6d", x"5997441c9345064d");
            when 6642793 => data <= (x"1e983094603d30ce", x"b99b6a525fb9356b", x"cd7f6852f7ec91b3", x"bf8065d51c4e97bd", x"e363e525a76104cd", x"7e1e9e1900c15f98", x"2640017dd2f6c764", x"3c29adf412113cd5");
            when 20012644 => data <= (x"db33f1e24b253ec0", x"43965e246389d40c", x"d70a8db3011f7a29", x"d75c1006acd22d28", x"1ab99b6ae13c2ec3", x"e653ad12fefbf0e3", x"ea7cb9f5915d7e2b", x"b823b300c656a459");
            when 12192345 => data <= (x"7b9a142566073d76", x"bc483bdbfccca684", x"af86b3b5b1264664", x"1d09d7a09997fb0f", x"2b88db13ccdec4c1", x"755bd169762ba575", x"ab693db7752cb625", x"f94dd0f2f2687696");
            when 32316803 => data <= (x"d010f3dead3cea25", x"5c5ed8219e8d3a9a", x"544cda044203a165", x"dea0a17d1c94ef15", x"cb985278231f0f2a", x"b79ff242ba86c8ee", x"81169084b5c6b649", x"438a1a439103f4e7");
            when 17889926 => data <= (x"50694b5270f322af", x"d9e6a07dc0dc5a7b", x"3b8be2de48c8b2b6", x"9bafb03327e2d771", x"ea84217bee1c8b39", x"330d090a646ff1b5", x"eed27b836c30313a", x"462702e7cc767b0c");
            when 941209 => data <= (x"77714a0850cdb6dc", x"b59ae21cbe087f88", x"07c13531603b2018", x"c155844cbb688df3", x"2b52f2326cd840e1", x"9f050855de757c04", x"f467ac19602f591a", x"24c505587d53c8e8");
            when 19558317 => data <= (x"87c86477a7e29354", x"10aab6d2414b6799", x"96911e97044c704e", x"5dd8b28cdff070ec", x"3c53e78d5659348f", x"beff80fd285c7f0e", x"351652bdb251ef8f", x"9d0cbc12780bd877");
            when 14102222 => data <= (x"b26a88d06f2288fc", x"7e8032d350704f3e", x"2ddfae596c444a2c", x"05387d44462c2070", x"ab446d695c8997ad", x"d844282dba762c7e", x"5c3c8603bbcfd768", x"964124d14c8e7566");
            when 11239042 => data <= (x"1076c3fb16105dee", x"230dc8dffdd63672", x"6bbf35a140154b51", x"6d9dd5d0e11efec4", x"02a5fd2fbe47eb53", x"4712e4d3aacdb67d", x"975d09bcc1fb6077", x"4a9453d4a638d84d");
            when 24169335 => data <= (x"7876f77f3c029a19", x"5b30b64f75194623", x"5a7105b387a8dc2e", x"8eb218f3d3697419", x"874ae83e3f1f03a9", x"805f3ae9ba5681d8", x"67c23122d6674198", x"eba90bbcb26360c8");
            when 28118375 => data <= (x"68fd2a2d92beca9b", x"847364eb5668e3a6", x"8a8aecf233736fbf", x"8dfb96b9127b4f4f", x"ef74b7003593ce45", x"c2cf02afe691854a", x"47dc2dd3befff983", x"358b1a289893c49c");
            when 14260411 => data <= (x"87b07621294738ca", x"76bf925d10d6576f", x"79019a2000617448", x"8815af224e645fc8", x"2658f3896d837328", x"5ff83160e2ad083b", x"89cf53dccab805c1", x"7bd5d0672ca08d8b");
            when 33023547 => data <= (x"6daea222d93aa05d", x"fb3859513cc4b245", x"4091c74b617f3dad", x"fb228664d058c5fe", x"8020f9f501ce5a9b", x"1c72a3cbacb98091", x"fee00e85c25e2981", x"3de8cc74b0d7b221");
            when 5059164 => data <= (x"7bd5d6a992568053", x"8fa41a4e6a230669", x"20689582163f57a6", x"7f101981d8a7ad98", x"18fc5e61330ef84d", x"9b5499728a3f395a", x"0bc3e2f4f4f42b53", x"82955fc44dc4f418");
            when 32149177 => data <= (x"73e828ba5982c701", x"bebed4c2c97bd70e", x"dac932ebfb41f9ad", x"8bf6d41be6392816", x"06100facbf510016", x"29a41c4ebe6ca978", x"5cfd367258a4e7bd", x"2165d7b1d8323d33");
            when 29280413 => data <= (x"c41f208f078fda77", x"7c3b5f00b24875c7", x"455fd9a324bcab24", x"b688b6a73d480d82", x"88897572dc9e8050", x"7c1d1de44962c361", x"51d9464d102cbcc1", x"b9fb349eb5da23e0");
            when 858190 => data <= (x"57c28bbb933e3b86", x"7fc039ce2eea7b30", x"9c68b18852ca30e3", x"d7ece45239f23ee0", x"b4f15fbaaf8244f0", x"fb45dc14e1fd302c", x"dddc5b8e8060cea1", x"dad1625928bbae76");
            when 27662930 => data <= (x"a045cb1fce8aa119", x"8d3903ae4cebd26a", x"3aaa219057604d59", x"5d2498767111c8db", x"8f8426d0fdcd7850", x"dc51540ec44982b7", x"01f30a7b843dd1a0", x"50912080dacfe770");
            when 13921702 => data <= (x"66d518ad9188e087", x"92ad2ec642e48f20", x"53e8fec52c242a2c", x"186f7d0b8823fcdd", x"b6e2df7c97df9935", x"3260bb7b6375ca52", x"60db71dbd0184db3", x"c3ce7706f57351ec");
            when 15796725 => data <= (x"73945fd394206a89", x"e63c90f21df22ef7", x"4cf754446e30e8ca", x"ed472a3312e668ad", x"13a11bf8b3ebb73d", x"b7f8326ae2a54f95", x"ae9389fa25f0df6a", x"7301514d803c391e");
            when 23162391 => data <= (x"f5767dce823aaa5c", x"fc64ad5d700ae39b", x"ed27df93a2d6e90d", x"7e7c0a4319903183", x"17f517af8d93cb84", x"aca4c14957882a60", x"1518550ee91b4d5c", x"6592c2fc92c67df6");
            when 11585857 => data <= (x"3ecd03c057889fc9", x"58b06afd63981ad6", x"7bb08a440e49e6f4", x"4ece26209377b8fe", x"0a526562dcfc698f", x"49916083888c93ab", x"2e5fb74210e06b03", x"4496f1ca7e7dcad8");
            when 26768583 => data <= (x"e1c9dcc6c2a7e620", x"045a490866ef4cdc", x"230c0273fd8f1abe", x"6da09fc9dd4d445d", x"94dfbb80fa3ba2c9", x"f53cba0be4d2a094", x"2e6600b5f158e297", x"534c493f2ed56e42");
            when 28002425 => data <= (x"29a27e6816fd6c9c", x"a722e0caf2acd7d6", x"634fac033fe04d86", x"bde80cb89e249c16", x"27067ce1c2260663", x"28fca6e1cd993d1c", x"3e32441977590ddd", x"f92538dbc3d295ef");
            when 12508836 => data <= (x"2a061c8f0d1c17ad", x"3248cb7a62fb3bcc", x"9b6f2e0d14a90c61", x"6c030739092d9b5c", x"f7020378c0b35f26", x"2313ca86772694cf", x"47e59e5e26c349dc", x"d62c78b80d46571f");
            when 29140434 => data <= (x"2c5b3300311a54e7", x"34f92fd23405689f", x"a1d3aea4a9544875", x"f2f8f0681aabc9d8", x"9af53edaf3ba41f7", x"958c069845194866", x"bd2bb5e18ce26db0", x"519d8b8550d6bdf9");
            when 6551370 => data <= (x"5095679d88f85eb4", x"71257256fc2af17c", x"7726305ec7690305", x"a5b11ada711b5c06", x"1dca99a8a39791cf", x"6b257fc370a2378d", x"d593f7d5eedb63e2", x"052ca673dbc25918");
            when 32862526 => data <= (x"ad7bc9c2c65be3b8", x"7e4c730fa3e5c79d", x"e378521f7478e802", x"4c0f545de8221c3a", x"a68e807d3a7b856d", x"c7cd3bdac2e30fe8", x"a91a5b5fcd871305", x"5cdff4ab284ba3fd");
            when 30020029 => data <= (x"8ae78baf3636a952", x"e98c19d25c4a3bb5", x"4cf1a76421c76903", x"1d75dc34a5538eb0", x"92471973f7f55daf", x"db8c23082d73bf93", x"1c3dd4a4c96ae12d", x"d90c102034115aca");
            when 21324218 => data <= (x"ac3729d4df4bc22d", x"c2ddc7e2264c718a", x"92363061c98df25b", x"54257baebfab66e9", x"5b842ae2f533fcb9", x"9fdc7b2a77d391c1", x"931f9feab4bbabaf", x"a585fa9f307a3288");
            when 811441 => data <= (x"04597e776ea8769f", x"98748c0eab7f4e0d", x"3956d885ea0fd4ff", x"80192b9d84717f11", x"d0336ee6e463114f", x"99b7d10064b32918", x"be4edce96fbae617", x"d3eb1e1650aee4f6");
            when 23751632 => data <= (x"64b12c48a0f4650a", x"6087f3e3232a6b56", x"a7c9dc5f7bc64bed", x"a4374063efde5b76", x"a2276ad7cebf3169", x"640410f416fb468c", x"4de0fc7ec5e252e3", x"c0da351b879521ca");
            when 33989730 => data <= (x"3bb38dac18c0b501", x"f194df06d779357a", x"0f2f6dc57ca49aa7", x"76fecf6a5b218feb", x"be597ba0075eb9ee", x"900d8d23299bdd81", x"f1b464b9043d8fe5", x"047b1b4efa4abc39");
            when 13254636 => data <= (x"cbf2b4f006bbc152", x"4ade14a5708bb283", x"92ff46a139fbf261", x"9cc548c4bf7c0e74", x"a2e93f3b3239ddce", x"f797581a3812648a", x"80af388cb191c308", x"1a2c5e51d93da588");
            when 17186318 => data <= (x"304eab00055a30cc", x"b4647a211b0b5d80", x"f5d7005d6a6ff673", x"08f308d5a72c89b6", x"062cf50bccea288f", x"9be0f0d500aa1fa3", x"69eb6759a19ad7fd", x"ee848a753b04e0e9");
            when 2122783 => data <= (x"c4569a09a7446b63", x"36eb1fb8f8b47b67", x"548bc00931321946", x"6a68b6e968d18351", x"9c3ccf957fc55a1e", x"bcb82c21512adc1d", x"d37fa02018ebcce7", x"0c125a7734a819c4");
            when 10690123 => data <= (x"30835a13674082e8", x"5508c0c38e4a4ec0", x"7ab126e04ed167b8", x"11697a734d227d11", x"f0207b33dc022408", x"24ba797bf26ae6bd", x"7598a1ec910dc554", x"d71d8975ff90d841");
            when 21895117 => data <= (x"e2ca17fa8f9619d4", x"b1e985bd434a04cf", x"a058956be6a069bb", x"2b378b09e591f076", x"9190671313d84a44", x"62160275c1cdef53", x"9529a90ef130db4c", x"f9d2dc5396b019f3");
            when 28055600 => data <= (x"91ae604105163923", x"d09d87158d2f4222", x"81d00aa7f34bcd2d", x"f20f14fa39ec9602", x"bfa2bc2c54920a1e", x"8e623759123e4856", x"009a0942638cb551", x"f75b5f9a7c9c681d");
            when 3524858 => data <= (x"ff03c52d6b8635f4", x"4a6f9def1c97c7e5", x"91edb5aa696d3bac", x"1508e6c6a5fa0874", x"169613749c12d785", x"f8776b4e1bde0a1e", x"0cd1592e493c8d52", x"660fa1b5ae01054b");
            when 19308132 => data <= (x"c63fd40a4cfae5f6", x"ab10ad6e19b59220", x"01cd9858b2833418", x"54f61a5b2a3c1122", x"63ec77f12b2a0313", x"3c3b29ecd46b3e02", x"bdf9006c86556cf0", x"fc350d93e423e956");
            when 9775515 => data <= (x"e200beb07a323e59", x"31b6fcaaafd4ade9", x"c5179f7385263f68", x"17e03c436de2d2f5", x"a6a850c70f8ccb63", x"d88e47511f3cd1a1", x"8c5fe30d67aa4f27", x"04238fe9410bae38");
            when 2837309 => data <= (x"10c6a808dd59b56a", x"c7be1e1b88c70412", x"dbfb680f3693958f", x"f0f6fefae58d91ed", x"4e4b19e663bf15bd", x"f4fd5678a31d3c5d", x"f52ea39976946730", x"6d38dc1071cf7adc");
            when 28669605 => data <= (x"e15a5bc370efcaf2", x"0bb6e173ca3ca5da", x"4cbeb31b480cddc1", x"603aa7c80b823154", x"a4c7f5b61229f0d4", x"61c1e8f8303fe73e", x"4058e2e8624a2d84", x"ea321c03803729f0");
            when 13124664 => data <= (x"450b5d5cc09409da", x"982a1bf3a17ac65e", x"d42a2199d8815df1", x"07e7b3e24674a1e5", x"43c01e18ee584231", x"da3da1a78506ad05", x"fb9250b84f1293e8", x"7789e3b6dbea25eb");
            when 2241873 => data <= (x"a57f220848cb52f9", x"fd110e9529e90461", x"ada2931083c425e3", x"d6270a14a5731c62", x"cf5ab786f8ce3edf", x"ebb09c1aa2a82ff9", x"2002eb9745307228", x"2dd939b0bc1110f7");
            when 15593863 => data <= (x"b55228f5b5dea9c0", x"19ac874d3ebdc870", x"85fcd60b8def2615", x"6eef72e91919aeae", x"a9e9503f43952754", x"6a002387cbc308c4", x"ba97ae332e0a081d", x"3682c975e70b4d71");
            when 12693235 => data <= (x"f93c00fd8d8d3f92", x"770535e9b6e81eba", x"a58c1d74cd87216d", x"2074dd54996e9998", x"bb957968a369653c", x"d7a805c76db82acd", x"9a0fd3c74a0b4877", x"806e4f7dc718cddb");
            when 2057793 => data <= (x"95cd761be75a9ae4", x"c3eeeeae9e06d981", x"c2333a4470a63d73", x"9da8b6802337d55f", x"7967a478724bd643", x"84c8b3d0b146bfd7", x"2960e01fa3461e33", x"5f4437400ae957d7");
            when 30952209 => data <= (x"7b8c12f28bfd0d20", x"190b6e9a2a460b03", x"ae5cd25c50340290", x"2ada9327c80a1ce0", x"a445a0c7b65bec21", x"2750f2a6a034f3d4", x"43ee0eff51a38987", x"c61a2f69abd74c85");
            when 26890155 => data <= (x"988d1fbea17fd714", x"d3a0421c2629ee8a", x"5b2f3c9e3858af76", x"8e7dc1cbbc55e5fe", x"3fd736f79f277d66", x"cb42edc248a2421e", x"d264198fe7daffe3", x"dbc42bc5ebb02337");
            when 15232849 => data <= (x"9be4e77807d70a26", x"de5c67b93be628e5", x"5e51f5862e130550", x"76d44c4bf8ed8dd8", x"a4bf6d1793c0ec73", x"898576f82a13cd32", x"c0330acfa010a371", x"c8da1865a7719d11");
            when 6584364 => data <= (x"3b9f30cd16c2d06e", x"fd7a82262e6fb622", x"f332906d6803b6c4", x"ce7ab600d348cf85", x"9848a8eeeed547ab", x"2522698a5464be65", x"dd65d9e2b145cc60", x"502eeca410854054");
            when 24361635 => data <= (x"ee717ae0b769731e", x"df54d2e8a3a70777", x"d680199d429b6f32", x"41f428c1d9f25ae4", x"b7920a3a9c69ad85", x"23ad0bd2bf49ff10", x"6de36f13b6da9667", x"32b858983126eda8");
            when 6020879 => data <= (x"e639767f2be2edb2", x"b69f8b3bf0c50b81", x"3d074518d4c41e03", x"52ad142fc4fba743", x"615e92664b112ff7", x"a818a30636492265", x"c1bb1b63eb894eb4", x"b9c9ec069ee6de3c");
            when 19959555 => data <= (x"8548528072107c03", x"23f123794f4151bb", x"bad41f4e0152f119", x"e40508672953e324", x"2e1f86ad07301cd6", x"de862f661c187b8c", x"0bb50847c94978ed", x"10a2e7019c554544");
            when 18775466 => data <= (x"2ca2554eb4aa0a0e", x"fe39f50cb694d187", x"5f1d1c485734d970", x"dd28e239d85673d3", x"9fef2fb5260fa64c", x"a0310bebde974a6b", x"dfef49cd63dff8fa", x"e5a5420322b4dc9d");
            when 10034640 => data <= (x"ae9af97b3c38c9e9", x"1302a9a6d039f7df", x"3b3c758bb5dec01a", x"b319bf3480e4d21b", x"a93e6c1e25f8a597", x"2e9a3f98e604eda6", x"2a7eb3df3a038cc7", x"78ef81f20a5bd5b1");
            when 10006926 => data <= (x"d9145892f26fb8c0", x"7b0f4fed70a2c0c3", x"a3d8c1661c3ee566", x"9420d74ccbb84cf9", x"d7e294ad19ff5fe6", x"3b4bc9fff431b190", x"d0580194b3cd5b43", x"bf45af31c33df786");
            when 19807148 => data <= (x"34a151f81dea8317", x"201431fec9455dd0", x"57bc5a107c5aed58", x"60ed44b545eba77f", x"d7e8ffafcb19b045", x"d6b392acc4d3302a", x"4d763f3838c3f3dc", x"067415df296448a1");
            when 23616104 => data <= (x"dea3c082126efeee", x"604aad5c60153a17", x"5fd57b81217c4739", x"27d3c33a0c0be18f", x"a73fe42a11fb45e6", x"b4d53d9fadacea3a", x"5b3213e9fe4866ba", x"1a9f042b55808f32");
            when 5107290 => data <= (x"3087216d0f12bc8c", x"934e37250d0c0de6", x"c2cbcaa1c4501cb8", x"88f00096fd5f91d1", x"3cfa493bdae87500", x"aef14c48e19f562d", x"6ea960c38503ded3", x"994f27dfe6ee9a76");
            when 15079469 => data <= (x"7ad3c62a626d7707", x"9aeab562aad6a326", x"f7f2305cb99787a2", x"81e775b139a419c6", x"f53ac738386298fa", x"c62cfb720097fd4a", x"0dc273a9a2ce9c84", x"af2a5bfda70f093d");
            when 1525485 => data <= (x"76294565c6b37b7f", x"5d4569bbadf2c990", x"f134d5df8f2da7de", x"fa31a5aa3f8ae29e", x"fd9123f6e7e21d15", x"18c524806e329eb0", x"55415de1a48a3a8e", x"1ec9dc578e5dbacb");
            when 18558186 => data <= (x"3644470ff5f0a43e", x"7c3756a753d66ccf", x"3355a8967026e919", x"299df48213694cf0", x"266e2783ed2f7fc6", x"5fc594db0f8f115a", x"8ebf129cd8764541", x"35ec3d7f613eba03");
            when 29095396 => data <= (x"1b665411d35510b7", x"0debe396a2398ffe", x"d83c978842d9e0f6", x"ce2676c88d0525d1", x"098496e353b996c7", x"02b51fa01509a9d1", x"4ca44d3753f5e64e", x"577c3b3bf6100981");
            when 23498831 => data <= (x"4eca7dff0185d2db", x"accf6dd15772ece9", x"8b30c23d4e184b21", x"85fcf4b2980ca01c", x"72791237c03e1b79", x"caa128746e93e55b", x"c4b23405b137b6cf", x"f1fb105881265e7b");
            when 31066072 => data <= (x"3a0e1cfa00b2b594", x"c77474667d176764", x"1e9abff4eafa094a", x"6ca70ae45c585f3b", x"74135b1ea68b5988", x"5169b515e908cf7a", x"ba56bd50988ac04b", x"f2b0efd01430f443");
            when 10394055 => data <= (x"882f5bf0f8f84a6e", x"48b0a2dc89e58570", x"da8195941a58f5b1", x"540a0b737caeb66a", x"2f64b4b302970427", x"b5d1e405d28e3218", x"cd4eec1ca7c48dcf", x"9e1e021aa0f897db");
            when 8349469 => data <= (x"19fe123eaa19f00b", x"12e470d5d8ff7960", x"bed4aad2342406af", x"3794610d1103900f", x"6876279ece48928e", x"ad40f55f95e49aa0", x"c029fbfd5d8a309f", x"dc7b6408d60ebd23");
            when 19754071 => data <= (x"67c2c7c25a5a875d", x"958bfde0b1e3e8aa", x"7c139a8f412c1444", x"f410a8af6bb33491", x"87699b5d10076b15", x"b98d8882cf25fc7c", x"326d4325d94d46f4", x"894ea6da985269c3");
            when 33852697 => data <= (x"0765206c55e80126", x"110866792caa2bda", x"02ac96864b4b74a1", x"3f4a99d226d12bc4", x"c4f48a041d595d7c", x"cd12b3e23775c065", x"4e2792f690a14207", x"0b3972e8a2168e0b");
            when 9239638 => data <= (x"f03c7f768469db73", x"d1a054648784498b", x"c85e005d51919c3f", x"685ed05f26b0c5dc", x"7de8f2986f2ad622", x"f6951fca859db47d", x"75e03740d07a244a", x"12b015cb2a18d817");
            when 31943640 => data <= (x"4b44049bfbf57143", x"6ac41b921f94a6bd", x"cddba5e466fd77cf", x"c036b8b220422818", x"d2e4739cdd66833f", x"5b46f9d2d7c9a211", x"fb52e03c1aa82c53", x"9802e7e95ee7d2b3");
            when 29657994 => data <= (x"58059439a0ae8395", x"cbc6620e18dabc4d", x"3ca2882b1ab8d849", x"78c68846bf79e7c1", x"6aa779952fd02a1a", x"c8c7811099bca813", x"6a45dcfe6766533b", x"483fa1835822a0fd");
            when 10745257 => data <= (x"43bda40c3c5ef1f1", x"22ef132691b09b00", x"5511cdf42cb126e7", x"fef1b78a7ee1b59f", x"458baa2c94fa7ec8", x"54260723d8cfae4f", x"1b8dbd79b6ff621d", x"7a242dcd80bcaf19");
            when 7479510 => data <= (x"65c8e926ebf3467e", x"de3b965bfbe1161e", x"dbf1e3b9411455fb", x"affdaf3f35e0bc4b", x"49eb17d5435f2f9a", x"c6d58269b8d36e33", x"9ed06fc5f8857136", x"87a744ac34f9980f");
            when 18597050 => data <= (x"225c76cd1a980684", x"5a89a6a3a6ad02f9", x"70df46b100eaddde", x"efc0b9aa9f96a3b0", x"c4aea98f8b7b7624", x"914a9a552d89d07d", x"0410b84c978c6c1a", x"7923e71b05fddac0");
            when 19808828 => data <= (x"68257141faedc69a", x"3349a2d00f8a6140", x"8b633a770a33bf11", x"65f15761e40815df", x"f0cc02c7d67d9dbc", x"418ea1857295754a", x"fcd107050d7b3691", x"b8fa0856e580ec4c");
            when 8759264 => data <= (x"a074f796e646ae51", x"b71cd49ce9f93923", x"1a66b89c9f457997", x"795e34be04514b35", x"3f5c1ee84e06b9ee", x"77827202cfeea69f", x"da2205c4122b002f", x"11e3e750f8903ff8");
            when 17633625 => data <= (x"abc97fb117efa016", x"68cc79009cef5b52", x"f005a2d2728ec7a2", x"8d52070c791df5d6", x"5426e61c292f3ceb", x"582dfb1d18324e23", x"d4d78e3c0eaacacc", x"415071b868236680");
            when 28560501 => data <= (x"88fd30fd8c6d750e", x"4fc93600091e9a79", x"17e7bcc50a22f8ec", x"308bbbee96640d81", x"0fa6fc2f0ec83780", x"57d5497f9e1f3e52", x"c33347a32575d6d6", x"18dc0db4376cb4a2");
            when 27454235 => data <= (x"86f0374fe6063cda", x"0f2154ab5c365c8b", x"7a0d73d0c27aeee0", x"bc1cc111ea0e8dd4", x"dd1bb7b7554b4922", x"cd0803886f6a5a5f", x"da9e7c07195df454", x"0fcda4ac5f69e5d5");
            when 14746576 => data <= (x"4c6edccdffa624f0", x"f075c69459b3bd68", x"8a9ab8a1c8c7676e", x"102dca9d7212e1cd", x"c78c41979ae6d17f", x"dd5bf8e075433d85", x"148770b36349abf2", x"f11b06e4fe4d4ff9");
            when 28185643 => data <= (x"a34831bd371b8ed1", x"d77089a006e9b3ac", x"9bd48bca934290e9", x"dbc41bb6aaf18a32", x"3f3b0593608a5ee2", x"0be8e8563534bba9", x"79fcfc94a42be272", x"e32991b4a2e3aeb2");
            when 5130709 => data <= (x"0c048ad6f1cbd458", x"699681eaeae565cc", x"9586ad7e96dad949", x"a3758e79fcb19ce2", x"756ca94433027544", x"5e5c62870f253ec0", x"f5897a63006948ca", x"473a338b080cbceb");
            when 33882945 => data <= (x"c2a99d9d1dc8a34c", x"eeaa7828e5b36c17", x"4c2df22a25167506", x"8b5f8acea10aa1d3", x"12a13bb00c0623d8", x"2c0b765b893228ef", x"29e1b8579deaa086", x"6c3a4515930d9782");
            when 14581499 => data <= (x"64f7fc15fc83b819", x"1e1450692a7dc2c3", x"df5946868a2950d8", x"b9521ef474b67409", x"e8d87bf1375396bb", x"c97e694139f85352", x"03c5d5ab395935fd", x"ee340b63d6ac0eaa");
            when 24544700 => data <= (x"8c3d7922db305543", x"523999b03004eda5", x"852db90dc8e18bc6", x"228fe95fdcc456f5", x"778eb32ae16dbfe4", x"c5e051df11985561", x"2992444b4db96029", x"15378d9c748d8054");
            when 14283410 => data <= (x"a387234cf27a66cf", x"7184a30fb566200e", x"c972418909392e5e", x"bcbdc29be73b84a0", x"f7435164c5250ef7", x"2d6051f48b34bc12", x"663de5b44bf51ef5", x"e8415b9005da5f43");
            when 25396745 => data <= (x"b011c49ebe97b7e5", x"14f325d0d4050785", x"1cac08bf018098bf", x"24506c9a59fe16df", x"792d766cb8f639b5", x"a690009706c515af", x"a3d01452fb9e5d4c", x"6a512c5c720fd43f");
            when 7267669 => data <= (x"f64f969acd09a241", x"fccf485ae16d0d98", x"be46d401299d1179", x"fa6f906be6121b05", x"0f62afed89f66fd5", x"94dba467c9545fea", x"9e9f88355c206a8b", x"3eccf35b40db0de7");
            when 28134407 => data <= (x"de6352ef47586a2e", x"5f2d72f46c823149", x"bc7f8390d008428b", x"24876da0646bf79c", x"0340bcc8b52c9d8a", x"566a4becc5c7b8ea", x"0b3b37ed421d2770", x"8ab6e15a07e9ebd1");
            when 28187920 => data <= (x"2045e18d94fe62f7", x"2a007c6513f5ed54", x"2863dcfd661f311e", x"9716d5a6744e958d", x"183e4ef8b8c743b2", x"b020ac673af4671a", x"587719afb3027d8d", x"a678782798f415a0");
            when 12992602 => data <= (x"f8af142e269c70bd", x"70b0a101b62afdfa", x"2bfb2cfb80b6e19f", x"b7f5e2f5a65b2198", x"b014a90825928e16", x"a4da6741703adaba", x"178214053a53f8c6", x"2be2554abde0db9f");
            when 26905446 => data <= (x"baddf1cbf3da4440", x"009d90a426af4190", x"78824c8048a5caaf", x"917883a814465ef3", x"ce98fb1fd1dffb59", x"bc6e9c69239adb46", x"86911ee5334a64cf", x"3e199aa47d4c8ba5");
            when 10159571 => data <= (x"0b7c9fb751dfbe3a", x"6b18c0b791053ac2", x"2f8f335f8a07ba72", x"711b9418be530cef", x"75d674b6a0b6df46", x"22563c265e354516", x"3048023f0531ecb3", x"e8d824098f124acb");
            when 29002443 => data <= (x"afdd796bbdb22ad7", x"f37fe7fcbba1354e", x"5bd4769c32348c8f", x"975e507008a5d5ed", x"d250f90d24c93018", x"75427e1a5a33e454", x"835c411e287aaac1", x"2fbfdd3e4be701b9");
            when 21278409 => data <= (x"891ee1691ac9a89f", x"625025106013e034", x"d03c8e487a0e69d3", x"0fd24abcc75335a3", x"bdd66cdf1f0fa3b8", x"cad93da2f56590f0", x"703de00372dcf800", x"a99695638027c02e");
            when 12943194 => data <= (x"25f706f4e01dbc99", x"63053220e12316e4", x"064e543f8ce96e07", x"3b658a19d97f3332", x"c867783610447bb5", x"456ccba54ae6ee94", x"68c1d75a01287fbe", x"6dc6a65d01382f44");
            when 20253406 => data <= (x"f3132c88dde757d4", x"d6e5da9ef744fc85", x"7bfb728207df3446", x"b930719eb10af9ad", x"ad68908804f5131e", x"7b01401c83057907", x"85aa4d5703d5f8a5", x"655a46e49c46e86a");
            when 12857742 => data <= (x"c30a574412cb6256", x"5f6e8217e60ae9b3", x"b98c83e52ebf9325", x"6ab299d3cff3a10d", x"7331f8db08d32e0a", x"55bad4ad02e8e37d", x"40decf8e5667306d", x"296266d305d803e5");
            when 8733468 => data <= (x"1c516ae66111f46a", x"859f8d229e3f217c", x"80d044955dbbd194", x"664ee3aab768f4c6", x"363131ffa7e94942", x"d2d00f091d8f23ad", x"e747f897e1bf8b86", x"56ed462dc8966e2a");
            when 24844662 => data <= (x"43ef512078a71783", x"7ae965f00a95d4d6", x"13bf28beeb970b0b", x"0283f42035cd937d", x"698a999158c2b5d5", x"0ab134b0d6cd8683", x"c5dd1a0244ea23e3", x"400aca42124a9793");
            when 8766579 => data <= (x"345e506e2fd6f71e", x"97871aa9d1291b61", x"1ae3e3c95093b26a", x"e0dd9e05556b2a83", x"ca1cdb96b769c7ff", x"f47429341aa4bbdd", x"7ecbb381a0b8e1b7", x"cc7b432a06d4a5f1");
            when 23680169 => data <= (x"9acb357d57f4e71f", x"0cbf1413b2d4de70", x"ca1e2d0d19ab5319", x"0b329330347341fa", x"1264f260ff33c067", x"98683d1a16902031", x"bc22aa1efd66da0c", x"749b7e983b0051ae");
            when 26157507 => data <= (x"4cdd6ed5905aabd8", x"d3ae505bea5103fc", x"008b750bd5024e91", x"8256b97e61ca59e6", x"9e31f4ab54912186", x"0e5961d1465f8945", x"2aa0b167e0d248fe", x"56feaa2712b07008");
            when 22750032 => data <= (x"08bff1936eff5cd5", x"64238f1ae227cbc2", x"c7fa7f044e4ee49e", x"b2a2b275054fcfe1", x"53ca33c03840f340", x"507018b2bdcdfbda", x"21aba4b9f533c0c2", x"f13941389e8a50bd");
            when 11043414 => data <= (x"fc96f714ebf69459", x"2ed1e65fcca7708f", x"d5d4a21aeaf36622", x"ca07eb039f1036f4", x"eb50014e5185cbcf", x"61686b731953e7bb", x"5925e4e86604e5f5", x"ecae6a9c90751c71");
            when 5921590 => data <= (x"35e5bf692bae34de", x"9d9c7a4e07783f7e", x"f554a3852f60fbd6", x"75c1ae80f2857ae9", x"bdcb6a5f8915ffe9", x"1309b9e7cbb144e1", x"f1b138ba2c86be57", x"24b9ef050540f62c");
            when 19890900 => data <= (x"e47db4cb99e01096", x"5a2d162424055757", x"ef0117bdaf562eca", x"91fa8859210bedb3", x"918d5e7eebd8618b", x"3d371ebb382929e6", x"932b4b3dcf2313ac", x"c3cab39bd4dde354");
            when 12097237 => data <= (x"ef8cbe68d28bf516", x"63f821cc2bd4ea87", x"378be648cec9d392", x"d591088f6d7d0934", x"e049998fe660ec81", x"250da092dd6c936d", x"aa8c497ef91439a6", x"e8215d08d53bb1ce");
            when 23782222 => data <= (x"f9116948b0f5861e", x"8aaaa091ea1c7661", x"8b7941ee9608fe44", x"288cfa6d71b6f6e0", x"956b777929a893f8", x"02993827acfcbaa4", x"87c74399e7a2ee4a", x"a2d0697480952383");
            when 15207384 => data <= (x"e21acc258a65129d", x"7de3fbd9930181ea", x"2da45d49e2c908df", x"f483a0be668e02f7", x"be272b61e4cab6f2", x"06de779f67369203", x"bf0ab150e145d50e", x"c9dbdbcfa9f2d465");
            when 14329952 => data <= (x"715dff3a9a414b3d", x"16a71b4f30af3a30", x"514aa0b24b40534e", x"034d8c566d9c553a", x"99c4dc859061288d", x"e84e692ce0e638b6", x"bd3dfe95ec3e7f15", x"b5946e5e01c80b36");
            when 3415924 => data <= (x"0e15371a90988c8a", x"46ed81aa157e237c", x"41e3d8a07a72ed08", x"0818a3c7dd4865ed", x"1201f2de51636707", x"42cbba29a729428a", x"25138d131a63de31", x"fc303d794e5ebe76");
            when 15904590 => data <= (x"17c075cc22657aae", x"f7df3333de3402ea", x"7a6cf928a0e8f58a", x"dd8ac527cf1e9111", x"34e24e96f39a40f1", x"9b9d2da81ecb648e", x"8f48cc97e6664136", x"a0be3847ca58ef80");
            when 5713700 => data <= (x"c34f15ff0e6d4742", x"dcea4b8b9ed609fd", x"ba5bd95cbe9cb126", x"df11975fd65820de", x"89a64d99680dd8e1", x"c43faf3f43410761", x"c95723d8422acdec", x"8d6035e9d8461799");
            when 21684081 => data <= (x"1da4cc28810a362f", x"41f8f7bc891310d7", x"578d1529265c0850", x"4b5835b4b546b568", x"42732ec162c92b7d", x"127cb529b36c134d", x"87b111b748166688", x"0db1b23543af50b2");
            when 24839660 => data <= (x"2487af8616561581", x"667c9ccd6ca4987d", x"7929b47ec60844ee", x"2d3abc1cb172d391", x"cbe22e79e2bc374c", x"75de52392df2372b", x"50757e3605160099", x"b75964f6dfd492b8");
            when 13799917 => data <= (x"2a3d1dd89f3cf14f", x"cd39277c93833cdb", x"1da15d13d1fb995b", x"ce38edba7d707259", x"0eba21cf74659699", x"2898eaaf2a5103b7", x"7c553cac96f8bbce", x"8f7c7337d1aa40d3");
            when 5491077 => data <= (x"9a85ecc570a1633d", x"b20d4c4e690ad734", x"21971df95b636558", x"df3903bee79193b4", x"b9591893d5d6e620", x"8c18a9155d594057", x"172b6d73260b6896", x"64ecf3be176fa8a4");
            when 16173997 => data <= (x"be148803db280b71", x"10f06253692e66e5", x"7ad4dc284e3d8fd8", x"9a4c146fe4b4d8d8", x"4d340a70676e4ca1", x"3c66fe7180bdc151", x"e90571317ab2e305", x"1d88cc447e73815d");
            when 5518844 => data <= (x"54e295a01c78f75c", x"22b8f5aae58098f1", x"ccadb546cdc7ddf9", x"ebe4fd3bdb1b931f", x"38f1e9a0a66ecc59", x"93a1db7e3cea1e6c", x"2bdabb52d1dfcd57", x"77e7c70d16d61cea");
            when 16642721 => data <= (x"6e5ad9044ae03d7e", x"6297326147e75d32", x"0a8ff85c13bb62ab", x"5eaef49d6ec2cc6a", x"316f5c32f08c055d", x"a483e04017826574", x"56c638b065eb2482", x"d63c7e5bc63d1127");
            when 30041712 => data <= (x"601fc625cc6af5ab", x"942a92065c5fd1e7", x"c9008d74f048720a", x"f511f6f3b720cd9a", x"0feaf0639be80e82", x"8d4f680b6dc46fe9", x"4b182f8a1621b6a2", x"28381df1c112837b");
            when 9808984 => data <= (x"d273ca89440d1fb0", x"a44d829a3f1ddc87", x"22f7153395bf5db0", x"d14481b1dc92746f", x"b8bc951da3dfcebb", x"b8d240282d73c18c", x"0bb228a57707554c", x"f353a28e1ff0bd79");
            when 2767226 => data <= (x"714f71836f7a7acd", x"c3d799c49b86d782", x"222fce81dd1b1d32", x"7f6eabbe05b68679", x"8938c537a5645b22", x"0b1475e0ae881b6c", x"4db8823eb1bd8379", x"8da6149097327615");
            when 27997071 => data <= (x"d8c04ccbe895f0b3", x"c8be061fd895a6a3", x"d8a50aa6ebb4781e", x"68da27e945baedab", x"30f2bbeffa06f8f1", x"3869943b2031700a", x"b35a108996112227", x"c4ee0d9f57f2a2a5");
            when 16099046 => data <= (x"3e44af1a533ae5b6", x"2798f87ec7051c8a", x"59d5f1c75294f96b", x"c467c91995b2b9eb", x"b22a1fa22a5c62eb", x"fcbfb89bd330b91f", x"a22f4f8e3c957c59", x"e760885d3a554805");
            when 3804641 => data <= (x"dfec4ab036156f7c", x"1f9c2891f40f255c", x"f687c6e89354a497", x"a7ced6a89c874b49", x"fc8cf174da27f598", x"bb66c8bccdea3dee", x"942181ab372d0e51", x"3fcef31e8448bf81");
            when 22518485 => data <= (x"9a90ba0402997e63", x"eb183227dee4af07", x"33b3d8a53c32b99d", x"7dc1c08e8137d2d1", x"9bf65374c2c9bced", x"69968b8e66e2d9b1", x"86fd80e699d7f3f0", x"25f757c0e2b14114");
            when 32006746 => data <= (x"0a7836a126d735d4", x"609c5c0f5a9c3034", x"3eb6c527cbdd9ca5", x"4ee029a595fa1f98", x"35e95ce1ae695825", x"acd6e27394c215c6", x"377b1102fd39d652", x"7d70fe08974aee0c");
            when 13872517 => data <= (x"d20ff3131a355beb", x"bf7a016aeea25a2c", x"7a07ca30f028d4e5", x"f00977dca4d60ffd", x"c26ee6a01200b16e", x"3eec83123f5e140d", x"91e643b8b2e580c4", x"7e34e94b5bb12210");
            when 15707841 => data <= (x"d484322f7d5c9c0c", x"11a7ba943071a68f", x"3fc6f80dd2b060d1", x"90dc9e8bbf55800e", x"b8283faeac920c49", x"2ea56ade6b80061d", x"8135ef83343d9616", x"a91399fc19c613ae");
            when 13940517 => data <= (x"621b6f682ddb1ed0", x"7f5fab7945ef27f6", x"ba3bfe27f350de17", x"3621d95d8eacbaa5", x"b3bf0c8b15cea8c6", x"790d74850b93c9cc", x"beed5518b38c1fb8", x"0115bc1b454aa106");
            when 1315402 => data <= (x"4ef0de4f0ade769f", x"8c18137a12dfe074", x"1bb1b40e027fcb00", x"8327e55b1f28d59a", x"3d044266e8d6a08e", x"38d405baf0cff7c5", x"50bd3b090203d7e7", x"5bb5c40b05608426");
            when 30767245 => data <= (x"49c74d4f6c1d1a8e", x"25bcf101a06edf35", x"f583b9166025d776", x"857923890be3db33", x"bdf8c7cdfb225ace", x"6d9d34a1eac2857e", x"797cb3c283ef1f34", x"413e03b6f1722f77");
            when 14248516 => data <= (x"344e407bd6ef1bf2", x"f69663d723550d6f", x"65345a11e4a61e82", x"49d82909543f2a1e", x"4a81b0023b8cc94d", x"eed9f87a18840621", x"d79d46160f00dbd8", x"b2eb390d5a7e36b4");
            when 29540714 => data <= (x"2e03c63513f9bed6", x"9352066fecb6daf1", x"fe41bb703d869e40", x"9b1d1b82871d1345", x"f308cbdd456cbc67", x"8e3a01f5e0e20206", x"32df61ebfab9b0a1", x"45875881eb508f7a");
            when 16184539 => data <= (x"faab76b96a878c0d", x"d3077ec54f5a82b7", x"b25cc60c8d0c0eb8", x"1b30402ca7ff0f02", x"e6e9860cc6c5d503", x"cb20f1e19565579c", x"fceaa3b89ec7c834", x"62226f694d441fad");
            when 24087839 => data <= (x"dc00d29d9ebbccb2", x"d41b6dad5fb1e2d3", x"649ca1d98043fb8f", x"89d923ab16e78f48", x"b46bdea856b5e860", x"da3303ac1959927f", x"ec6aa5ab12742c26", x"58311d6c9a05a9dc");
            when 12814491 => data <= (x"5b58f92348e193e2", x"fa62da6e81f1d530", x"f0b8cc0923c7807c", x"4ee7d57bbdca0c62", x"4e1f4c8dedb6cf72", x"5735b9a16e5d46d7", x"e41f96b661195101", x"441cd2bd1ad7cf3e");
            when 31280261 => data <= (x"09b24acfb4711134", x"9ec1fc3a1a22e460", x"b4671a81da4c2c57", x"b197225dcfd28f92", x"f565b2c6ba85a5ea", x"6596d5cc9070424b", x"2f9db829d6a8abea", x"8815c915260c3d58");
            when 14287540 => data <= (x"2bbb08c114872e49", x"69bc673b5f8bfd39", x"bc4036c6d8cfc2ae", x"4b02dd8ca851e62f", x"5ff25002e3dcf157", x"f44ddfce3b25292e", x"06216f21178b4986", x"adf05dbe9c13edb7");
            when 3766503 => data <= (x"8f3f58211fe1d929", x"3747e622aec62f59", x"d7a4f2dc6f55f3ae", x"368b56698b165dd0", x"105d608789bdf4d3", x"cdc9cab47dc1b73f", x"4aed669ccbde033e", x"ef28a57bd9304ac6");
            when 25297094 => data <= (x"b8aecc4e14897192", x"8ebca24a486947a5", x"01705cc41877ee83", x"951099daae3219c1", x"ef879f7b20afabfa", x"cecc0498c60d3271", x"5bce92d138e6f6f9", x"2b887e9f2c976efe");
            when 13114242 => data <= (x"ee7611a1ba9e618d", x"ee2f33d2b047366d", x"9fea2563f11d21c6", x"91b7b4bef9c659ed", x"6978089d1e56c970", x"5cacb6def96001ae", x"96eb5199ff09bdf5", x"41eb97cefa492828");
            when 3365882 => data <= (x"b74064b747b7fc7a", x"f4b15a2a9f218960", x"aa04fc8ef438315e", x"4b606432f5e6d30c", x"53b89691ed36ef27", x"68e8a8aa8b38a929", x"0e90783f5dc196b5", x"d507e809f691e82e");
            when 20440024 => data <= (x"7ecf303f48a3bab9", x"20e2e4656e6c2083", x"6e7e953d9c145a97", x"0887f71824181a09", x"0ea6d7bcd7afe7a8", x"08083bc7434d2230", x"cae5550987cabd87", x"cb92d4a1e84ccb4a");
            when 23966415 => data <= (x"e8f3c8cbd9b16c70", x"ddf14e3bb87675f8", x"66b92f12ffa88c35", x"fbeedd1469cfb68f", x"063562d4ee63ec30", x"2302e927d9e2b826", x"8a584c0a8ff90aa7", x"046f28afde54d16e");
            when 20750601 => data <= (x"32ad6736a701e27a", x"9f1c95817ad72b89", x"a1340a40f010b31e", x"0f77dc177483e5c7", x"f597cb3ce5f8bd51", x"c86ecdec32746717", x"97239520015671c0", x"a40a6453110056ca");
            when 32957522 => data <= (x"ad5be3854f89eee6", x"8e5823450559d2de", x"171a1d773721aa64", x"f91090293f586ff5", x"48f213e78787d4e6", x"4b481281e558cf0d", x"30230c1991fa3dae", x"bd13e3b249d67e9d");
            when 23212598 => data <= (x"530802ce144c77eb", x"c6749ff815163b3d", x"62041293e1d56388", x"31ae11c5d61a2ed6", x"921c71f61ca4b431", x"3e5d1f64a7c18db0", x"bfca340954817f7d", x"624048b820ac7c5b");
            when 32174800 => data <= (x"4d977c5b78a4e657", x"aba592dd9b44501e", x"c3e595d1681d5568", x"5240e390d3173d85", x"ad08e88f762a5d1e", x"d1dc14e4b167651e", x"9bf81ebbc3e8e9c9", x"62fa77800b007b11");
            when 1232074 => data <= (x"b158510ddc7abfa1", x"fe0c881324b1dcfd", x"623c3f9b1667939f", x"19489d0930e876cc", x"00713e22176de5ee", x"1f34e8c3694f0c23", x"21cbbddf33217ec3", x"a59a276209c5f009");
            when 21082784 => data <= (x"5bd816c32ecca60a", x"ef9a14844b1fc9aa", x"fb5549b828800b7a", x"53c883b36ce83d05", x"1d6dfbcddc25c292", x"e44757ff118f9435", x"0d35f6903c88a412", x"ff1534bf137383e0");
            when 5197098 => data <= (x"494782018e5ee6ed", x"e2e22e5f91bddf96", x"fc78476cd88c5548", x"9f90f8900cc78a7f", x"7a679d4eb79b82c3", x"f62294807729e7bc", x"83e59c5dcc777b09", x"e18d5441b884fccd");
            when 4667097 => data <= (x"7b517dcc42b91c9b", x"c40846047d22f189", x"d5de2fd990cd01e6", x"faaca446d9d8f611", x"20c3c6bd8ae638ef", x"d217c98cda9e6bc2", x"c54d656151c3ac2f", x"30b7d10505037831");
            when 22467145 => data <= (x"67de05ae4fdba9e1", x"119ed03768941079", x"cf880af5c0fdf3c2", x"cd8f5ad982f752f3", x"55da3cf9b9d8513e", x"1f006bfdecb89d7b", x"ee3f62cccac8aa7b", x"74f7a252121441c2");
            when 13669552 => data <= (x"c578ed2258c6433b", x"02724378d78f83c9", x"c7034c6c1e259ebb", x"f75bcd39d8ead58a", x"7049b95b2011f387", x"2e9478a608826a9a", x"2ec0aec90caeb91b", x"43134ab0b6e5b342");
            when 29118984 => data <= (x"77826f2fcd9cd556", x"a8b5524ffe275904", x"07ad47fbb06d8910", x"0d1487c230bf97fb", x"8a820bc51219105e", x"68c71cb0ec475da6", x"00726827c82e0d92", x"a4d688bdfb4e4160");
            when 21547586 => data <= (x"9fada1ea763201ff", x"62ca1272e5f3f5da", x"14cc99561556fe00", x"85027594aeffa811", x"23f9f38110cf13f8", x"2dae7658a6147948", x"16b23cc77c63745e", x"060f7902d131b490");
            when 13730376 => data <= (x"6c6bd3ff450f252c", x"d118a5b5ed7b885e", x"e263493658879dfb", x"9a5d12e0022cfe1c", x"d4ff188e08217ad0", x"708c95522790844d", x"8ec440224a6aa300", x"ae2366ed572dbae9");
            when 9609731 => data <= (x"4ecf673552021bcc", x"2df926f7d026c350", x"2f4e0f2444a22054", x"20f74be47a4c5786", x"8aacc51b55690cb6", x"e4ca67676e514c41", x"bc576a2f55086f4f", x"7b73b93f2805e44a");
            when 30299900 => data <= (x"d732ca46eb7856d0", x"63273aed3e99e533", x"7c41a03f81d2fe61", x"dcd052e69bcc8e35", x"0c07f24845bfd472", x"7628b5ba0b2b5404", x"c4c282985b4b2add", x"e3d6d9b070901016");
            when 28128225 => data <= (x"491731ad4130df74", x"a9eeff4de1fbca42", x"ea5fcd8cda3b1e9f", x"56ea01eb64c6f800", x"cc1519844d62e05a", x"5fcc7c4246598a42", x"134cd7f4e6bd0a2f", x"fa956740192fa420");
            when 30763586 => data <= (x"326c6695ce6884dd", x"0f1c8314171718e3", x"eaec559b95cbc3f9", x"15025a4ab22aacdf", x"97e42d8777dd9ccf", x"b1ee75fad076593d", x"35cee7befc8675e0", x"500c4b58cfd576d9");
            when 21352981 => data <= (x"305f6539f491f54e", x"6354c33d66d6bf62", x"c4b9894c92f3e842", x"cbedbd9c8b6f2b19", x"9ef5b531522b9cd4", x"17355bff323170d0", x"385db9b01f9858d9", x"064ce03ba63e7d5f");
            when 7846684 => data <= (x"2baa99fec72994cd", x"bc54234d4cb0544e", x"1fcf681968606712", x"af67c9693b5c58be", x"7abb570f3ed5c7ee", x"ca1bf0a6a99e3f3e", x"8a1155b14967e840", x"26f7246f78d115cc");
            when 12860538 => data <= (x"684ddd7ca0a08c96", x"254a1b8e89507657", x"cd08e49ffb5ec7da", x"c6263ac74259a640", x"183f4a35a30b506b", x"26413cb1211f6d1e", x"acca500e8f2be6fa", x"2268283971e84308");
            when 6021740 => data <= (x"53246c3513dda2d1", x"7c4a77a501f2e0e8", x"a0522964fcd4c291", x"d95a6211dd4cf167", x"182645b555449f83", x"5f699bb2460b2816", x"dba04b435a33dacb", x"6eb58413dc48c41a");
            when 4420015 => data <= (x"7b3c54aa87070206", x"4477b78cb92fe425", x"3b79b02250c6de3c", x"586677ece333a15c", x"d77134f030872f21", x"1ee01d47f7f4b68d", x"083040a97f7d616c", x"34ee0cf3ac2f7177");
            when 29681790 => data <= (x"d198426d1c1c9607", x"850aba135b4abc57", x"49ce30a0d69e3d94", x"680e6c2212a0517b", x"6070c3188acc2584", x"8db26a6d0a562aa2", x"d7e68d737fef6d64", x"3a854b63ea311832");
            when 7162040 => data <= (x"a136070968389370", x"8474929557489745", x"399b721c7c73a658", x"71e0469c42d223ad", x"85a4d08ad4df56a7", x"7352c5454b2b5296", x"33ed37d4abd30d5f", x"b1ac94000941c845");
            when 18258138 => data <= (x"07f82958249a9092", x"3fc1a73acb353bb5", x"643e75abbdbc0637", x"13db7f9a47d4db51", x"9099da59b8d5b74c", x"0e2565f731f2750f", x"b9c8df10b17c4777", x"6de06e2827664691");
            when 31554189 => data <= (x"3b2e86758c2c306d", x"bf89e8e939179b0a", x"bfe9140fa9c07315", x"e48be1b2355f7358", x"35377373acec4753", x"a5931d5b2cca2f44", x"c93b57a5d92dce51", x"7caeb2a633d42336");
            when 1252831 => data <= (x"19b7f2ea00499de5", x"da514d0f454f8748", x"b033e3e02063df20", x"36afad1bc6fbf189", x"d1c4b62a89ee41e8", x"43bbd2d30e33f69c", x"7fb122c04a672516", x"71153ce50af49012");
            when 19333064 => data <= (x"f8f027951f2dbb66", x"a22a8d8bf34c7dc7", x"5ab118267bd86d2b", x"702c0b664f05b08c", x"9be2aa70b6b01594", x"a1d3b9109819eb6f", x"9989db34e203d50c", x"7e4a8e96a6d39ce0");
            when 26826545 => data <= (x"50f9707bb189eb2e", x"0f16342f5a4108b3", x"3990748f7a5fd242", x"322ce7837174cac1", x"543dc002df1f62a7", x"d807d3132f638658", x"a23c57ab583ac783", x"82fbe8c6c8634a73");
            when 30993797 => data <= (x"988f28b48d4e6eee", x"9a032531fcba2f3d", x"8c6296fa1bfb649a", x"9f491671d8aad223", x"03aa219d38834c3b", x"8e5355e6a3061a67", x"5cbfa9fe6dc9f41e", x"a9b3c0d27f1a32bb");
            when 13037242 => data <= (x"8b44d148531e41ca", x"98d44f8183faffbb", x"fcaf127f2ed800da", x"9e9784523f9325cb", x"0874b40d48cd8ccb", x"eef520232f17f4fe", x"e50e1d96b525a657", x"c264317d8f570f50");
            when 6039603 => data <= (x"fd08beb5543c35dd", x"376cf5847455926a", x"be2eacd2363cb7e0", x"e68dbf2c4a95986b", x"064eaa441c0634bf", x"25b38426c641ce94", x"4032a3311eab1868", x"6ff7d88f69e8d530");
            when 31675309 => data <= (x"c41a61a90e4d555d", x"99991a9b6327d27b", x"8d771b493f1c1084", x"d3ef6c0ea04fddb3", x"b0a2bad5f7ca3522", x"cd10fa0039e9fd06", x"350bd13027b4cb8c", x"341d9e59f569089c");
            when 21749301 => data <= (x"3739603b989b5ae4", x"dcf1a37238ace757", x"ce95a7e86c03dcc2", x"5824d3803dfc74b9", x"5051f69de1fe50c9", x"2e22bfe183755265", x"58e4a0729c22e9bd", x"2cf6e714ffb41b12");
            when 31955343 => data <= (x"9f27a2152e42e49a", x"cdc6f29db766ff25", x"96423a0af0e1b036", x"0a0b38e5a59ddf5b", x"e3b9dcffec2799bd", x"891106f401c01e57", x"3f7445aa20fd6ad0", x"442accdb246b4048");
            when 33299158 => data <= (x"d763b5f198565910", x"95ad1d0cb67b8602", x"927ff707d8584130", x"68be861a79ad047b", x"f967845c454857db", x"905d27a28d41f5cb", x"3e905cd76a8278e8", x"ad20480d72073776");
            when 30569884 => data <= (x"948026b230935211", x"ded8d1452f8ec56f", x"dfe7f552b3316843", x"522078562972191b", x"3e043201480e5733", x"716ec59bf475ffbe", x"cdf5e794277af363", x"0e119052728e01de");
            when 11277112 => data <= (x"45306c38df2fd578", x"b717edd39c255015", x"e0de5842f279c4c8", x"d358cc90fa79a1fa", x"a0c3b6449b3cc48d", x"baae6d2f3ec2029b", x"56a23b30871e63e4", x"3a8b77d69611dd1f");
            when 21848401 => data <= (x"644d38d3e9e516b5", x"7bb8aee6b09707a7", x"fdcd9aa6b0393eb2", x"85f109c11d9dba5b", x"e33e55d0165543f6", x"2b88a4b60584ebd0", x"c0725a709d2beba9", x"cb21cb7196b8f219");
            when 23726599 => data <= (x"9cbd5bd4c38eb64d", x"4efd1118f940a39e", x"001d2a4e7585c2cd", x"ba8be770297100ba", x"5a1403ede834c197", x"4aa8441ecae5f196", x"ab3a88e6e703bfbe", x"5319ada91fa9ed8d");
            when 25720420 => data <= (x"a2fad6a1a7db9b54", x"8c6dbc4ebda8a94f", x"23a9436bf19900a0", x"7c2896549212f7a8", x"8c8ee9f3901c23c8", x"81078e9894bf178f", x"97e1b329d1dfbd14", x"cd8b6f94a1bea35d");
            when 4898775 => data <= (x"e65f057b769c2ba8", x"4d75a5f5b8a997c9", x"a462e7d19f35e93b", x"69cfbf5ee8cc4b58", x"67e2000c9288ff62", x"01eb30de85884f66", x"a78d90fe85ca6e90", x"14d0e15d72e37768");
            when 33238254 => data <= (x"2e041ceac216471e", x"edd53157f7eb4cd9", x"f11982a472579360", x"29afa80537971377", x"3b689476b2463a4d", x"7228bd1f7cba656b", x"3c1e7a09ea46a1ba", x"70b8603256208799");
            when 18133047 => data <= (x"27237adf0705e999", x"760bc4bbb4e0dcb5", x"f988385afee078e7", x"ab793a4baf48afb5", x"350bceea01b1df75", x"96ac284ea0183cd8", x"6d21d73ac7e789fd", x"b62279035b92ba1a");
            when 16657705 => data <= (x"2d990ec70231d0db", x"7d17a50ebcc2843a", x"a66f2b151b2c8bbf", x"ee2763f2b33e4749", x"522fc3f1eaa4e7b2", x"9d8704906f0fa703", x"bf18d749cdc2d34d", x"12805db09316a2bb");
            when 24228670 => data <= (x"c909134a4df0d5eb", x"f9ef98dae4b99db4", x"73a5583c4b08ec6f", x"58f75218b4d83ed6", x"0debb1bad5175cf2", x"9d606e5163c2244c", x"70c44add2498c277", x"fce7224d023a2b36");
            when 10129229 => data <= (x"296c36b967402594", x"dc33b4df5f7bf68d", x"26eaf1e40b7d3145", x"d34b8caa0b281714", x"b40ad61b760d25ee", x"583267374381b353", x"88d4894216d6fedc", x"c651727813b20c8e");
            when 21729489 => data <= (x"740cb1ebc88fae6d", x"b6357546b15e9616", x"cbe4e083d438038a", x"fcaa7db653c9e823", x"8be0da4ef0590e61", x"17076464b9d58e7e", x"ff2ae74367356147", x"ac543ef10018ce17");
            when 3967176 => data <= (x"7b0bd0521e02b28d", x"5e03001aea23b52f", x"781fa8fcaf6a5f24", x"2e18198cd447d703", x"f85eb05ddd8ef046", x"65622e33203552c2", x"9b8016f69e54792b", x"4e78b62525ab278b");
            when 4459229 => data <= (x"f0a90351b08c1009", x"2162de1026fd9650", x"4cb119b69d04576b", x"2b0566bbf1fe14a7", x"8448160e46f1f7cb", x"f79acb0cc83da02e", x"f1077710203596ca", x"c7993b321442f333");
            when 32871385 => data <= (x"b17d3d453749d987", x"c0e9a9a3046683ec", x"78c8621eb7ac9b36", x"963d319404338cd0", x"cc0e3764e65a36f6", x"e7104cba86f5eabb", x"80152905bea7f06b", x"abd15d162acbc21d");
            when 22606761 => data <= (x"6abb3d6c3a173445", x"d35033b920fa210c", x"4c35ddd890920a9d", x"b9b2e449fa1bb937", x"7fe2ef2edb79e701", x"cc8cc59ff2b13ac7", x"f3e0c3075d7af529", x"54883c4e39310e9b");
            when 14338800 => data <= (x"d1a9481f4489e206", x"40ab902a4a1790ac", x"05d1b4d114ccc5ca", x"74fad7c71811ac67", x"266480c26ccbf49c", x"566fe584617882dd", x"c45f93dbe28ff841", x"a7b075d59a07c62f");
            when 29379008 => data <= (x"fdb59e86a9440655", x"84f29d5f3e10e61f", x"f3d18ba37acbc37e", x"134095855528f856", x"8f099bddb76cae48", x"27fea6e125a5019b", x"11d9b10b9587a2c4", x"2c9dbae4020ed41e");
            when 30520214 => data <= (x"8ec2588d1c2d227c", x"bee418cced77fa76", x"9d05a80a2ba0ccbe", x"08c66a86c550a6af", x"2b80858cb0c9d13a", x"72f550430b411f0e", x"1543d51b281d6ffb", x"ce99921f34371be0");
            when 29006511 => data <= (x"4d95f34c185db800", x"705b5f6e831bf439", x"6faf071ab45c4bb3", x"4078801a0c636423", x"28432749c877cca3", x"ee10784e5b557893", x"b0cf794b3ac0048a", x"70ffb761b47be650");
            when 21215086 => data <= (x"d4e7b7242ce59bc3", x"777d1d78d05cda9c", x"01c216abb3d529f1", x"f5efd9d86ddde8b9", x"594da29b85e91df6", x"ab92dbf719d07b3a", x"374a62c8208bec87", x"8b3d33d9d865e9f7");
            when 25660301 => data <= (x"76d927aa65225b8c", x"a6d906f30535019c", x"53cfdd3ffb817b8b", x"d065a8e63c34d5cd", x"aff12f5c962aea39", x"d3aef548d41e161d", x"35dabe47396e1ea2", x"772091b3fa654945");
            when 25029583 => data <= (x"7db429310218b060", x"8b9cff16eaa4253d", x"0901db296a5c4478", x"05e339616177cb0a", x"4657756306f6cbc7", x"764478af98d97373", x"57b9150f5bf99b60", x"cbbc363d6bf8d32c");
            when 25098483 => data <= (x"4ccf8ae4e355a319", x"8b69513bdbd2ab26", x"3f5c2ec8d74f620e", x"a9d1cc239588bfe4", x"de9f444b7039b8c6", x"c5d6a31a92aa8f08", x"a0cb42b7d9440c10", x"686ae83c148a0696");
            when 6397548 => data <= (x"795e38e8025910d6", x"ecb840b29c9c8f71", x"77703dc096c6937a", x"84aa0e93c37e31d6", x"701756e354185a2c", x"027ac0cf06e376f3", x"ed3ca42e53d90b4e", x"f8177dbecfc4c68b");
            when 6414356 => data <= (x"e907a201c68696e2", x"e28b8c06b8055c19", x"df772b8ab5dece29", x"4de8d3ab416677e6", x"d56c419c94b9e876", x"42bdb1708b832860", x"0b2228078eb3569e", x"9743f7f0f6ea3e2a");
            when 10587021 => data <= (x"d2082dfff76aa0ad", x"30c171a0f3d8a57b", x"ea781817217e0d5a", x"07cc8ba81c1f8773", x"ff6c1add18a365a9", x"888d49ecfbea3550", x"a2c6b172d3782638", x"03097e8747436a9a");
            when 19025355 => data <= (x"e99afb762d75478a", x"65d7630ae706eec1", x"f1697c6dc640bb54", x"97e1243fe142d835", x"626aa337e2c3e9da", x"494061de0efd4f28", x"17ee587c8516d374", x"8f4e980f25807e2c");
            when 12768454 => data <= (x"f042efd7ac3e8554", x"64fcfcc5ecb363c9", x"dd92093efaae9d1d", x"7aaff4cf62d08887", x"6136b1a4a2ae7d1c", x"e265d6b7993e5a08", x"36da4ae53faf09c4", x"0a24617945b24fac");
            when 27984416 => data <= (x"e10a1a340bbfdc0b", x"0a9ca9453406a67e", x"60c201179575baae", x"84c1d5985196a220", x"7df32e9a956f05e1", x"65b6f0a754166285", x"b10a0f74b6d0f06e", x"422a04787d11fdf8");
            when 4631070 => data <= (x"3ad55c0ab67f3636", x"014dfe3bc2f847d3", x"cbf55dd2969be258", x"f0951329774a6440", x"d297bbc6e3853ad6", x"9a99bf65650fb326", x"761358b1607be9ba", x"1a8701052eaac47e");
            when 10829941 => data <= (x"92295fe6456f6ba3", x"44d0e302700b53eb", x"35c66929305e43f6", x"a580d4c972fae35c", x"1dd5e4ff6cdff123", x"86f15301bba35d30", x"f0318161be31e758", x"27c70eb0b80bb3e0");
            when 4945971 => data <= (x"e24ad24a67c02b1b", x"380bcaca3659660e", x"0285f900a374ce20", x"e2ae5518cc692127", x"047bb7b89672ea3b", x"4dc4c13f5a532517", x"651d1db0b4f2ca2e", x"e3616f108ccd2770");
            when 26865610 => data <= (x"1b212308fbac820f", x"5df89d1bca0d5590", x"5c9c204e7c755ee4", x"c0c24b0bf8990942", x"07222b6c1ba3c322", x"08491efa43a1acf7", x"1f365358399cf83f", x"dbdee312f7af60f3");
            when 3424138 => data <= (x"f68d65c44c422fa5", x"7ffba5c252f48e16", x"446ed4043d9ebdf2", x"6b73f95ea94acb35", x"ccb09cd0ce224dd0", x"581646db9a86ee03", x"8fea9d0e3558c3b1", x"9bc80555ac589733");
            when 27975242 => data <= (x"1f77e0b9a12d9e92", x"062e4941e74a5cba", x"c8c87d723333e9f6", x"b906ba9464ec0aed", x"5473866cf4e13a54", x"11ced567e1dd10e9", x"553403853e161271", x"8bd94fc2b36e2531");
            when 2715305 => data <= (x"759722a9617e3e1e", x"90f53bfae6639d5b", x"c245a65df5120505", x"7c745546ed06904e", x"af981b7310abbb1c", x"ab5fdb74f65717cf", x"280ab2f3f20672af", x"021e3f4739e61270");
            when 15169635 => data <= (x"aa9c784e2196f968", x"a0309c70fc307609", x"6be630fd921b7104", x"a56f157bb1e3d4c4", x"96104324badfeb26", x"bd8c07bf9330c010", x"1e44c7b812497235", x"43c670a0d9dd31aa");
            when 9949333 => data <= (x"a07edbbefa050841", x"aeb75b32242a4e70", x"991dd6462d7100d0", x"8374724d570b2f30", x"80170c0581c2d6ea", x"cc1d04c256788097", x"ddbe1df62f026804", x"858e8b43f10123f8");
            when 14705201 => data <= (x"fdbf429e1057c500", x"6f21a5f13c2bd5ca", x"8b6886031abc2cb8", x"447ddcb12c10645b", x"0d2ec8585a9b88f6", x"053bc7c23e89a591", x"cd581d83c47e0b79", x"cf2060ab219a7150");
            when 4885014 => data <= (x"7e1151b691f2c97e", x"dbf5657cda322753", x"2e16b0eadac7566b", x"0e40e5fc32d40b30", x"bf64698ecb4ba609", x"202e128a43830ff8", x"ab3c23183760a94e", x"d1bc736ec7423f12");
            when 9779865 => data <= (x"d8b47bdbbd58dddd", x"db7f76de74d60de0", x"2caa29c3efe7e035", x"beed0727383a5909", x"f32c048b1658233b", x"91661479bb63f96a", x"673395db6d12346f", x"85d0f83d276e3726");
            when 21134183 => data <= (x"bac36e3e4e5aa95d", x"d440b584b5b82235", x"9adb02129213ccca", x"68dd7872440db48d", x"f4e11340ce0fca4e", x"1997b9345e84ae8c", x"06663e53aa243c09", x"80c27012708fe2d5");
            when 4457333 => data <= (x"020b6df731dd8ca8", x"03b2c3a343293b47", x"ef1b9e0db2552813", x"eead25a0e27b58f8", x"b643dc7a85925006", x"c5d0581a541a48f0", x"0643c386b6eb53f6", x"bbcb06773f31139a");
            when 18482679 => data <= (x"801ff89cf085dbdb", x"d16c714b86956f51", x"d73480db9ed7a4ef", x"a9f9db101daa20e7", x"86e7e7326f0b800b", x"9deb1cd8f8e243d0", x"505d71fdad17b970", x"ec31e8d0aaa04283");
            when 32823526 => data <= (x"57e03a278c1db9c0", x"b8bd8cb35ba2535c", x"af0815eaedbfc663", x"8a18340d53b6ac45", x"e05adec05ad8cc73", x"f93aad02c1adb079", x"1ff5611d5e2d8223", x"1e6d39c809130957");
            when 30509957 => data <= (x"0d51111d4a9d8c7e", x"205b17c0c75dc96d", x"7948731de8097f71", x"5355760c886a090a", x"8f3dac5e3c045062", x"edfa9ef105a0135b", x"9dca37308b24b74c", x"04d8896f5be532a2");
            when 15758222 => data <= (x"4d19c810f6ecf91a", x"a7bd6528cd44311f", x"8d00c4991fb46a83", x"dcd69d709fb2ad12", x"da700f2a6019f8f3", x"09fea6f48e2195f5", x"a69fea48843a8b9c", x"c529818069a246b7");
            when 2544973 => data <= (x"2fdb709a4d1713cc", x"625ca4af7a667858", x"562e5fd68f6de500", x"2a5142a42cc1bb79", x"f57cee783ac80d13", x"1fe84657edab2bea", x"c5d87b1cbe8d7072", x"0e265a827b26e900");
            when 17762553 => data <= (x"fb14167e61bfb7a9", x"c96eae68c823b539", x"005bec858c05a00e", x"274d4d0d124df595", x"e6593a33ccfe4f8c", x"00d938ff26750e2f", x"b15835a2cb2a2a19", x"0446a38880317278");
            when 32029442 => data <= (x"9e688c47f2876103", x"b193e5a53e5011ee", x"27348c76f71d33de", x"7c071212d30dbc77", x"4000d0da35605cd1", x"2c86de81c78ec601", x"2d531dc0887faf6b", x"50cc0c057ede3bd4");
            when 29961255 => data <= (x"6ac4f42ebe91aeff", x"4205c984bf82016e", x"fec057b9b8bd78e3", x"1dc3c6cbbdbe0487", x"6bf2455d8b227937", x"630dd3743e930396", x"f120d1cc7eb20808", x"42658b99e4ecaaf1");
            when 19038457 => data <= (x"56df8cccb362c96a", x"4f80194893e7ee89", x"023944d2428567f3", x"26451fc040551e08", x"4926a0eeb28ea255", x"cef0af72e2e4f65a", x"216bf0598364e8fb", x"556443aa9ccac72e");
            when 8204544 => data <= (x"3c4daa33e976b8ff", x"e9dfc67be4374774", x"3faec9a8d31cb9bd", x"d38cbfd0f967eb34", x"b8dee32d0c9750bf", x"28e0b3592ecd5b1b", x"a635c8b3d931042b", x"dc18b79aa8ab71a3");
            when 3321769 => data <= (x"5094eb3c8aca53fe", x"3e6041debbb57f7c", x"7d5e5a91e179df9f", x"4e91a2fbb8b8298b", x"26823b67d672fe56", x"2df8ad6afcab60f3", x"ada65f315ba70ff9", x"1cf692b6ff4aeb61");
            when 24462873 => data <= (x"e73e02bb2aef1b31", x"28f9f4153306f9a8", x"381d1c1665de3454", x"782a891435209635", x"9e6893818222a0d0", x"21070bc96e100156", x"d9015f95cc0c5818", x"7d927f6cb21a042d");
            when 15624642 => data <= (x"d8f6d4258ff9f3d4", x"840085a654c2325a", x"db9813b2eeb1df48", x"2549d3a7cbb34ffe", x"2b6dfef64e570e79", x"1b6093598a01566e", x"6f39f86c5eb6a9f6", x"2b970558507b55f8");
            when 18386435 => data <= (x"b98c30a295823b2b", x"bedaad951ad1a709", x"1c9cbb542fcbaf61", x"ab0044181b0352d7", x"cb0e4afe840cc9ed", x"3e462ce860d44a7d", x"1e6a38d480099f1e", x"4c1a9b4113cbc09d");
            when 1290224 => data <= (x"6d6e09f5d3c673a1", x"863012b7de8f97e2", x"aa9043cca8dc6706", x"bb828ee0036974a3", x"afa747a2d0ceeada", x"d87d01bdd747d239", x"c84799db7b18c48a", x"ba011a839b0aae5c");
            when 6216141 => data <= (x"9aea8485cff835fd", x"c8bdee6dfb0a0e37", x"7c98b9981a3ab163", x"ef5e7cc6a6dd8bf5", x"d7ba44ee5f52d1d3", x"0ba3537be542e414", x"f22041125036559c", x"8b04669aa35f6946");
            when 9859934 => data <= (x"19ac5be403f9cd43", x"1f61b0b5789473fd", x"78ac70a6b414dcc8", x"b869b43843a1139f", x"b2e735601b1391af", x"683952e6ace7d6eb", x"884d1eeeaac06295", x"2b40a051c3779892");
            when 33071331 => data <= (x"1c999ffffafb8060", x"3967c91b2dda2f63", x"4d08bc42364f480c", x"a8f73465c0d05796", x"143dea016a1e8c40", x"785f8e905eae8b2c", x"a6bc8070ecc06212", x"f83a1c89ed4115e3");
            when 12712220 => data <= (x"66657e708e7b3848", x"8ac22ad49edd04aa", x"5ad3c43575892624", x"f20221c271e6d31a", x"44d9fda5277039a3", x"3b0737459fe77dd8", x"c2f7f8263f7efda5", x"e1785142529da671");
            when 14041486 => data <= (x"e4da9cf4496ded71", x"3be989a3cac34170", x"af5827a38ba25b17", x"7b393e32714fa1bd", x"33086c602dce9929", x"a476bf105653c308", x"55a7ecc9864473b4", x"a06b348341bae384");
            when 18502382 => data <= (x"08437ab3dfdbeb75", x"a1c3f373ee808ccb", x"bbed7292625597b3", x"a7b6ca01ef0a374f", x"d3200fa973811fa7", x"47c1cd0ad39d8fb6", x"256efa9e76c88c6e", x"5de4733137af9296");
            when 27087356 => data <= (x"ceed7798042d719f", x"22dd4a3a15e6e789", x"63a2962c101d0442", x"d3cac4b59be74863", x"bfd1978ee6d7e6f5", x"1fcb597a5f019cd1", x"8fc8f33760086ef0", x"63000a7714ad6952");
            when 6146128 => data <= (x"c76d3a3b9cf93d64", x"0f87a54bb16e2d7e", x"448d9f841f0e3aee", x"6eda9ea56b961f06", x"d53c38648bf5d77f", x"719c6bd1ad39da9b", x"878c321b8cfdb63d", x"c53a1b5be2c884ad");
            when 24713943 => data <= (x"6c560b1fe8e8ca68", x"7cf76cb3421224a5", x"e55d0a2b8095c270", x"5c7e689863f57e31", x"25b1758ba7020d6f", x"31122a95ede01bef", x"b81e1864f9270f4e", x"61911d29528910ea");
            when 30277637 => data <= (x"1f80d3a5d343f4eb", x"908cc9eeeeeb8b9a", x"2a30505c8b3774ae", x"59c2d05f7991ea1e", x"f95f3d97d2882662", x"54dbee7fef80603a", x"27b4b11436238283", x"27a597cbf0309e63");
            when 9163461 => data <= (x"7247329388a554a3", x"804013bf598e7e5b", x"4523c5ecdb2d65ec", x"59d4aa2e9fd7044e", x"90cd760f393129a6", x"2762f5c3b6d984db", x"1ff2daa16e0d3874", x"7abc95837c1006a9");
            when 8304712 => data <= (x"a84b46e453cab740", x"e410f3e543cf628e", x"3e12134e46a9dc8a", x"8c2ba5f4a0689a55", x"e627309478bbd675", x"0bbd83fb692cfdaf", x"94b8cd66a0932a6f", x"1ce389ae82a2b5e4");
            when 13490839 => data <= (x"eb556968e681de8f", x"e2265487471116b4", x"4226fee357289297", x"4e8113e199465a61", x"c0ddad4d9bc67460", x"5d3daea7a9e781dc", x"2dfd5afdf80edebd", x"0841f1f444bacbf4");
            when 21879152 => data <= (x"fd7566e19dac2497", x"ea2533a27c3fc7b7", x"55f5ce1d9a8a4042", x"03191f526eac7b0d", x"5fa2740f40143edb", x"08932ebc68cf4ddd", x"535bec57b1aa201e", x"27602891ca384cfe");
            when 22290614 => data <= (x"c9ca07f4627c46d3", x"ac1c301bfe97dcea", x"04b73bd42ee3e353", x"24703d78123684dc", x"e3d527604fb62a8a", x"6ed02a4e0367407e", x"e330103d32ca5ce3", x"8c2de27bf03c59fd");
            when 28152845 => data <= (x"8e0d69c07ff9b756", x"7a7e29b26f13433d", x"7657266efe2a2294", x"97d5c203dd86cd2e", x"b6dfb4fafe419906", x"006bc566afbdb16d", x"abaf6e5202a02d2b", x"08f35c48548262c1");
            when 28259996 => data <= (x"adcf0f1eaf38d7d5", x"65902be220a4b06b", x"54b3b13b9aff1fcc", x"dbd55bf017a92f84", x"3622bc1a3daa2d7f", x"e9e4193d743b04dc", x"8104c7046b12cba2", x"8414f94444d9f045");
            when 958825 => data <= (x"c24bf007b152f13c", x"c37bca1e36d8a08a", x"01eb4eea5e187d5e", x"6231575e96b4075d", x"e3a71b14ec288c85", x"9bc561a4c1e60575", x"457eed7e1eb258c9", x"01de9ea6ab465b1c");
            when 33873413 => data <= (x"490b5a5869426612", x"4c72b9793a5dd630", x"3ee05cc402590da8", x"978259011bf554ae", x"bb8bafaf882822b3", x"640a3f653dd9063f", x"a05823478f6db6e6", x"cb32f0d9129e7861");
            when 24129973 => data <= (x"bcc7c735cd806eb4", x"58fc81d68c3dfe50", x"f757fcc6fac5b0c2", x"3065aabda1eec54a", x"374fe6680d84aecb", x"ddfcb5879bbb3e34", x"ef5917c5db1aa6f1", x"ddf37100f762ca18");
            when 832481 => data <= (x"d2fcae9d51ee7fd1", x"cdf08b48629776c2", x"b4311af013d70b99", x"b5253c0c9b400b36", x"38452df3819d8e62", x"0e53e52e1df3fd43", x"e8db76af999a2c12", x"b321216b0fbbd04b");
            when 21620215 => data <= (x"cb4a0e238f4f16b6", x"5a9028d73e1fda97", x"2a86b9ade3078484", x"e791ad845c365ce4", x"949bd1e390db65e0", x"e1ad3d5b0582e67b", x"368d1a2ef9f02a70", x"9d3817166d7e1358");
            when 19626924 => data <= (x"a5652c8d38915a5d", x"2271126a9b373fa3", x"60ad51205dbad94c", x"56cbcc62d62bdc0f", x"d4b7f830a9bf57f0", x"58b6b1f6271db325", x"8225c62b71c9a093", x"1f7cf8e481970c7b");
            when 21261126 => data <= (x"8e1fb34668ad78a8", x"b1f9851ea3300420", x"47f3941d975acd56", x"1089485b7c617142", x"baaca7ebb38ba95c", x"02833f3bbf944f4e", x"92e9c4cae63f26bf", x"9efcb2b710e907a5");
            when 13229302 => data <= (x"240cb6fc1cb57536", x"c0f9ecc62c5137f1", x"16d87a5219efd11f", x"8cb9437f0ae22383", x"85b5e8324320f12f", x"597413fa91085731", x"b15dfc211bb8ce90", x"152eb5cacd833a56");
            when 25101996 => data <= (x"3d6585c70f9a9072", x"ed3ae1b2c5e103b1", x"9e5acd347352a8d8", x"c7f5b4964d364ace", x"5e6ad1e4b5e32dad", x"9191edf02c1f1931", x"b11423885e7c6e15", x"5d8363b37ece075a");
            when 12493486 => data <= (x"0e1d8a39aad237de", x"aa8916725bfd7da3", x"775514268cda70eb", x"6809f331de1243a5", x"b1cd11f2636cea7f", x"5c79e94b57a9488c", x"9767b6ba30690323", x"f711cc39d11227f5");
            when 31777873 => data <= (x"e546887c288fdccf", x"d9f5c46c77c3021c", x"ed9ffe65d8b3b44a", x"450ab861400e1189", x"5709737d876624e1", x"5718a538b5e5b00b", x"d20db1f0f7185372", x"a79076bc275813f8");
            when 6118857 => data <= (x"50d1641ae0f0661b", x"63638ed67096bfdf", x"538c9e7db00b1073", x"fb580773e03cf94b", x"4914f9f10ddbdc25", x"5ad68caf93a3d73a", x"08124116df25e15c", x"2b4c52f8cd706305");
            when 12905522 => data <= (x"30fc235d793758de", x"5f5229bf05a712e2", x"9650cafd0788f57c", x"f854b7d9ba994b9f", x"1bf9d271b55643e6", x"d5a2ce9d0faaa8a8", x"e12771b486a36d40", x"55e6e7c61f3f7a66");
            when 26101093 => data <= (x"da6002dd90845446", x"a046d7534f52e9c2", x"5b2c3410f6aaaeaf", x"660f45353298bb2a", x"25d7d622e3cf7340", x"c80e8c1d2f79070f", x"674f547cb3a2f1ff", x"74e8a7dad1bac70c");
            when 28196374 => data <= (x"988d5194e15f6639", x"a3a83154054df6e9", x"64a574321ede45bb", x"6bdcd158298527d2", x"67c10d8ce2227ad5", x"88f5d0ea7990d3ad", x"d7fd9b578e997521", x"1abb0ef237013ad9");
            when 12235701 => data <= (x"a9ac7f5a6d1c4340", x"76ca66a7ff7ff062", x"5087788718782628", x"217ab77c381f1eb7", x"82b3622b7812a1a3", x"38be55ae56a0bb06", x"dfdeaf8117840b57", x"3290e5ee04efe719");
            when 10482119 => data <= (x"72ea41fe4ef7506b", x"ce80b1268a869c45", x"8ee5d43cf050a867", x"bfddca1a794bd971", x"390563df7ef4d100", x"b73be6f601f6a38b", x"b54318fbfd16ee66", x"5fa73fda34f29c07");
            when 3470364 => data <= (x"5d6b8affa1192c7a", x"b8dd90ab623ce7e1", x"9d441fdd43fe3ae4", x"86ceb37e8db50b3a", x"6fa38c627a66e02e", x"00dd3ed1fd25e569", x"036867552f00ce34", x"fa1415f996f21309");
            when 25380398 => data <= (x"0e666b3c69208e3e", x"77aa3f432294eaf5", x"a12319c54a090836", x"4e9706d3fedee1dc", x"001a5d3bc6776ad2", x"246b4a3185751554", x"85d02282e7f82b0c", x"c0d27b765845f82a");
            when 33543052 => data <= (x"8e1b4ecfeb4fbf4d", x"29adb874942bbf06", x"1947716d1bf58119", x"a1896f671e78edb7", x"41be2fbc1e2fe4fd", x"0a2e71a8b14413c1", x"21a3ae67ed072ef5", x"a6e62428294ce0fd");
            when 23511061 => data <= (x"bfd5c77c9e93fccc", x"810484126cdfb23b", x"1bdb286f3106d6dc", x"ce27b9e531ac4bba", x"29d111e69d1734b0", x"289fb4e1c0717582", x"098aaaa1e97cc175", x"285082d7a4c0a528");
            when 4354979 => data <= (x"72900e99260ba6dd", x"82f75b8a424b93a3", x"7e300c99a400ab9a", x"8381a4054b25322f", x"80137145a8ec75c3", x"bc84f99dfaa18ec4", x"3bf65200a2226202", x"93f249db7debfc7f");
            when 22776819 => data <= (x"af95783929afe842", x"0714f39eed63639e", x"0378ad6fefe24c56", x"2e82afb3405326e4", x"c50e1ad5be91e0f4", x"a48835918b566016", x"f430eceefd945895", x"36f0c929ff3e56f7");
            when 30880467 => data <= (x"66314c8e2193f3c1", x"c896ddf8624608b3", x"766c9d935540baf9", x"06b4e49823939c8d", x"df850ebfa37d2bef", x"db2bd2c49a45d3c2", x"1785c198f6ec63cf", x"3d2f0476fb5866bc");
            when 26622357 => data <= (x"9eff8774db7d5ed4", x"4f4900429f734d64", x"7410723201ae40d2", x"3381918506fa7896", x"5e8a2914477074a7", x"89430ac3908fabce", x"a50bc25ff7d55a41", x"9b1ebf11a046edf4");
            when 3447538 => data <= (x"5ad20fb18075f35e", x"0a5c19668059b110", x"a48154b09d72355f", x"b17fa62fe165a3b5", x"f3fd4a9737e8d8ea", x"0636c55855e6061c", x"f68ddabcaf874430", x"3a54153086673b52");
            when 20709324 => data <= (x"3317face9df0fc6b", x"6127fc8f301d19ed", x"aaf7ae6ab183a9db", x"7457200bb867528a", x"6c901d66ac5495e4", x"425a89f3ffe6b539", x"2b70adf6841c4573", x"a1e41e07c2ffd1fd");
            when 6710997 => data <= (x"ede9252111371724", x"6d6c00bec7b6c2df", x"68c1ba0c819347b4", x"d0e1832b1a9fd03a", x"21f475415664c2bd", x"6dc1d9e9e2049e4b", x"3b4fdf114556d5ba", x"cbc08dc6d8982c67");
            when 4435980 => data <= (x"07c9a9877989226e", x"484fb59e039b4dc9", x"b8e7ab806f2524bd", x"e87c5764c905c77e", x"5a69d2a3b2710179", x"a1c10071d7d6d4df", x"cc23a1aab5f70494", x"6885c1863078c741");
            when 3293647 => data <= (x"085fbb2d9c566526", x"674d1e4c8aaa3899", x"d211c9fa79edb5c1", x"b30cb3205399084c", x"8e3b6c891758b170", x"a3f731e9c3238caa", x"79682d5a9ab29587", x"dd8c534ce65fd476");
            when 15268849 => data <= (x"a6f55bf394dc4eb0", x"ffa71ddb2ea1e2bb", x"79976b5478a14149", x"9c5abd598530ce44", x"48f2c9c56faab7c0", x"34eb1c69e73a6c04", x"a29a0f24fa26ca41", x"c5913d40672f9195");
            when 8011456 => data <= (x"3eb4176de854ad76", x"ac2970fc21b09882", x"ef90fea2e33f6838", x"2bc5c0f03a0b1451", x"0378bcbb93b04fef", x"b22d803487ce403b", x"bcc2a79047d900b9", x"63ca50d672a4a8b6");
            when 6597720 => data <= (x"32da60cf3bb3ad7f", x"29cec959affbc70f", x"f4a312f0f8822b18", x"d552f2bc9f61999c", x"a8cdb0b572131543", x"6c5511bb779d7795", x"1adb76b358484aff", x"0bce107493b6a312");
            when 3359470 => data <= (x"50513852476a15b8", x"f07d2c38a1031c67", x"8c457ed74e83c735", x"21f6c9ca1f278944", x"7c5c52b4ced6c110", x"127ad5d4e291b119", x"fda734c0ce96847c", x"674b2c1d54e2c0d4");
            when 18768032 => data <= (x"af5a604c5ac34bea", x"606e2bb1cf88fa95", x"265178844637d87c", x"b52b13ef3a455458", x"37c134c67ff81d8f", x"a0575f2560afa453", x"370b7e915057b9c3", x"a57e4ad2d3c62594");
            when 3800674 => data <= (x"3a2a22bf69d9d1cb", x"f092634f735d5ed2", x"600d4a734600d321", x"f6d3f0a137c51f88", x"d61cb3b7c0203d7a", x"b6058b3334d9921d", x"a29b4f7bd8bc0947", x"b2fc04d05716b616");
            when 5999607 => data <= (x"f440bc15981bfd8f", x"a787feb388ed25df", x"11ba33ec96acd5a6", x"e079186411f6122b", x"6fb531b468603a9c", x"ced3e8d73b135c64", x"f74ca57bd60afb21", x"c5090d1b557eabbd");
            when 21631801 => data <= (x"11655344d69f26de", x"a1cef5be8db15d90", x"9c9483e83a79fb9a", x"6c5c467ae05c5c79", x"3c3ed8cfce363397", x"e0a82033c00b8c8e", x"b39f6b5c793ee786", x"07d39e5633c2648c");
            when 26593199 => data <= (x"6c96986daace4123", x"7f9126c6bd19f220", x"a01f5ab7291a2863", x"6051478d5e26e859", x"abb1b4702f826610", x"6f378db882735d1c", x"240cba0b5471f71b", x"79f213044300fed3");
            when 4628448 => data <= (x"a66f193eb874a0c3", x"1ecb796eeea9de5c", x"eb5d68ee4e2d62a4", x"e573f1baf30450e0", x"d511bc477cf2bc1e", x"d7e6df475b92374d", x"c8dc87d02af60b81", x"e6e6da25dee11ca0");
            when 1631022 => data <= (x"20805f0d8da26a82", x"b99f302b4742a164", x"720a2f1eba846b7f", x"5bb3190cd24387f9", x"cd41b19b8d610de1", x"0b5fa9716185a15f", x"12eee680e6f3d648", x"fe5cf08460322efa");
            when 22527776 => data <= (x"01575775dc616446", x"b766d3502227d724", x"6c8b9e832aa94fc2", x"27ad3f89b8cf3ebe", x"d8885a0e8ee535e7", x"61f45deab51b306c", x"daa8e7d9e74ca079", x"6308f1b3bde6871a");
            when 28590712 => data <= (x"f013e81a0ae5ad6d", x"b13d102a99981c38", x"eb8829b80e9eadb4", x"d1d88880e9c7ea9d", x"80a8750b4b9ec0c1", x"9a7b3e0f96fb7358", x"eca7f2fd86c44a46", x"08bd9863124ae675");
            when 24385035 => data <= (x"804a1246b6e4b91d", x"5c66584b31a1b452", x"ad12d312b7374769", x"e10e2f5ea949cd36", x"b057391572be8233", x"ba10470c503bc012", x"7d8aa67472d23d1e", x"1140ff0a5cd654bf");
            when 8282558 => data <= (x"90ebb328131d18f2", x"7d58c81fc6effdf5", x"41ee806ef4fdb58d", x"03d531b95975fb49", x"c92f85777ab4d108", x"0a86373a925a9ce8", x"221750afed8dae5e", x"d9b5a53213133c11");
            when 9549653 => data <= (x"c5c20b71bcfb8623", x"94cf775f3a41d60d", x"dca66ce65114a99c", x"751d57ce66a0de60", x"c9d2d470802fce6a", x"2a1de260ef6a7533", x"2903fc11965cb4b2", x"a06ec593dde0b713");
            when 31314915 => data <= (x"95f2f5609be3a7cf", x"f4d1d0f353b9e5a9", x"5908f144bc2f832d", x"2f3333a480ffac6b", x"a9e4ea8df5c5586f", x"398776d8f68a529a", x"bbb251687b8da12b", x"6192a62f92d2352c");
            when 6011694 => data <= (x"ea5951f379a4a351", x"f3f2aa7c48f6ed60", x"cf359506fd881976", x"c4f043ae795997f6", x"a0ae5b6e437948b4", x"01ac596a59d26bf2", x"0d989907094b3b1c", x"e275d877db20d3c7");
            when 28188150 => data <= (x"f4692ca2f0c04b4d", x"b17835b68ad1654d", x"92a9425a71a09b03", x"7c84c56dec1f1aa8", x"b5e1177d04f7f415", x"f6eaa3be66792a95", x"576ebb6e01ae5226", x"33da7204cd4e2f32");
            when 11787805 => data <= (x"8eb055e7afe71204", x"53a59c6f1a964253", x"413b9605561de034", x"840bb618f6941907", x"a00a47fc4bc2e1cd", x"8869447ab9253e13", x"a180d4b793de0785", x"7593206ccef1fccb");
            when 14516470 => data <= (x"e3083f2628667f53", x"89fa9705edade64e", x"10073f262a4f5f64", x"44d124fe33238849", x"a7bde268502d09a4", x"ca9b39a63056d1da", x"9b7c4ff310b851d1", x"b404e90d03e71c0a");
            when 3361245 => data <= (x"2a50a7ea9fc69705", x"d0f15bb000b453d2", x"ba9ab87896b7e760", x"c558418f1585fe31", x"f04607275e667824", x"7045f007772830ab", x"40879e256df56120", x"29890ac88f100646");
            when 33300454 => data <= (x"21862c4d7603bb0b", x"20a5e2132da1783a", x"ba0f733aada17130", x"9eae8c8369e44b9d", x"7eb0a3ad195679f9", x"d5c9a4670473f970", x"c49618d65b0c28ca", x"5810735fe254974d");
            when 15832426 => data <= (x"3508e9b43103cb31", x"ead77b15b0975a71", x"6b18a45a82541223", x"9f33448aeee17f4d", x"c8a41dd396bd37a2", x"2f962a76d0d961a7", x"76baacfebf5ace22", x"e7768b232286cb6e");
            when 4789479 => data <= (x"308a696d26ebd22c", x"a6c7c455c6321a37", x"8ac81464e6eeb7e5", x"e23a81a4cde9bbd2", x"072e7c3f34fad31a", x"6ccf0812d1c9d616", x"8ba3533934d21f24", x"40610632ca8d5b8a");
            when 27795892 => data <= (x"dd3e3610b2628a26", x"fb7d9a0761abf577", x"4b47466b7fe077c6", x"c0647e8fa9fe8b1b", x"110dc87642d87429", x"ecc5c820f3e035b0", x"48c6ce45d5309f52", x"d1afe0cbd00740f5");
            when 23474072 => data <= (x"9a85b03b963f6c1e", x"8b10196ddbb8f287", x"4390a6282cd8c24e", x"877659e293cb96e3", x"57d55bfeccda98bb", x"65cf15c0389323a1", x"c31e2c13daac6b20", x"cb5d4ae5eec0ebd8");
            when 9565403 => data <= (x"48368c51dbdfefb7", x"c114a597285927dc", x"677dea3e26a35f44", x"26d3fc41f6a6db24", x"efe7bd8ed5bb120b", x"bd76a5cafe7795fd", x"5a557f6ebdf0f449", x"e84118819245cc43");
            when 20881742 => data <= (x"7b7bea5f06ed72dd", x"98ec7e6d51a2670e", x"0169b6de2a80a1c1", x"60e29a2e66c58c71", x"00b37f318099d96a", x"fae4aa45a0e5073e", x"b3e7c63f474cc6df", x"af6419743e079955");
            when 20076240 => data <= (x"7e288244fdef3f0c", x"5778270ab6a5179c", x"f06c7b42ffe6f912", x"19c5510e43d7402d", x"db5c7d4107d3c630", x"2ad459f07c0bb62f", x"f24136b5c025a59b", x"45afbf3aa49e3181");
            when 5518443 => data <= (x"9cd06e815f79f776", x"daead1ab92577ea2", x"da1f6082a43eb270", x"655cbd0af29a99b0", x"ec70054dbc538b7a", x"2b88514cee8654d4", x"e2cea69adedda4f0", x"8506cd55a588fe95");
            when 26145178 => data <= (x"52ad86e2ef787058", x"229c5de13e107c7c", x"0e281a03abc9bbb8", x"5900cb1b0c5e0218", x"d74d14c1c6fe4dbf", x"ae4ab06d7dfdc6ae", x"3bf7642139eb13ce", x"dd1450f8be445baf");
            when 32683354 => data <= (x"1e9b0cea353e162f", x"ab87ebe844e3c9f9", x"2c7ab4a974d80eba", x"718c14a61972b7cc", x"bae0cc482eb9b8c8", x"6890d2c5caa9cfac", x"02f016404156d8a7", x"b371e7c9ed65155a");
            when 528560 => data <= (x"bdd5f3f33b6ea744", x"312bffcf56ff812e", x"c12fc6cbeb4fd1fb", x"14d8b66df46bdb86", x"2999cef549563dcf", x"4ef2390fb924422d", x"72f97dc7dd0f6079", x"c7da75706b4052e7");
            when 25191426 => data <= (x"266dad90d25fef2b", x"932328bd4f0b2b36", x"9745c9707243e455", x"98c0525153ae7d42", x"227091f530908f17", x"c5af405261609baf", x"262272b17212f964", x"37b6f3d724cd67e3");
            when 31423439 => data <= (x"a28ddb0d0489b4fb", x"c8e41571da84a33f", x"df0ec1b2c09a1f88", x"058211048b0454fe", x"2d806d1cf3ac64ea", x"7e7c91f71c7bd0f2", x"7e8daef2c44adc87", x"5301c7ef0f3640e9");
            when 8826217 => data <= (x"2659eff8697e7c56", x"c9336417ae9d26a4", x"eb678b7993439185", x"16f5b10231a627dd", x"49fbc856c2600fbf", x"298f4f7c4dbe9611", x"1bfbcd9c80f8dfb5", x"d314234ebf790e68");
            when 15223398 => data <= (x"72c522e1efe5b2b2", x"ef3399f66bab3427", x"c1d88ed28054619e", x"63704f7e165bcc26", x"0ea01b3adf7bc167", x"bc7dc70d364905b1", x"8134c0cd67a057d3", x"c859de2b5a2371f9");
            when 24930867 => data <= (x"a37c3c548caeaf48", x"434f00b218416f06", x"ce4f3e4d837b6f7e", x"66f3c039263e4dea", x"6cf265e58aaaa05f", x"e4b67aacc7546efa", x"b3b5cae372cea429", x"b9dad3c400abc84c");
            when 24263132 => data <= (x"4a48fdd650a4f4f8", x"dd838e50e7111bd5", x"0f26d39683ae9f0e", x"8e2445e1a9856240", x"62f8a810611c6577", x"0d451029768afbb2", x"76a297ee3112568a", x"22c1a7e6c89899e4");
            when 23774368 => data <= (x"19012edb718bf32b", x"cc70a8ad30877c9c", x"401f6853d88f0c31", x"ae7d75f90d73b92d", x"ef6a69d157d2a6bb", x"311fc1057e96baa1", x"465fb684682c8373", x"652d826559eba509");
            when 12755859 => data <= (x"f3b81802e5a8f453", x"abe30e3eef5c6a3e", x"615c6b40181c8b83", x"c80158c3a27f2c69", x"e8064555b0a1720f", x"60f43f4f61dcbf15", x"dca8c32a4e248d3d", x"16a674e50281a8fa");
            when 12734932 => data <= (x"1b63e43d2443433d", x"53ae938d1a5436e9", x"5aa5246783f9ee44", x"c052147c9d837a40", x"7d84dacf4512f28a", x"217c0d52c1cd08ea", x"5d9934367bec074a", x"c74f3fe89316c9a5");
            when 16060408 => data <= (x"65ad4bd40a8dc618", x"78ae7c77c26c7e7a", x"366f78b037b88116", x"c766e502cf17395d", x"2f4f5738c40329cc", x"593679d88e27b770", x"3b7ada29fed86302", x"d6759a6a53b6f523");
            when 18751129 => data <= (x"ab6b3ca6a447ea46", x"ddbeb1bc18d6d875", x"e51e38f3f48f126f", x"9a95c2790f562ac5", x"aff4959d83505bba", x"e96670e735ab55ad", x"9e1d44bd5bd48d08", x"9f31089bf58f64a8");
            when 6862654 => data <= (x"e0905d5bad799274", x"10595fb55f4606d6", x"961a10d861995395", x"dbde0113df8ee24d", x"a7c2b6c0ea30c73f", x"e615aae8373aaed7", x"71b4da1e5dd7ff0a", x"52fdb086d84fcc79");
            when 3321689 => data <= (x"61fefd203742ba9e", x"a603f141547f1817", x"665f2ec8a3ec183d", x"3811fa90c36681a5", x"292f5de2238fb1ef", x"516085e7c6a17f33", x"7bc448e51a057acf", x"a69d414c06a0b9bf");
            when 8304072 => data <= (x"d87652ae1d81b426", x"c42bf9c0cc32ec9d", x"6349f512cf32c60f", x"553fb1222c3b90c2", x"de6a21d400de977b", x"ce80339c29b1c293", x"5fb5b7ac440aeb3e", x"6d5774b51a34a0fb");
            when 31991790 => data <= (x"8faaa7796edf2e85", x"731443c77f17de93", x"22b100521ff94dc1", x"7d21a56a23aef41e", x"0d33a52c696f8ede", x"d3d814e9dde58e2e", x"c5eca3404779765f", x"b66db16d715ba59f");
            when 22602507 => data <= (x"bf5d5e8d8e2963ba", x"e97fd2aa5f8a102a", x"f587dd38f5da5aef", x"2251cfd54a73e821", x"181b09ec69156628", x"fbf20c49a885a87b", x"b788719cd3b68b3a", x"f5f89fae7695c48e");
            when 24025903 => data <= (x"d0e731bd44b6199b", x"32c5810af78df9c4", x"71694f420c770994", x"f7a3f9ad4554737d", x"133d0c95969c9707", x"834e7712b03dcace", x"ae4ec9990353620e", x"3490ea7d2fbe976c");
            when 29393417 => data <= (x"c47505265512817b", x"566c124558e5d177", x"8392b93f412a87e4", x"3a683851a43ba795", x"eb668ec2b1c563b5", x"ed97fc53fc025cd8", x"d7b88d897f3ecef5", x"694e8ccd6a9b0982");
            when 33952504 => data <= (x"9b6bff29f3ed3a0e", x"7e4095ca6f48b18d", x"0d1778aaa3f9ab5e", x"023acd57c50fe4e9", x"587ec2cbd3181de3", x"062f3c016f1d13a5", x"64efcced413c2c0a", x"4e32ef69de740f8b");
            when 27596702 => data <= (x"f0e6f1a0cdd7de1a", x"330245e6a3d1ba81", x"0113f276a1f7d138", x"cfeec531ddeda49f", x"bc8774d3a2ac0345", x"a6e379e1d8840efa", x"96a881c5c0566994", x"71c9d15254e3996a");
            when 19612587 => data <= (x"14256f6841043167", x"f74cfd72060b69c6", x"8af2a0e19d49ec33", x"03392b25d6247db1", x"dcb1b37a78f6e11b", x"8bd89cde7482b00a", x"e875b028f1a05f22", x"abd0373838be4346");
            when 32423537 => data <= (x"3f24dcc0239edc9b", x"e2ed22c1c90c8085", x"cf728f93a08185dd", x"06828712e6fac7f4", x"e4dbc66465af3722", x"7da54661671f19a5", x"b18032e9bb28a891", x"079643587d61f00e");
            when 2647388 => data <= (x"e21b14e234de0174", x"f9e1c3e079f378ed", x"8ae23fddfd9bb189", x"a81c8eaa30a550b9", x"772f9cc4cad395a6", x"d611fdc6abf0b0e2", x"ef4552038000780b", x"a574e1a8a79158c8");
            when 31407062 => data <= (x"ca2b163f0485e235", x"6b762b1080a6f5c6", x"19d5a4f99254b376", x"225ec93231328d31", x"b2cd88e2907fb5c5", x"e1b36c67101f064f", x"d40413759378de5d", x"c3e2eec65aa3d9f3");
            when 13894041 => data <= (x"274b732da0aea940", x"459c57d6a52a6c10", x"7ce79133895b0e13", x"2ff56144151bcaff", x"b85be76a4e0c6b18", x"22e397880512ff0a", x"b2dc748ca474a756", x"cf1fcbfcd3697b81");
            when 11141288 => data <= (x"a0357be0466c66a0", x"54e293c2987d795c", x"576c7d3d50b48268", x"fe5a13264419b340", x"14d1cb5c81d1a63f", x"203278fc29b98150", x"819b0408e6c38b21", x"e2daa95f3da10b36");
            when 33102218 => data <= (x"11b4a893c536ea87", x"f9db355dcd6be9ef", x"5a9f0fec6b102406", x"bdd751ac61afcb5a", x"09f4c64c97f33e33", x"00c6bf78356dd541", x"a52c5ddae83f801b", x"a37ab64ab80b7905");
            when 2048106 => data <= (x"4497795cd50e3185", x"2360a2a1735ab21b", x"7654e872517a839a", x"14e3362d2725b95c", x"f588c41fe61e5120", x"53cb74fd7d013771", x"d7c3fd36828411a9", x"5c2b39b7fa64c791");
            when 19766872 => data <= (x"d618e78573ea0159", x"aabcb8a23631168f", x"14d8acccebfe6804", x"7d5eecab2bb31caf", x"97cc0b92d2c00851", x"4e10919ea9f50405", x"e0af9794ac77d93e", x"015822c396dc63cd");
            when 4281912 => data <= (x"0779c29d532719b2", x"d06e4455858ef46e", x"5ca32f821fc18b9f", x"3fd0c4c48fc80d9a", x"4fe73d72f7057379", x"3214d7ee672d0141", x"2a926d5d98e40fec", x"2095ad30d1b1a850");
            when 23820035 => data <= (x"481205579825907a", x"68623fb085942d50", x"a9b3bc2bdbec941e", x"f5dc659216ba911f", x"927335aa41b6eaa5", x"ddcdaf2c5e3d975e", x"06d943464671430f", x"53d090b5eb65424c");
            when 22452893 => data <= (x"007d49338cf5df7a", x"bd47f3cde2ec0219", x"aec3c7c582ae8d83", x"821e867d5004668e", x"dc529dd5e138b1f7", x"b58a0365fbb9881c", x"97105a6d105aece1", x"9dfa610efb96463d");
            when 33813935 => data <= (x"392a082b1ff96d8a", x"85941be082e77947", x"ab52e763cdcc14a3", x"284c461db5aee771", x"da319b9aa9839d80", x"5938ab030332dbee", x"77073bcf183053e1", x"7408a94713ee1838");
            when 25195025 => data <= (x"cd02bf0bb2258302", x"fe930b486fe883ba", x"5c6437616863421a", x"94db42d35ae8ca8b", x"c8de9cc6da07dc0c", x"259f4bfdfd7047b3", x"11e636836329b4a8", x"956bfe28237ae62d");
            when 31210963 => data <= (x"3c30ab3b07eaeba5", x"e8ba4b3c75afc1d8", x"3aa54f91b60099da", x"950661598883196c", x"65c6456cb5eaf83f", x"0fae51e36d0c7e43", x"cf2cebc0f26184fa", x"2f39b98fe68ffd7c");
            when 7158073 => data <= (x"dcd428ea7ba2deb7", x"1c90205bf20d6b8c", x"7b2f97c43479216c", x"053789ed6326ce03", x"1db65690029a4e13", x"a510bccc314335a1", x"3be523dec54f7824", x"f9afdadce41bef5c");
            when 19203170 => data <= (x"27e9feed1ccb3a13", x"da4ba71811292f81", x"c8d212f19a4fae75", x"bb9930f71f9ca08f", x"1e6c109f3f9880a0", x"0ba4241fa1a4ec5e", x"aa09d74fba8e1478", x"9597f3b142d5e598");
            when 3566397 => data <= (x"302e46c22861663b", x"7f30f25e643a5df6", x"55dab0c7ff8749a2", x"3ca1bc6a76d99efb", x"e58fc6ed41f5cb3f", x"4ed9602b9fd59bb8", x"cf20241980eee99c", x"cad57ca6ea57051f");
            when 18012397 => data <= (x"e129a1ecff9fd62f", x"1759433df7cdbf68", x"65ee9afb2b0baa6b", x"7a870b4270361d63", x"52aa2f6a05ffbf5c", x"e2d1e05909e1cf26", x"6929fce4643d0c39", x"939c00db79ecec9e");
            when 11146391 => data <= (x"a10a7bd855c1b4c7", x"46f468e4f484e272", x"1387aa7f65072219", x"223faa355cfa566f", x"a5acb9d6e901fb5f", x"d7081834334b6768", x"c4800b1d07716180", x"35b6cd1ad071b229");
            when 13803414 => data <= (x"bfcdb6d462ed86e1", x"3f60e28428ab4e0f", x"717488b712d04da8", x"3b19cc5746db9c05", x"5267e8b94138ac6d", x"60760e415423de14", x"37f3469c8b28198d", x"5d0b5e3998cb8b17");
            when 14080149 => data <= (x"a4d0912b5cf33ef8", x"865766f8ed2af867", x"074db710abee5948", x"fce8947b2de3e1df", x"f450d7102f020c2b", x"d400eb760e79a3f6", x"6b2a5c49c6932a8a", x"5c3aeca8f2c6b91b");
            when 30942225 => data <= (x"ace8fe65f91eb531", x"ded45d575580dd43", x"d7bb1442ff29f901", x"e325cb5b3db95b94", x"0c7d9d5334b43dd8", x"3511aefae0625f3c", x"e04e3d3f9d943d4d", x"bb3c2319a8c377fe");
            when 4067356 => data <= (x"a67db7758d40c614", x"5fcb247f38ef6fe9", x"ad55ce15dd9cc299", x"15d79e628aa0709a", x"22d51d4d1772ad1a", x"102aca7cd6f5dcd1", x"5cd1802e95acb0a3", x"c1e18a16fe209caf");
            when 22290207 => data <= (x"eb34d1339b548ce3", x"a5e4e6368e608420", x"d9f8839a34cffe57", x"a0789f8d4626df4f", x"b3ff10ec7dd5fb9e", x"328611c149f7a3de", x"73c6734bc414c574", x"bf8e3b527e417e66");
            when 11316459 => data <= (x"e69e3d76032b7ae6", x"29384bf2db60acd6", x"f2ed715d7616caf0", x"e771ab549fd8d79d", x"a214c8682e1bd3bd", x"9144a7b29b6766ce", x"39474e8be86f4969", x"db91dcf00294f7f6");
            when 31950052 => data <= (x"f02a3e0911ed9b1f", x"5564c80cd7000941", x"3493f016905c05c3", x"ef1d74bb4002f1ef", x"d9fb2727e356d584", x"618ee6e6c046ec85", x"6433bbc1f34cf78b", x"0cbfbf0a1ac33f0f");
            when 9195015 => data <= (x"7e5eaa27506eb946", x"ccfb78f42e11a1bb", x"5b2fc7a246316d4b", x"9c55ea436149a0dc", x"498d30eb4605fde8", x"bba247b71a63616a", x"e17c318b686047c8", x"f2fbffe8ef91c3f5");
            when 5643964 => data <= (x"0453749c942c4a5e", x"865f6b05f94ccfd9", x"c22e1a4cb224914b", x"4751093247d28de2", x"58281117b6cdd79e", x"d68c525ce207df29", x"b6253ce971463a9e", x"3e6a4d60df452cba");
            when 8471833 => data <= (x"aedff1d866d30896", x"cf628721e72e1389", x"80d8f227565f7dcd", x"e7ad8793451dfc11", x"2144bf81b31fc075", x"04eb5ddabec91f15", x"e744e0cf21e98657", x"469fd15ebc99f0a9");
            when 7605174 => data <= (x"f19bf2029eff9fca", x"6665ab92beeb2cbe", x"5e1db12befd09ca0", x"ccfd1aa3f7d7a7c0", x"6fbcbc8e8524e021", x"afeff54e4aa4ca83", x"882356ca921e3b3a", x"48b23c1f730d3332");
            when 11909880 => data <= (x"4798bddeb5b801bd", x"f621e0696cf6f317", x"edee23c03c8bfb36", x"e4474bf5f979b62d", x"efb8a05fe40ba5b1", x"d1b50386383713c5", x"40d503487d4acf7c", x"1a1d2302086de8cf");
            when 1834288 => data <= (x"c4bcfb78cbcc2728", x"dbb847d9834cf96f", x"04d3ef5aa819c623", x"21d3b16f6a64871b", x"0f58902d2754cb51", x"c80365085b2f3b59", x"6f1baa721fdde9e0", x"3cb69080eec09c24");
            when 4111148 => data <= (x"1211008ad4e6c485", x"660be9108f4737a2", x"5c690d03e3fb7001", x"91b8b78a04d95279", x"77d291a7c9dfa124", x"44af2e073c155981", x"8642c28e553f80d2", x"1d131535cf98e9f8");
            when 15073971 => data <= (x"f66ab033ed06d65f", x"b6a1df45360beb4c", x"561f06f44302f40b", x"7076fea70bd67924", x"2801df1ca5c74487", x"d75208a5ef9efa74", x"d5c89b8d6844eb36", x"2afa10e4e1365811");
            when 22009731 => data <= (x"1d1a8a45fd1c0598", x"5887c513d4d254ab", x"eb91dac79b09c64e", x"1c6b8150d540f229", x"ba4910d11f62869d", x"346b301b495b5d0c", x"7f749f9165ff08eb", x"a953c61828deb0a0");
            when 8009240 => data <= (x"7a814d852c8cabfd", x"7ecd0cffeece313b", x"ba36099598816f5b", x"143ebd679a2d3f02", x"5bf7bf774d5bc44b", x"c6a33d0735fb29ee", x"e583e30e80ca54ea", x"5258d654c40841bc");
            when 17400757 => data <= (x"e1ceab3c448ca3ab", x"ca93aa45f3f64655", x"41de1c0d63f91365", x"18167e1c68d6df54", x"edf03049accff2ab", x"70f66987f23ada1c", x"1fa85d23f7feb036", x"ffb5678e55238398");
            when 2437797 => data <= (x"224ac86e58c1000b", x"4bd1aa8f836d85e5", x"df7ba4b3651b3497", x"581fab3096ba6976", x"e5b6f77a6c639472", x"c5fdedc58d75605c", x"da036c97a56f608c", x"51c94e2a8ddf1969");
            when 32028863 => data <= (x"8a02c3d2cdbabcf2", x"f8e2db53fe42ac02", x"11d35bc8ab97ce0c", x"5dedff631e2996d3", x"6c7d7395f209d6df", x"ece4d2a18a67bd05", x"44780dabfdc34e60", x"31d9d5f28631fbdc");
            when 1194275 => data <= (x"adf1e9d340a8019b", x"ecf197eb99c2832e", x"7b5303f4067cbfed", x"8b70e0355710f1c4", x"7d0debc916f152d2", x"a34ed9f0ebc288f6", x"74efae7247cc0a6d", x"b8b8803e9291b55d");
            when 23282767 => data <= (x"8197a6b6484f5c39", x"2b8de04507fb9fa8", x"1fe72f9656fb9ccf", x"d486a80032663747", x"e7b6851ba1a17812", x"bb7272afc6a81045", x"a1e5056ca1a16626", x"bcf6baa6b96c1ab3");
            when 16231389 => data <= (x"e9b8e2c5ebc68716", x"6876eddf6cabaf2e", x"fe42b1c2545f4a6d", x"65480bdfa38cffbb", x"4bfe131338353efd", x"af1f39499960ad9c", x"1d5f97382bf4d9d5", x"736be64e87f7a455");
            when 16457994 => data <= (x"ebd2c00ea616afa5", x"32c9ef4e1ef1de6c", x"83945cda70bef25f", x"3f9729e3b5639733", x"7a7b6c7d8015831d", x"49cdceaec60e2b67", x"9b45abd683c67fb8", x"919ae295d6595a3f");
            when 16651251 => data <= (x"93b860f2557fca12", x"664331c3995fe7e6", x"043d3e330495bda8", x"bed8fe097d648fbd", x"778cc5d45393485d", x"5a222b207d5143a7", x"f9839c0a1c0b5a27", x"357c0315e7a31995");
            when 12567799 => data <= (x"d8179f3d2d310fff", x"5a0a916f93f07693", x"09fbd7abbba10676", x"6c03cb3e54194881", x"f332a0449569acef", x"fb57ed8bd63de0bf", x"f70dab7dded8cb5d", x"a921e5b612ffa3b3");
            when 8167267 => data <= (x"d414570c0b1d88de", x"a583d3abf658f91b", x"239174268febc4b4", x"d25b467a052751ca", x"cbb4a4e615a62d74", x"a47ff4f5d98f2981", x"64911add3cef3236", x"b3904b660cf5a36a");
            when 10665957 => data <= (x"d87fad5636a09205", x"9fc738b222f1c548", x"7d0c2ea33f32eb32", x"ac81d5a07c6be433", x"470554ab3c8db852", x"eaacb0919275df2d", x"becb8c2a2a599ecf", x"d465457c6374729a");
            when 26758239 => data <= (x"d83a3f5101adb487", x"9ccd4a1b382fa905", x"b57b3d30a78c6b75", x"811cce90d6139739", x"cd0512e21aac0e40", x"b6ac44766ee01cad", x"3e76c580f628abef", x"ce2a8dbc50fe97d5");
            when 1869364 => data <= (x"d8ad08415b543bf4", x"484fd8ef94c788d7", x"af8415de86977ecb", x"04855212a100038d", x"6825809f804fc979", x"4adfa4d508bde611", x"51cc760f2f4b9eeb", x"e64ebc0ec609ea19");
            when 23611108 => data <= (x"14b6f91e9c4f6196", x"6cc2d23e3ceb6369", x"6683be2dc10ca326", x"9ba4f0b8736b9f52", x"b7a8fd46e55b634e", x"0b630ce34fccd26f", x"cf7673aec630b4cf", x"64388b2c658ec1e2");
            when 21209567 => data <= (x"c21f6355e5afdf07", x"e686f1de13287b39", x"54f2048bfa9acb48", x"ed763b716a443f49", x"5ddf539222029c9a", x"8179a48af195ef44", x"d6dbfd1aae6e2a44", x"d352959cb42a9dbb");
            when 28159149 => data <= (x"dea9bbebe5c83245", x"83ddcf3037ad0dc3", x"985538c56718c230", x"a03ca4a611222f32", x"2b079361b1959f36", x"e10197d326255b97", x"a313daddba7878dd", x"c54e738113975e5c");
            when 28112677 => data <= (x"2df0aa3a1da82af4", x"c7542a645521e877", x"f22bb705b43442c2", x"204271b5ca465fc1", x"0c44356f4115d901", x"f64bfa4b5fb1af54", x"b94294a6f00931e6", x"4da6b54931e95080");
            when 32365268 => data <= (x"a5a37d27594cccf3", x"f6af3630fbfaf889", x"3d611d1c059e1150", x"4ac733ef0085af9b", x"4ab65e975ebe8f2c", x"58b8f04ba2704f35", x"b40699ea698cc6bc", x"edb4792e6b0880f9");
            when 27084667 => data <= (x"5091c9a78a09fb6b", x"149d01693d7510e8", x"1c57f8d3e4fdb6a4", x"8530f3644a314afa", x"73c01f4196c8f480", x"be71e2222e19dc47", x"1e4b1212765d1b26", x"302cd6db7896f32b");
            when 2299930 => data <= (x"285a9b722c973da3", x"def9b7d8ce39b4ec", x"c14da614582f2eb4", x"a6fa1ee6b39f6e06", x"f1d904df6faa55a6", x"5134e2838915a837", x"f067361edb13880c", x"0e55ffeb6c9c726e");
            when 22807837 => data <= (x"e707b59693498ee6", x"d34293e3f149ab8f", x"23ad18c2ca89629b", x"b02de7432d3a34b2", x"7ba3611d5e173034", x"555e779794aade83", x"1e0c0a3669d88442", x"35c605bd40985ad9");
            when 30266169 => data <= (x"70078284317ce6cc", x"be594c914d9be0d4", x"dee82b2574916833", x"c021e3293f32a08b", x"bfac15e4539bf8dd", x"baa9e75ba3f57b0e", x"a1be164c76e89b7f", x"df9770aace57a0e8");
            when 26827746 => data <= (x"9e9451fda3b083d1", x"8c1f56ebb257db13", x"9e82170fb77a9e13", x"8d5f270b21309fe7", x"db948ff9e35d73a7", x"a922237b57e77e93", x"e826eb27ced3edea", x"a5dfa3527795038a");
            when 24831420 => data <= (x"2ac39c9377fd1d00", x"42d75c726cf21b85", x"a980e82534a2f555", x"b941c56f070d800c", x"a80aade5be490775", x"9e109e4a7371250b", x"6deb60ea2f205b35", x"474edf0f877c3909");
            when 11225950 => data <= (x"dd33d8a5b0232f0f", x"56016653127b5c49", x"a76039146795da8a", x"ed091d9b06b7f260", x"b4249f1d9a266169", x"f8050d0c2da93de5", x"135bb30614b7e167", x"be37c0129254ad9a");
            when 31698596 => data <= (x"0e12cc58b5e84914", x"283167745aa00df7", x"7fa570b13ca03c11", x"ec2da8172814da8b", x"626fd861f314943e", x"1cdbadd6626b4892", x"5401bef8d852a959", x"1b2c18f0994e8c7a");
            when 24601806 => data <= (x"90fb3f8ac7a4c090", x"40a599044b720edc", x"fec68d820e1972c6", x"9485f05506b0c01d", x"cfa544475686894e", x"359c90b7731459c8", x"1f8c6c79e75bdc3e", x"8e5d45068f2e46ad");
            when 11507594 => data <= (x"4b96a47efc0ee8ee", x"b59acb8c76d6c2b1", x"4f45244e7622f90e", x"2629adf6ad70db2e", x"6bc6ba01aa0e58ed", x"b4507048d982c570", x"03d9118974ebdca3", x"857069657cd4e62f");
            when 26945869 => data <= (x"3ba1336c692674f7", x"e81c2c14c6de71ae", x"3efb8f44fbd57f7a", x"dfde4edfdaa6648d", x"5320b12ef98d6501", x"bcc552b5b16dfea0", x"527ab29402c8ac55", x"77d7c1d72dbde6cf");
            when 13186345 => data <= (x"912fdb05a98b60a1", x"63cf9be1559ef442", x"b401fdec2d7cd293", x"403c0476c17bbc83", x"cc738d0bff4c2493", x"f905fcda3ed17202", x"6d2bdf049f1a704c", x"91a5051386bfc023");
            when 29070806 => data <= (x"362b2049c31b8349", x"2b474ebafe2662d3", x"113f13b251bbe94c", x"54c8c5f7a99fc680", x"d85e014792b562ca", x"35284c3f8a1deb52", x"acf9e71017956dcb", x"b26eff14d8004f35");
            when 16271402 => data <= (x"ab46fa6eafc8fd89", x"0dc8c41d7817c4d6", x"e6283bafc4079485", x"3651ede314d415a4", x"99c3c4fe21d5cd2a", x"7d3cbe9558c77dbc", x"accacb9b0213cc10", x"24c634257b1d0898");
            when 29471334 => data <= (x"56e7a546886fb7cb", x"26743db9f514100e", x"7819cbd1a5cf3116", x"7c7bad685709be25", x"77dcbbff660f4ef9", x"23a88dd0b476e930", x"f63a40966e301cae", x"238545997a449f4f");
            when 11688796 => data <= (x"a37b4aa7cdd28696", x"a3593c3d9497963f", x"5ce5ce174a42f36b", x"db3e7e2871bf345d", x"ad10e050e5668622", x"6d51708ca9987364", x"9384bb51d2692708", x"047d835a365b2f25");
            when 2692091 => data <= (x"b865c6ab0fe3550f", x"6a27e1da378557c6", x"a2a016f2e30d9142", x"cb518d7e3b73b54e", x"0f0c3ca2c30b2536", x"516bb711bdc9f78d", x"7c15dd29ebee1618", x"553d4ec53025a7c0");
            when 26400497 => data <= (x"9f95e3ef482f7898", x"958c9a6d3af672e1", x"a90ac7eadee6c055", x"13ccb379e8adeda6", x"1e49e40cbad7ead5", x"f10d75b910c688aa", x"9d6b727bd996bc72", x"3ff0f2deea4bd658");
            when 13463620 => data <= (x"c3495c0638f3f558", x"0d30840af7dfcd33", x"5bc0c2fc8b5e8960", x"5bde14c2bf061c70", x"ab3e53ddc2b829c3", x"da940c01dc7caa9e", x"5bb01b22e7b08ad3", x"2ff4dd2c81b8c224");
            when 21142960 => data <= (x"70a7eadc0bad98ca", x"eba5e25442499233", x"7c6647ff0089f971", x"89039447dd158e76", x"49a44c639f1f20fd", x"da88dabda3d2151e", x"7f6563cac4a37259", x"43d9bfe4ac09201e");
            when 31617024 => data <= (x"b24dc738d3623b0a", x"c7dcce38b017e894", x"01578227aa70921a", x"4d8f83cbe9e2e77c", x"18fccf6684fb01c8", x"3922703640f0f11c", x"2ee91b6ef86b089a", x"6f2f347080c1e8d0");
            when 13619072 => data <= (x"2454c5e261265e94", x"299c1c8933f1b9ed", x"211c575b2bf05280", x"ee063a6fa3775910", x"7ff620d191d06184", x"0be9632b567df5fd", x"4673ea76912d4065", x"e342e7cb4a1b2108");
            when 3762408 => data <= (x"7c0d5694808a3846", x"d15d3b9c4f5ff947", x"fa231d38f25841e9", x"e201bc945707ad11", x"1cb2d9f6f8320dfd", x"d37d5cc3e9b1223f", x"d6fbd78f6e50809e", x"41e74bc021ef7121");
            when 29665016 => data <= (x"28b845d731609915", x"900b256037b21817", x"f15de80deeda6e47", x"814a6bd1db4e7ee0", x"aabefbf9749bb2e4", x"4c744be325c13c72", x"7a81e9957cf7ef4a", x"2dc85c0397044fbb");
            when 866960 => data <= (x"6ea313892f3176e3", x"eee59ec32486f3cf", x"ad13d12b1bcbe42d", x"d6d4f0581e57d3ba", x"6b2a8c88d69fcc08", x"62f9cb9059c7caee", x"ad2ea041fafe936c", x"96f2218d4322f93a");
            when 6321934 => data <= (x"b69ca6e34a4abf59", x"6ffbea61ffe8e119", x"a15eb0512f060cae", x"d1ab1a61c36315d1", x"105173412aeab22f", x"7fbda17a4ea3f721", x"6b08f4ae853b2063", x"b6703d49e31136d1");
            when 21740862 => data <= (x"57b7dbf635e38fda", x"873cffaa4066df7e", x"fd744d06444309c3", x"e672438db68d5311", x"f595c481c646b39e", x"5b50fcff9a920e6d", x"9d02d0c1781c41c0", x"85ca8c8c53b1727a");
            when 33026714 => data <= (x"85c0bea166246872", x"d27595a18da441c4", x"f9f67ce874251a51", x"5fc955d1632e7799", x"b79d830a69330d98", x"51c66aea31d1dec5", x"abef77e3fb7ab6be", x"b3e1257784079033");
            when 11321495 => data <= (x"694a7e66dc889712", x"72c606033ce42264", x"0232e930d4b8681f", x"0f74dcce90526b7b", x"b37ff574e4f044d5", x"d72ce84ef97ec994", x"c6a293d59de52f61", x"dfafb18fc8e282b9");
            when 6150626 => data <= (x"f3a633eba12ba1bb", x"3cba1ed9f2f4c2b5", x"40e9672ed887db40", x"5045c6e63b663dfb", x"0165a718e20044bf", x"5424fd8dfdec672d", x"4a1aa0b0b3d6a854", x"083b6ee00f767740");
            when 12751872 => data <= (x"19db061bdd2890ea", x"0186d1bc40c1c6a5", x"5ae1a3df967f55b9", x"3230eb0fe7640abb", x"8088749bc98dbc16", x"7ee215e9574ddd16", x"7a7b0526a2681b38", x"108f3173604be7e4");
            when 20107838 => data <= (x"87a36b013011add1", x"35c94a0b430a3e10", x"29a56e713474324c", x"6e195e0112a3fd64", x"0039cb5cb8d686b1", x"028a07d6cf34cedd", x"801b5bf2c597d172", x"70fcbc1ceb5229b0");
            when 12529395 => data <= (x"606fb9d4a3a10e50", x"080a0e4f3b5ef76d", x"17e839f11fa3891e", x"600b30670718cda1", x"607e6e5b830417ac", x"e24d7c3b0a313fb8", x"8f0024cefb77e437", x"ed7260a594108cc4");
            when 33765645 => data <= (x"50dc328c6a13a9a3", x"f89d23ce2cc53273", x"44f2917ba8e0a68b", x"5a1cc40de019a422", x"d7fcbbc68bce1d88", x"7c00f8df65fd16f0", x"2a0c2f1c6a37974e", x"07b9da1f25f230d6");
            when 1018201 => data <= (x"c110da2667fd64f2", x"cf70f336886b09d8", x"76ebdff8249f3974", x"e4a6e0c367e6763e", x"fdeddbb0fe65de9c", x"5ab4faae38da7f28", x"db32735a7880e405", x"1b1ec1c2e675998a");
            when 12412496 => data <= (x"42942fce0689e32c", x"ee2acd6be576fa5f", x"fb831cd6e16911c5", x"c0f869a3e4d0c357", x"b703a8366557ca63", x"283497dc147bea65", x"d8335cb5139fc352", x"09914d2eb4e08815");
            when 8828704 => data <= (x"0b98719e7f949c1a", x"7ad382e654524a44", x"51868476bfebd501", x"5d0e53792325785f", x"3a49b8ea74ba0d7b", x"4c77ee363c6b2f87", x"9d39493c7a12359a", x"a49efca1d0d645e6");
            when 27948630 => data <= (x"9a962531b2707832", x"dba7ab250aca49be", x"9a62686622e43582", x"eb0fd92b197b046f", x"6fe58bf4d9ed19ce", x"40e11d21aa357d20", x"83c61d9b310830da", x"2a3174cd85636173");
            when 31306963 => data <= (x"5a0517971d4ce73d", x"33de8f262a700175", x"ee78a5fb25b4c427", x"9cea803ec61fc4ff", x"3473d478988999e9", x"09029d1d36cd903c", x"faaff0364601eb9a", x"f4be415b4662125b");
            when 8250718 => data <= (x"b105960c38f080e4", x"5767571507c99199", x"6f41c2824f3c6b93", x"1864d4bacc2c71b9", x"3da3ca7663741cf6", x"123866d8d21745e5", x"e74336fee96f3b77", x"dde57c78c05b5ae3");
            when 13163249 => data <= (x"1d24b6b606021d4f", x"bbf749c5bc9ecf37", x"edb46e77031e0d19", x"197404128f32ffcd", x"eb6b6a563cf77576", x"063fa544a442e101", x"90e3d24f669f8c32", x"1926e67174468b26");
            when 31422050 => data <= (x"a0242b241dc8e88e", x"94946258f6194fc1", x"09b0d9ce4677c148", x"3c39ba2dafed7fcd", x"249bfc2aa9782c6a", x"58073ca8198bd0bc", x"851ef176d6bdd2d8", x"c6b5af65a63ff420");
            when 31750590 => data <= (x"917aa19ab7177c3c", x"133d2f264fff5748", x"77bea427c3f747dc", x"5bd3fac4ca30e6e2", x"8825012b576dadcf", x"82109a4558a3aed0", x"206c0a6735da054f", x"70b79fbc9298cc63");
            when 27212296 => data <= (x"95a6c5631c470ba2", x"a14c1027dc57e321", x"bf26ad85c624f5c9", x"3b28c77961942c74", x"4510326e191a8066", x"4d26d5131cab4d11", x"f026bc73877fb12d", x"788c1b34d2047c77");
            when 7039234 => data <= (x"b99334ff4d4d6a97", x"e3e115f546a7d2f5", x"35acceb79220110a", x"2e3b1aaede7dda4d", x"ccc68293b90d5a5d", x"6dff26082a66714e", x"477357e8425218f4", x"6e99ac3b8d71f5d7");
            when 25950347 => data <= (x"f8c1f2b76126dded", x"deb55ac25aed6b09", x"02390e44367c89a7", x"c9cfd61118810d2a", x"08f666bcec5f7b6c", x"f4f46c23639f9ca4", x"48e9e29962de7d7d", x"f86f20ad1bc17669");
            when 22894153 => data <= (x"38212b02b57f3fa3", x"36fc2a276cdeed65", x"8971daffa117f61f", x"91d147af7d489bfa", x"6860af80f2e3c7ed", x"d929d0ea629b219d", x"a2e12858dd8ebad6", x"69c32a9032273bed");
            when 10678784 => data <= (x"a2201aab9c463b6d", x"bdf3a854484dee68", x"f3e3132a5503760c", x"4a6692d80b1e41ab", x"884effad57f31433", x"eac7dd1f01818843", x"3af06339a0357178", x"14fc9a20df81921c");
            when 2013693 => data <= (x"97ed3d303172500f", x"3581ecef75ca7f64", x"febd2f3b2d2376ef", x"678b882104103495", x"2ebb026cddb5c907", x"1627dfcdf7cdbbf3", x"7599d1190d881eee", x"2db9123b7510e69a");
            when 23919881 => data <= (x"8d9dfe4e6c17d411", x"4d19b017c1d1d1fa", x"45109084d364eb1a", x"4388104cc4ded910", x"7d911d87e2752a4b", x"6ca1027c82b15a36", x"56872262ab6be59c", x"63f1848fdb2cde32");
            when 5718403 => data <= (x"d45468da29adca4b", x"66e0b10cf3891d1e", x"e146718868e7b8da", x"3a72682fb94a453a", x"2ad89d9051b97db7", x"6281919446ff70e1", x"d1fe7d38837d2eeb", x"e7c7215d29b3081e");
            when 20384326 => data <= (x"b4cbaef1941d8ec2", x"4952d51f8e4cfc35", x"6eeaab3aa3fc0b0e", x"92fcd7d1b7d4aa44", x"e48fabd0b7824c03", x"3969b53199df1b9e", x"f2af1dbfe00c87a2", x"c7c71fa36ae89600");
            when 21071330 => data <= (x"ebbea31e6b4609e1", x"c2a3b449b35e0591", x"2acfef0ca8e42123", x"29891afc377d7619", x"ef6231d712781b26", x"b61d8d17416b561b", x"273581e3cf45bf5c", x"a162e03dea177a33");
            when 18270932 => data <= (x"2b188a91fcc24a30", x"cbed2915dfcda5b0", x"17a00d90aa329451", x"4b48c046a28bbfbc", x"4beaf54637a4a71f", x"49d619b1153ede7f", x"321422522ba5f088", x"a6a1db88a445cb8f");
            when 31060027 => data <= (x"eb01b04eec7b69aa", x"5592511cb16124ed", x"21e4c2645013e298", x"3f55fe855c5a7a09", x"ccd48ddf9b954f86", x"9b387677432700d5", x"f61baf224f304e65", x"17a13635dc361629");
            when 21085015 => data <= (x"7a5aaad333cba107", x"5fff801e8220046e", x"95fdc900c29bf2d5", x"74106dc251298d59", x"bfbc278c85e7db1c", x"f818b7ec04f9fe7a", x"114712782b46cb9b", x"bb04d7c48615d87e");
            when 3493840 => data <= (x"c88a7ae57d466e11", x"b36905ba2d440ddc", x"7e66aeb2f6ec95f0", x"a385b55bcf5203c8", x"660cd21dc2e5df83", x"bf092a06d0c10e91", x"a2a290646df49750", x"04591c9928166510");
            when 31136408 => data <= (x"636fefb453e2f138", x"b67828902434304d", x"8d3d51bddb164f3c", x"ae1ebd1607f073f1", x"a5ed471f86cde82a", x"6bd165d532014d75", x"b44616bbbc6aba68", x"7bcf8e5617f1ece6");
            when 19151433 => data <= (x"ccd1af711efbc7c0", x"c338a2643b640632", x"928f6253e940420f", x"47ee3c5f78b605ac", x"cb39df64cba72f5c", x"7a9558f8b89cb69e", x"e470ab5c0b973b4b", x"4394b0143a018803");
            when 9365454 => data <= (x"8f72922e9cee01fb", x"036a16b40a07bd3f", x"2144bbc67209167e", x"557f82313a9ae3df", x"d8db3f8459e19b86", x"2e0054c476b4bf84", x"13432671db3bbfa6", x"94523dc039937e26");
            when 22355375 => data <= (x"40f25ff5a99a9e68", x"70d2c6b8571ca316", x"4d6d7d31298d5f2c", x"8add80cc3f4b6a66", x"52c7a96baf5951e5", x"abe0771d04629b1c", x"2cb4418b6eeba569", x"33bc1eea52e875ba");
            when 33899998 => data <= (x"d894576a5b28c82c", x"4d9f010947fc251b", x"d93827d4b2d5a198", x"ea2454797f9a6792", x"b214a70c93598e74", x"57a7ab04231fc46e", x"2229492725cb0ea5", x"6eb439808580753d");
            when 30754149 => data <= (x"30a2a47504c4be7e", x"5b97ec4c9e97963b", x"f0feddde183c093f", x"e285ed395ffdfce8", x"6ec31b7830abdc44", x"0d8aee2336f2500f", x"9cac09c7b2a9244f", x"bcef48cbe7d301ca");
            when 26545084 => data <= (x"28bf61a8daa3a8b0", x"859b919f51537e1a", x"5844e0a92a4c1d49", x"6aa68889815170e6", x"4542dacf4336492f", x"ecba89106eb3d41a", x"74978b3c7071ea51", x"84cdb36d18ccf013");
            when 18038242 => data <= (x"696f71fce0f69861", x"f817a05c0e9a3a0c", x"3e7a7947ee2b9e01", x"d4e6bd79aebb3c81", x"e5f0f195e23c9136", x"4bc256fe2bdbe835", x"5b4aa36a96bc01a2", x"d51766ef594ee16d");
            when 4349163 => data <= (x"96a778699577958f", x"63e506b0ba42ec96", x"ba2df2f0dd72c7ab", x"b2f54163a4d80b06", x"9ff11a011b8ba343", x"dc0acab25122ad10", x"77d68a4a014edd93", x"bc170428525060a3");
            when 12046900 => data <= (x"3dd479f7281778c2", x"a5489711503c62b2", x"df553fc68f3b87c8", x"b64b72f67acacb71", x"87945a0a36c6f0f4", x"5bd1a2d196a1380a", x"d44d5bd87c0d5265", x"45ab333413e9cdb4");
            when 3060291 => data <= (x"08cdf0ab60fa4b4d", x"1f2553c490d3577a", x"d302c78edc3f2523", x"5127abb50eb9af9e", x"7131e56311b8b903", x"0d47f79030c43879", x"e8b31bd235f2347f", x"0d795b4ed860e389");
            when 16839956 => data <= (x"0cd44573d7c4dca2", x"df79c04b06525300", x"6caf07499676691b", x"f059c3042e7d5ed1", x"73a182005659425d", x"19bcccb4032ac5a5", x"2ed789b489dd9b8e", x"6bd284c49c32e949");
            when 4907561 => data <= (x"051ac4ce6cb469ac", x"d160e2ed39493e14", x"c8b8548012bc26e5", x"9adea6439b7b105e", x"508e96d8db3542bd", x"71efb3729eaa855f", x"113068fc9b41b857", x"2add0aeb65bb1d7a");
            when 20294002 => data <= (x"41e8e75bc96c4d3c", x"7a40d929d1b98038", x"dc9d1aa0d5ad59c3", x"88aaeddf978077b3", x"423d311e7cb291b9", x"5288aafd38699e42", x"378f32b91976cf20", x"320ceb237404e7ee");
            when 6591888 => data <= (x"68de8339b0ebe98c", x"3c12fa822b772e28", x"ce18d0860c0c5504", x"e67f9d20f31276e0", x"2ab4eab7400b57e9", x"a6d39a79e52ef2b6", x"ae0bb9d97d2eed46", x"9eaa6fb54db62ac9");
            when 19307477 => data <= (x"2aa9061bf22f129e", x"2da8e10486319ad7", x"930e696b5730a001", x"53e2f7d449e818e4", x"53cd822304ab10a8", x"e7991b838162c019", x"eba8be4eeeca8184", x"f8f209da09ef2943");
            when 8942867 => data <= (x"4110be452ac17cb9", x"3597fde8eb3b1e3d", x"b1806f3f55701a23", x"8aae0bd19074d1bc", x"913d997872727636", x"b1ca05ef75be0f41", x"df09b1fc1b908729", x"58e09eb86601b58a");
            when 27727414 => data <= (x"614d8708c7b681d7", x"2ae8c07eea97c0f5", x"c4349fdb7dfb55ec", x"14738a9b3c28b0b2", x"24edfac372d30c51", x"ed2eb2b22ce941ad", x"ff6a83d82a593baa", x"fb3595c6d284449a");
            when 23577562 => data <= (x"f359c863be2c1023", x"64a0f2524b59cae9", x"65977c16269b5495", x"a0b63a2c4bbdf4be", x"176688c66dedc12c", x"d0749d069c00aa19", x"e5e09c6566b362ac", x"31ecc06bb33c2b5e");
            when 9188285 => data <= (x"c0d22fbea644cfbe", x"87e23a834579c1ae", x"261eb5ab18b4813f", x"fb3c7e30492825b4", x"efed38d10e7b2d7d", x"c6edb873f7730b31", x"5047a526f167ec13", x"4cf6aa3b0630d008");
            when 3785465 => data <= (x"c762eda8e151b7c5", x"eafc00accb88c746", x"7ffa6962f66aecf4", x"30cc8c1216329ec4", x"4e3f46533ccc48d7", x"515f51e8a4c22367", x"72176e7d998f0b3b", x"14d3274adaa121c9");
            when 32063298 => data <= (x"738265ef1b1e01f1", x"98ce779d865ad401", x"8db9abb738d21b67", x"53cd0eac5d8bc225", x"d9c4694019be76c2", x"509a22e0cb466094", x"146f27a5b731b738", x"db7d100afd4a3f8b");
            when 17873822 => data <= (x"9583dbaa9fe57aee", x"031600c1ab181d9e", x"c8e4a00fb4fe79cf", x"372afe737b8b417a", x"a32042d7d88783cb", x"35ec8d8e888d225a", x"98130330990ccd48", x"3975adf08808458b");
            when 7965479 => data <= (x"cdfc93df66e1de1e", x"037905f078507325", x"b0de95f5829a100f", x"3cf62259fce1692e", x"18384dc365bdaf94", x"b9c9b213d48ec7ff", x"39269680f2af41b9", x"960b6921396d56f1");
            when 5183735 => data <= (x"7b3fa90b8114521a", x"028357d4b5b62aac", x"be27c8106da0f15b", x"f570aaa0b030b467", x"d148a9bcdaffd713", x"4da8574611439271", x"b95497099008452f", x"5afedfb0ee7f5945");
            when 11896464 => data <= (x"0eb0a6e490e2323b", x"4a766ca9a988d3cc", x"b87087b88ecc4d90", x"51aaa534be528cd1", x"acf83b7c765d9c38", x"c7ba6d2ef63ca8a3", x"62305935e986f9ff", x"28578917234ddd72");
            when 30496708 => data <= (x"4acfd13e8c6980c1", x"6e9a90aa918f1928", x"5166d62270287182", x"1b7b045b7461e253", x"200edd20081f5df8", x"4c94c86cc7c295f4", x"f5e357019deada2c", x"cf0a5800bf27b344");
            when 25407473 => data <= (x"2bf93dfef1950bef", x"97b9e5adb36df1e3", x"70b898e5306810ea", x"2d7fa43e2352ef1f", x"69677ffda1b31227", x"d095a0e9ca78474c", x"3a07754703967e83", x"d66524b37d7b5c3c");
            when 31595360 => data <= (x"ded22b18c1068128", x"28718edc2a15ca77", x"dbadf72dc0c8541a", x"ecc5a16a68a84fe1", x"674d297d173dab14", x"e8fad043a8ca737e", x"c85c8060dcade94b", x"e64dd39c40209d9b");
            when 23851464 => data <= (x"49e2839665889b4e", x"a8ec686a736d05dd", x"8ce5af0d4fec0705", x"1109204857cd0614", x"9291561052c9b64e", x"e23d4a42d6a2ae80", x"dfc39f3a300c5ad1", x"5b0fdb48906ee418");
            when 17194305 => data <= (x"cf8103bf1c0223b5", x"bf16f58e91c49380", x"bf9c67dd6746632f", x"b3c1c4fd9b58ef4a", x"e1397da658b9d378", x"4c0b364fc37b0fb3", x"a1cfdc504ed5b3ae", x"8e12a43cde2308ed");
            when 26568472 => data <= (x"8208b6495d72f325", x"26f82a2c44b52472", x"e0f5137df12f46da", x"7d9552a07d2d4d7e", x"7e862ae2b6aad253", x"49642a496648c9fa", x"05ac92d92d7d4959", x"f284c83f9ad5efcb");
            when 30195756 => data <= (x"90798899b476d8cf", x"0f8e6c1a78ffd3a4", x"c7bb1f2a4a45b603", x"60475216483c757e", x"4959d4cc15c71d59", x"6668b77b6e193e3d", x"2248a223d5fa5671", x"dfe29de35f2e956c");
            when 9140037 => data <= (x"3dcf4cb0e54080a1", x"1ebe7e53bb922a71", x"0b7551e039d2d110", x"c847f593f9b8e925", x"1a2ece23f88b73f0", x"7514992844a3c9a8", x"9afe542e7716f084", x"30d223516257df27");
            when 7046755 => data <= (x"67da7d7f3934d2f0", x"814b767a3c8de006", x"7e416e177e2b2cd6", x"5d840044376ef636", x"735943802145bc11", x"cf32da6f18cad018", x"80bd771a20d6f976", x"c2ac5145be1631f6");
            when 31174753 => data <= (x"8d72163d9952d170", x"969f13c1d936de6c", x"b073aa7417f50d29", x"bfdbd960dc9110d5", x"e1e5dfa70bdf48f4", x"ea3158392e8f6aaa", x"ad17fb3e778e4402", x"267e186fd75b9526");
            when 23229982 => data <= (x"fa5bd7849b7719db", x"835a9baefa57635c", x"5001a5983c6aaa4f", x"9312b8ec8dde63f1", x"a8d7fd8681a03788", x"6fe23ee234493660", x"359539b3d93bab79", x"075febe90c9050eb");
            when 22758903 => data <= (x"84509de0af03793b", x"4a528e659cb98ae3", x"393b2c7367a6b7dc", x"d2d604008cf7bf9c", x"2873676c8881d7ca", x"ee3d723e4a9b77fc", x"3a3323237d7ba973", x"d965d5472f13f2d2");
            when 15626555 => data <= (x"e33a7f3085830c2b", x"5bec0574324507ee", x"f15b91c03945dc1b", x"b88676338040c82f", x"edd09938f61605c2", x"ba5f58fdf585ccda", x"835e8c58fa96dea0", x"9dd2d333a3cac0b6");
            when 10764964 => data <= (x"84d03429bfde8dfb", x"2e975ef560c9b7e3", x"3b4410801a012094", x"0ff0932468bd70c8", x"05c182ad0ef9dd48", x"009d66219aa0ceb7", x"c232e654a6489877", x"e45b8adce5650313");
            when 13398189 => data <= (x"2b8e58707e1dde4c", x"0823cc1f776674ac", x"930e50516862f993", x"f8aee760831bbba0", x"5db835c8cb3f8827", x"90238009dffc9c89", x"7738973ef2b9bb4e", x"4592da6672f1bf1e");
            when 2350503 => data <= (x"ae9046bcb6637a27", x"27d675696a14900b", x"087108345f189784", x"142cf4074c01f445", x"241a2f24734d8dd7", x"9571fe2f8eba60c5", x"c2cb7b0c0c455210", x"154e2b7a70502003");
            when 25295514 => data <= (x"dc9889697c1456d9", x"24a9234dc0e92cfb", x"e483d97da10ca989", x"24503adc775cdd72", x"997a66d2aa3d6ad5", x"532836cbe8f846e9", x"3318aa9d33423136", x"4d6d2af796949636");
            when 15433315 => data <= (x"8de7609329b2e505", x"5f7431f903840633", x"9ee41222727aaa8e", x"b096a0ca85cd7580", x"4e891afd7ac06dc5", x"74704b4033b8f570", x"33fe216ff96ad680", x"17219d19d1d74384");
            when 14333313 => data <= (x"2c2521ce3600026e", x"bb9361d2795ff3d5", x"4690fce74d786d33", x"c900e4ca86384321", x"a044ba08c3d47881", x"593c1c65a4e2cd06", x"7261aee2fee04635", x"335dcb01ff1450c7");
            when 29838298 => data <= (x"9e57e57293f0b67a", x"ae08aaf9a4a32833", x"287baeeae119f7b9", x"c9c662ff42ea8fbe", x"6f0319e9ad97ad8a", x"855674a1d80615a7", x"90ac5eae7b8cc9e1", x"b5aec9f1e4bad077");
            when 24414997 => data <= (x"e2ca4100bba8411b", x"4af0c6b0e5cf3079", x"e46b997971c00fbe", x"5c2f9fd92c92465b", x"b9046fc2409bb15d", x"da56a06db88499cd", x"c24ddac59a04efe2", x"e935ba836af1693a");
            when 23097857 => data <= (x"56a72d1062d91520", x"6003f8b96a578782", x"863024632bd16b05", x"82e37a6800ad3732", x"d3ce1764e0cdfca3", x"657878f2758e246c", x"d3ce152fa309396e", x"2ed10f2818988375");
            when 3154062 => data <= (x"29a7989d253f32c7", x"6c27939c6032f4b4", x"e98061fc21e2c288", x"bf7ba381fb8b279c", x"f231a8ab6869a856", x"3b155cda1eafe681", x"014d2595fbe15b10", x"20e6d0b2ac400eaf");
            when 11416690 => data <= (x"9e4b058c45680902", x"f073d2828be8b787", x"f94cc33d86fc2284", x"a8441a477596798f", x"90fd018211e2f366", x"7b212c1eeb01d207", x"c5729a74792c3e95", x"c461c37c1153900d");
            when 6428273 => data <= (x"fd18459a3170e7fd", x"8de4f59516b61030", x"c58d44e09bd8f999", x"fef41b89e2ab9628", x"586761e719382dfb", x"eb148b155f88442b", x"0af1c12e7e76f506", x"6ee2a22df7c06778");
            when 29158933 => data <= (x"b0ed91b40591e161", x"d517a76bf4085c87", x"cbba9b147e82c57f", x"cc8716a3fea71ff7", x"c139c084fcbde96d", x"3ac0f3c2a7d4c967", x"fa0b4742dbb237e1", x"5504633ecf1932ec");
            when 20886618 => data <= (x"7caf6f0d53097e2a", x"17acf77e0793060e", x"27c5cca810519430", x"51c20dd65caa5cfe", x"74010bcc0c6bf49b", x"ebfe53d7199f8809", x"7b043d32d3676d5d", x"d0df3e209d5793a5");
            when 16586634 => data <= (x"f6a800ff691364a6", x"19b05fbedd23bab0", x"6f2507020cc6631c", x"7a9734e1a01fae85", x"878e005cf4b3523f", x"a50e48051d14d502", x"81c1da20f1207f32", x"383586249476281a");
            when 9975679 => data <= (x"c5738f8837775ab1", x"26052767341ff7b8", x"8825c30784843d1e", x"458d06dda98e64b0", x"275afdab32bcbe20", x"9f08362a1c970d70", x"2c139e2bbb883a71", x"1e891cfc3c5a8af9");
            when 16501306 => data <= (x"eaf7d997edb616c8", x"08a2d092cb2fbae5", x"eaf4ad276032c1df", x"b485af09ea925f7c", x"824a8731739ab1b9", x"81cd0580340a105d", x"dbda0c8def51aa64", x"04ab1bf0bd2472cb");
            when 33071548 => data <= (x"5cbb9d59af7ea02a", x"20e34c47be19f732", x"df549b9c02e8fcbf", x"580f6419e8e7b86c", x"ad91aa418debe32f", x"796ddf9686ec8978", x"c45ab72f10a47a5f", x"953f0acc27c149c0");
            when 22358189 => data <= (x"3ef437cc0ddb15c5", x"4a713b24d3bf40b5", x"30c5631ec49120e4", x"3267e37d84ec9ce6", x"0bcb8bcb701ad906", x"312a7af205be8652", x"ac412bd7cbf5c6d6", x"30a43dced7954177");
            when 5833231 => data <= (x"458b37d454161034", x"4ab17c566514b825", x"123a4ce677445473", x"9f43dfcbc0da4d27", x"2f1ae4caf01d3183", x"06530c442e61eb8d", x"9be9953262c6f00e", x"398900afe2e6197d");
            when 16075993 => data <= (x"419305e1429e273d", x"9b2d2c47d60b114c", x"b6abdf77806189b3", x"b4e3c6d37188045e", x"2bf3fae8d1c3ecc5", x"369c9a5ec4681392", x"c8f881943fa941e6", x"bb4950a9f43e054c");
            when 22648643 => data <= (x"b16e96dcb1e4e8fd", x"d462fe55ef167393", x"1a4ff0448f898c7b", x"90d965c5c99b9435", x"d985fbfdc035aff6", x"eeca7afadc60e7eb", x"877418084fc57d94", x"b8a958a3ed651bd9");
            when 17393561 => data <= (x"7050c53b3c7a515a", x"2b35718dc952f25b", x"f0ae0cfb308f4b4b", x"115516de83683397", x"e07f927269824a7d", x"b08e399ff92131ac", x"bf57c2d775ef2176", x"12c5c3025a044cad");
            when 15070214 => data <= (x"90330a90afd6eeea", x"a3225614430d0dde", x"a2b1d94b38c92fd1", x"6d6749c22c0bb0aa", x"790436c089430a84", x"58c3af0d8dbb1704", x"3926ec10e672e387", x"116671dc6310256d");
            when 2323787 => data <= (x"a0d8e307d37847e8", x"ca73e9ea02ebc8a4", x"30a801619c34221b", x"c3ada05323165754", x"1cbdfed66bd09690", x"91218c43b216f118", x"efc4b66e96220432", x"e2f242bbf4dbc34c");
            when 26438177 => data <= (x"19de2533f011cb7e", x"b2eb7337a1411747", x"2e0ab7eb0f951ef9", x"22687aec5c6b6bfa", x"4fd69b791cc75fdd", x"59a1d31e9d19546f", x"8b5da015625f2dd9", x"3859bafee9a77cdc");
            when 31189163 => data <= (x"91f4495b9f251320", x"242b54648be52dff", x"46392e4884ec84f3", x"dff798c54e892710", x"79f85c656ea8a8ef", x"8d6b73bddb15aca8", x"6a3ea3472b99dedd", x"2749730c93111306");
            when 22557836 => data <= (x"18d73cc3a4bcac70", x"e23b5e45cd636170", x"05c33ea575dc4390", x"c2ac2542e9947e46", x"451c09ab7a20f609", x"fd8a65092816fbf0", x"efb09d0c4b1e2f3d", x"e139afc7922cd725");
            when 20510960 => data <= (x"a405d9c6a6698ee0", x"f7258645942d4dab", x"c83b306a468ec760", x"192cb096584b1333", x"dc45b50b7edbea42", x"d82874281510209b", x"e8fdb1aeeace3456", x"e0589acdd1b19a52");
            when 32401925 => data <= (x"7dda01c70f6f300a", x"02ec60e1c485e3a9", x"3d3e2756637695fc", x"9d1f76972b398f3d", x"ea1bd87e1d05d7fc", x"09cda417983f67b0", x"ddee81d0eb724c2f", x"8f1c0393530d2663");
            when 16682757 => data <= (x"aa6585df41057ea9", x"8f539d74b366d720", x"0c08b9edfd24e1bc", x"aef6332d49fa36fa", x"52fde6e0381d80cd", x"84d6a9155efbc1dd", x"082670ce2fa662ea", x"c16b768e629ad324");
            when 17126294 => data <= (x"ee51c62343a4ae05", x"079784eb826006c1", x"5d02ecd9d3af0161", x"47b268298ba17006", x"036e3280e9c50234", x"bb9c0bf95276dc66", x"061b067e8e331ec2", x"36a32dc3f7794dc4");
            when 33598623 => data <= (x"ca42cc9d6580e541", x"d55b77682cbda220", x"ea989f86a4fb270c", x"3d39b8195bbb24e8", x"b4dcfa7527adb7f5", x"5b3ba7d0c4eaa632", x"41e46d9c0a46e64b", x"dfe16ff38936ef89");
            when 4016904 => data <= (x"7228366db29a7e92", x"30be894494dcd85f", x"9d6c5cd71c969969", x"bf69bc65e6e86e43", x"014622c5b0f5a37f", x"0e86167959f1b70a", x"1887a96eb3ca31bf", x"b3028f4e53c8fc31");
            when 13281439 => data <= (x"1b6dfbb2b35e194f", x"4992546ad87217ee", x"abf6c75fef3e8479", x"288eb856cbd0c1b6", x"c1d987addacd47dc", x"3a0c46116db9367a", x"8973dab8c6ec6f01", x"e5153ab7a119c98d");
            when 11049400 => data <= (x"6ac1f7df95cc91bb", x"95996e481a4f424d", x"b08c1158d8e472d8", x"a7f4b369ac1b1220", x"93e0981b91c1aefa", x"b160bc1fe47b19b2", x"d532c04d2e4c5da9", x"c38171f0ca5fb994");
            when 23754277 => data <= (x"8222ba30aae972c7", x"9bd609b0708bfea3", x"41744ff09569f83f", x"df8a4e133e7bc483", x"931193d7c62adc62", x"1067218d0a64d343", x"8b7fd0d85d03c703", x"62e528ab6498a35b");
            when 17105387 => data <= (x"f613c95e0eea6c61", x"fd3928f29d59d8a3", x"b291a624b1f920a4", x"473b9bad2992a0e2", x"f9d3d51584fff769", x"49eb7edc276f4e60", x"9ada93d6b1cc7542", x"d8a8742480da560f");
            when 15154271 => data <= (x"2dd7edb0222e95ab", x"e82c3201af5a5f39", x"22711610cb39222b", x"6e0ced3fc8b49f9c", x"162a2c926a46e05c", x"80ed4984bdb67a1c", x"88505d1e081cbb90", x"ba55fc65a63720bf");
            when 3236147 => data <= (x"961ba05231cc7859", x"e85c18dc834a904d", x"687d048f1c537f37", x"6ad93296da444661", x"90fa47f1b2d511cb", x"bb5f12b790cbfcf2", x"6fd21398e1104ed8", x"b00d24c634642c92");
            when 11500342 => data <= (x"cfd5bf813c86f055", x"fd2fb78477161125", x"0a7f6c6633202ff4", x"1493cd4c9c5ba6e6", x"0724f84da986c3df", x"a4006d288cd23f8d", x"07bd0c3da68dd793", x"69296839446279a5");
            when 4704390 => data <= (x"805ebe8f39745a6f", x"02cc6cf2f076e855", x"01bf51f0b164f103", x"3bd720662130b38f", x"3bf5d6de4b07f9c9", x"051805d965cce9d0", x"1c16adfb9842c229", x"4952ae2039c59239");
            when 6179677 => data <= (x"08a192e550c85941", x"2539125bbca09401", x"1789c72d01668565", x"9e807b6515acdc4a", x"db65ab59e3812f87", x"d99a1b69e269930b", x"69618633e660e4b3", x"0c78a3bbfe0b8667");
            when 8801992 => data <= (x"be4ac0b862e0d198", x"d36988cbea8ebe12", x"e54648d647b98a56", x"8329335243d14668", x"ded088888c380add", x"bd04f3cf2d58e43d", x"da32b364c1ab9428", x"785aad3e5ba54e61");
            when 27530487 => data <= (x"3cdc79c5dba83c9d", x"cfc700a0afa35c5d", x"7b3c3270cf605702", x"82ba4d7a97449694", x"04d5296b650543d5", x"915febb82c2962f0", x"7fca1e0f6bbefd27", x"4e998595417da14c");
            when 22950457 => data <= (x"df11edbdb4817af7", x"568c7705abac5838", x"fbb0c7a926745e19", x"f07572191802fbc5", x"0a809dcec766aaef", x"717eaf0d385dc594", x"f08e5cb80b00fbc5", x"f4736ec63ef97438");
            when 28274704 => data <= (x"278b62f4b0abdd58", x"b8f4b4f8c751ab18", x"1b40195efb93a314", x"ea598d435cb6f948", x"8db549d9cef1b5ce", x"fdee9fce32a8c988", x"9850bafaac2c2479", x"7aab840c0a87257b");
            when 1177338 => data <= (x"9c857b03f04dd9a0", x"89ba1fda554cf6ac", x"ce3b2e4fe88f8ec0", x"20cef02d070df98a", x"6d80621563d3b2ee", x"1587c11ef745e72e", x"5f3f97c557079468", x"3939f2a4ec2e7cd0");
            when 6409668 => data <= (x"05fb0185bb499ff4", x"1b29a2bed07d288c", x"861113833a427e51", x"f6d4930b5ff1e411", x"be3acdc0d2c024b3", x"626e1832fcdbb106", x"a0516ae021a8a318", x"34a012a9116529b4");
            when 25093745 => data <= (x"9b9dbbf35c50ec42", x"c5275d4c0d5a5d86", x"c9ef86b93a6218c9", x"567b8cf1acc093e2", x"7fc3430826d5e728", x"02499fa9e8ae4a9e", x"57178f7d80b511a8", x"9de1af446a528368");
            when 2657755 => data <= (x"740ae75faedcf8da", x"ba3daaf528db8d74", x"9842c2a318ca75cb", x"f731402ee29a47d6", x"104831fdf2f3af85", x"2216eb3a0c3204a9", x"b3261e96bef63d54", x"7b29fc8fdf8ef14f");
            when 11536158 => data <= (x"815967f5b85fe9ad", x"93f6195b27d2dd67", x"7c598439810a4c13", x"539979c8ced57fbe", x"9b360ec51b5b8146", x"3b6556f0b385f0f7", x"80f915b89a836338", x"abe981505fbf0a01");
            when 12867590 => data <= (x"6ed712e6add0944a", x"8f3c7942e19d9e96", x"c4ada93e3652e4ed", x"768d1c42ef41e55e", x"754a0f74160bd063", x"b77eaf71f1e183d6", x"c3d2015057d54091", x"6ef67c3dc18d4431");
            when 27739827 => data <= (x"428b5b02bd3508ab", x"d5576b3f5d878a82", x"ec884538e6eeed78", x"0682fcdf2112f7f2", x"0cd991a6f944ab78", x"5288aad85be6e8e4", x"3818cdfbe76dd79e", x"c76729d62d1d1f14");
            when 19945596 => data <= (x"5e40bc2d78147c7f", x"9cfe8fd52b37bc73", x"8908149333834024", x"15b2f7a2ecc04240", x"f217beee1297d99a", x"60dd6cad95300787", x"79f4f2cb8c19189d", x"a598533cec3d1b08");
            when 9123717 => data <= (x"2af7799dbad7ff16", x"d1fb67da6f03f2e3", x"1b11c5a7f896ea29", x"226376fbe4b8076c", x"059c4c3938e48c8b", x"a54957bf3c4e6f9e", x"c965ad8dc94637dc", x"a9b174c41d3fe702");
            when 6930006 => data <= (x"687043977a4824c2", x"c8c0377101cdb301", x"0b3a3311f037e304", x"0cb905fa943d7cca", x"6378dabbbef9bb5a", x"3cc204ebe56b8b9e", x"745e02a177c3e24c", x"9ac47c5ff1fee66d");
            when 5902821 => data <= (x"a514fd77d146721a", x"d7591e4e21ac7a18", x"126a842e4fffe74b", x"2bb17301bcc65037", x"bebde6468fad307b", x"426648a9c2cd356e", x"5a2d008033577591", x"34d87e588e6cbec5");
            when 29216829 => data <= (x"9313c7df798b2daf", x"b05a1c7aaa886a2c", x"6c93e9b336e859a4", x"1c281f5a67e3b54f", x"737c4b16a250a9a1", x"cb472c0f332fabe2", x"7394ae1c3966c969", x"84abadea93e23eb1");
            when 23615793 => data <= (x"b8b0f1409b325ba0", x"044caef69b623ecb", x"7c91a77a40d2ad47", x"100b62ac7f64afb1", x"02910c53e46717e3", x"f657e5920087ea81", x"81264dd744c4cbf6", x"bbec116961290730");
            when 2326007 => data <= (x"b98183d8236fef83", x"275da013f32fd490", x"f9a0c0c49281527a", x"a8b154c2853e032b", x"1a3d7680a0031122", x"b42322bfe2390c4f", x"3dd54d73e1b8f7be", x"ef0bfe2a56a3d647");
            when 3265020 => data <= (x"d984434287a7a3e6", x"4640dafceeb45221", x"4143a45f41e4e445", x"03f91c85383414e1", x"0d02ebe993b130b4", x"d8b0abae0e52f1ca", x"469021842eb5ce28", x"82cebd6382e84eb7");
            when 30462239 => data <= (x"1d29143efe46933b", x"9034917f413b3d43", x"1a9f4ff0489dcc13", x"2bc7e306fc6ddda1", x"f97d5163c7de66be", x"8698f17fdf7efe36", x"a6058f61577548a7", x"4748eec35710e3a4");
            when 24699856 => data <= (x"ca3306a189deb0fa", x"2c7287d7a49149e8", x"8e96f2b84792d332", x"79b47d24e679c712", x"f550b0a3961aceca", x"aab33f213232928e", x"71900406da3177d8", x"16c2cbd64dc8b694");
            when 34066713 => data <= (x"d5945333530d5db7", x"5f5da45cbb97f75f", x"4633b1db653f8fbf", x"915f4662feb6a975", x"a9b7e16626e8aa60", x"461dc65c9ac87bcd", x"32dd5a40ebc32995", x"0bca6ee65967bbe6");
            when 26913099 => data <= (x"1057dae02d9c0067", x"ed605c42ff261732", x"dd4c5a4931a7577a", x"48299f27bfa0da4f", x"7330c56e4523fe77", x"ece8bb36c3c058cf", x"26a3800c3183d867", x"749b0016a8aa301f");
            when 16725237 => data <= (x"6a130fba9e6692dd", x"8a76c07e08e08b56", x"6d72f80aed327277", x"2dc2902c03392d66", x"62438a6e1fa44e61", x"3924ee911300d7bc", x"1f1884e56cbb2718", x"ee3bd14acb580610");
            when 3086189 => data <= (x"627add66bf889b57", x"a2f877995e4c6126", x"9057facf76e0bfa3", x"1032d8d8f09c9fc9", x"40858789f27933a8", x"e513b60d3f03652d", x"75302ffdab374be8", x"208d372a9783f24e");
            when 9704520 => data <= (x"d533e87d19427c5b", x"ead9f4ffd81095d7", x"90714f20b80c2513", x"ec4eb29f7715f25e", x"afad579ffa186fb5", x"6a329a6970cbd5fe", x"cbf778a02af58e53", x"5ab2f67e522f425d");
            when 5745119 => data <= (x"e1a434d841d86a8c", x"71acdebac8da3036", x"ae2314782a2127ae", x"525718a3a5f9a917", x"70ba85429204f573", x"433023377b881b36", x"d43ccadb6fdfdba4", x"45aaf26cf01d723e");
            when 3149163 => data <= (x"63a3ef31ca0d3bf0", x"fc583aa7581e5929", x"c40d4a26d58867c7", x"f651a9efa3000314", x"d517ccab33badf05", x"b70c5c86a99a1483", x"045cf9d796e204bf", x"7c5249597fc193c1");
            when 27064944 => data <= (x"c3c09bd9890e91fb", x"ace56ff525c8d732", x"e2cb994450b9de0d", x"4a9e82dd4194402a", x"371035f5d9ebcf33", x"2a6299365723de9a", x"e14eac03fb9e794c", x"d98afd5340b51b79");
            when 29242224 => data <= (x"34561fdae6eaeb5a", x"304a2c1d79923741", x"48a95fa9b2a6bf86", x"d3267ecaa9695233", x"ae2a5bc03b2ac254", x"0b5eebdea632491c", x"99f77bbd97f15af1", x"bfd81d661c8903c9");
            when 21636732 => data <= (x"fb734cf462556451", x"f52e63a3d3e4064a", x"c1e29ce1ff882a80", x"d4130588c8485c97", x"32c3111cb440d696", x"76c12947e2723cef", x"491b1f4bae875e1f", x"aebf733c2e385816");
            when 9544081 => data <= (x"984e18b4281bf059", x"f13905b62da19e21", x"cc8a1dc440fdfc1b", x"7245edb24daa0677", x"09aa0dc05d361fb1", x"0a20cd3dc8d52d9d", x"e65c266786b23cbc", x"00c5d4c2886537a5");
            when 1441572 => data <= (x"b57d7e15708214ae", x"9be569102dd841ad", x"57f693dbb74f19dd", x"6a1c8a22cc952f8d", x"d4f9ddac3a4ab18f", x"7adeef06a2f943a6", x"bd433bb8b18d7072", x"79d6c9ee5eabe5bf");
            when 19187914 => data <= (x"22fabc1fcda37645", x"5cd91fdc1c2bf93f", x"3a8dd493abad94c5", x"ba1091e3f58cbe15", x"a7d627f0642b5e65", x"5fee4a9a4f3aa14c", x"6f54363ad7917992", x"98e3265523d39ec6");
            when 27596807 => data <= (x"1e5b76e5f4ed0688", x"8df4b43f2790fc11", x"c5f1c1b3ea55d4a3", x"adfd707efddffe04", x"071ddfa131d34ebe", x"e56a37b710395871", x"00e57b566476c49f", x"bde70c9ebd2fea74");
            when 6940209 => data <= (x"da149924c9652e5f", x"a216b6eb386568db", x"b228deb8cb11ca4d", x"a7e79ce8d785004e", x"af2a50a09e6beb2a", x"021629dc68aaf805", x"4edc4e83f5082065", x"da963d8b012d9e1f");
            when 28196597 => data <= (x"294d83f7306f1346", x"d6eaec3cd8132615", x"3bf95461fb879b40", x"f9750730c29fcc54", x"a7f2231b101044a8", x"c7056e83b52f6204", x"05d620d881fc673f", x"afa4df27d537d688");
            when 18557983 => data <= (x"15c42149bc0103d8", x"37f73c403fcdeaf3", x"2f354c71fe29e128", x"87bd3125cadc833b", x"7164196fb4f1a9bd", x"54e1f06b37fa1aa8", x"9bb4f00166058e85", x"73633044bc88c527");
            when 1649365 => data <= (x"3880f5e728dab6c4", x"053340ece535fa8e", x"714cb9888f1edacb", x"783ac5f0719e68de", x"b896a662715ab17c", x"0908d545b8bc8408", x"6d048d99d5dc34b9", x"68b42943d4df5ace");
            when 12375310 => data <= (x"8700e0fa6c56df57", x"245509a1dd35dce8", x"c76734243bf4dd9b", x"5a1dba32b0fead32", x"84ba7ea9f2dd0bf4", x"8ff23b661f54817d", x"d3fb72f69db78f5c", x"36596fc19d14dc91");
            when 2084807 => data <= (x"b6ad3d3885f8a996", x"f18fff43dea1ac26", x"28ed1f47d70ec487", x"d206b42d3f9b1240", x"0623c4e76e8a42c4", x"333364b27bb02b3d", x"b597ca06360a7809", x"fbde702ab33f250b");
            when 6652039 => data <= (x"1171edcf5e6ada34", x"bd317944dd7e9211", x"3649398ecfd5a8e1", x"d6e4f0c13b161aa0", x"ad247d1efe51c0dc", x"791552b4e224fa32", x"cb6ac451812a3704", x"00be4ac0021288bc");
            when 2177399 => data <= (x"708bb73eff2ca205", x"5b386d2b462550cc", x"7e8736c62742daaa", x"826ccedf84acd55b", x"5d2f7dfefdcd7372", x"4b7823e24203e521", x"b75d619203cf8955", x"c8db039dc87b3b23");
            when 4521691 => data <= (x"41dc1fb478fa3b37", x"5977b41d95143cc7", x"7bf47b084c2812d9", x"4fc26db844b746f5", x"2fd44ed3988642a8", x"4303d836b0ba3e27", x"2b3d35c7565c592a", x"95ae852ccf0bade1");
            when 18451888 => data <= (x"345112d605352c26", x"556bc21c53baef52", x"e62792d76129918c", x"66018d998c74abad", x"ee58eba8ae593be7", x"a515024cbc35db02", x"2468535689b06fe0", x"673777bfe8120489");
            when 19084473 => data <= (x"4360cb4d52d704f9", x"13e2ed2089acece8", x"a18a1f3858102c8d", x"9e1c4ff32f3d6679", x"94198f64a940bd84", x"74577950ff46a9b7", x"a81727499ff7d0f9", x"c70c795517dd7502");
            when 20998991 => data <= (x"4c44bc4fe15b29f5", x"ca4e3511e1850ce3", x"c1182eb529ebc7b0", x"ead619c985e4038a", x"618b814d4760c853", x"2d1f866699adeff3", x"0113a624fb303e30", x"5511a9c5845372c6");
            when 7649510 => data <= (x"ba190fdb5ba4f5c0", x"34c8ce39247b09e0", x"ebf8e4d6d227574d", x"7ff944a298ec2f5b", x"19f071c8b4437727", x"f72ead1142834dd8", x"12319b4a1901bcfb", x"398f1a4806040479");
            when 22980156 => data <= (x"6f40f1c2b2760485", x"8db0256b9a47653a", x"50088699dbc9b9a3", x"ae52dba43673dc33", x"248480780e6976fe", x"7643208610b033e5", x"39d01fbc0cd135ae", x"6270229fac0c8c73");
            when 21974654 => data <= (x"0d6c4fe5b4d3934b", x"da416009fa4957aa", x"cd4637c3e9326004", x"c87b5fa7558a6583", x"99cd1b5014733e86", x"7973f71fb66d99e4", x"d4a8d7ab5fde5d81", x"cd75fdab412a5d75");
            when 31905320 => data <= (x"f6527d1d5bf9804b", x"7381d3a9e4d26d80", x"b315678bfac684cb", x"8cdc222e62c85f12", x"275aa6f4d9fbf57b", x"e778d992b1755609", x"15169e8a096bab32", x"75ca693c347ae3c4");
            when 27169539 => data <= (x"84577e314c99c585", x"5674950240b80bb1", x"5f56c6d7847fab25", x"f8051934cd470947", x"dc6998d60a07ca80", x"1b0edf39aa6e117b", x"e787411744ff1ac3", x"f3dcaa7805e2a620");
            when 6264176 => data <= (x"a4dfc7168ea9d1ac", x"6d54f33c8f29079a", x"e8ed9b6f5da1d658", x"ed515c729b9e2d53", x"c1e01c671166d193", x"41dd09009b8d441a", x"1e0116c7570c28a4", x"c40afcefe426235d");
            when 33787186 => data <= (x"0d432e047d3b4c70", x"6807aea308bb2596", x"af9ac88afd92eea6", x"542dd2a82215bd36", x"7db8c1bda9e4f95c", x"50d5d9799ce03e1f", x"e63ad8d0e8ae1309", x"c7d79d5c4eab248b");
            when 27656388 => data <= (x"35d26218caee73e7", x"bd1fbb4b07a580a7", x"71c06eb7a0087e4c", x"25bd2ee841f21884", x"fb6597a74a36257f", x"e511d3765680941f", x"e2362bb88338364e", x"5a9549344f4cc866");
            when 13732923 => data <= (x"ff82c04ce4eb59b6", x"29051090477ea121", x"53ae6c4a06b1a06b", x"2821dbbe87eceef9", x"4f7e1cf7e04d9690", x"122f8d676933bfe5", x"3cf8d07a8d636150", x"ab1d8f83eac367be");
            when 8284234 => data <= (x"2e79c13f8a8f534c", x"09e69da326577aea", x"42598b75238756d2", x"5eedb0ed56d829fa", x"545567adb1673036", x"e431c0a6150af8bc", x"889163a364c81fd2", x"886341657f516c47");
            when 26596016 => data <= (x"60a3031b83546b4a", x"906bd18bf1057b94", x"66f0b22542ce40f8", x"f1e798bc500af39c", x"51923afe50ed4edb", x"278658556f3e07c4", x"2d231d840558a798", x"9bd290a710e66805");
            when 5145452 => data <= (x"4001092476ee85f0", x"df27830f01dd954f", x"5e74f5b0eb35dbc4", x"a921e90cdb7f84d6", x"539606a123d5cb2c", x"a5bf198d73beb963", x"47b2dbfa39ac6ea6", x"b6848a3510e205c8");
            when 23216011 => data <= (x"2b03a47681a3d837", x"6f0271cdef6ea8a7", x"24d4abbd5fbb6d6e", x"44517b6fc914e7e4", x"00ff3f78b02b928b", x"a88e66d82ba9994f", x"ef6c51c4ad3d45b2", x"95d53a837b186a40");
            when 14946862 => data <= (x"b6d22b4eccb02522", x"90a4b5aa0e2f94aa", x"ddaeca09ac5c8420", x"944bd9dee7a2a013", x"ee61647fbd5b696b", x"73175c7f3fba4723", x"d53c1d54c8e0e432", x"a3cd04b8530602a6");
            when 7281897 => data <= (x"d9097da95ee7da52", x"23402889bd21ff4f", x"209d57a00dfa4a87", x"02fbc74fddf3c7b5", x"2e375a89757b651e", x"a5da30fd3e0c0128", x"a46bd9c03bc24039", x"776b4345d668fac9");
            when 15976395 => data <= (x"684d2e520b3e1a4e", x"a5d69eeaa82b93ec", x"0872ef4db990d81c", x"5e23f9b85ca26755", x"25300ba8bdf9fc99", x"91298e7d09dc81e2", x"7f593e12b7a2e61a", x"bcf6eb6b0722615f");
            when 10957806 => data <= (x"30d4408e6ff7b035", x"8e5b384432d64293", x"5c760b41f1989d14", x"9be75f42c39c4e0c", x"e4b1428339be6e77", x"732fc0b64efaa454", x"083af95b86f3eb2a", x"1497bccf8e41be77");
            when 7951265 => data <= (x"b6133f733a76bbb7", x"ebf8136b06b35560", x"3997aeec9c821f8c", x"b3a6dccbd7f025a1", x"177cc3788f80b912", x"badbc2a70af11439", x"d7c0dda82ff59c2c", x"2d8960c1f7745458");
            when 2043398 => data <= (x"ba6b3f01c3213302", x"c12661fc496492e8", x"8dcaa7d64e6bfea5", x"0d91e3f1637cbf55", x"01c5e0cacdde5f65", x"157b8adb2793f156", x"7514f782ad6e45bc", x"e844bb2b3bcf980d");
            when 19595129 => data <= (x"fb93ad56f7d6dddc", x"2b18066cc01abec9", x"28b0d324fdd31bf5", x"be4d8b3e1252a966", x"92bd56456440afe4", x"d757e9f1efdb9985", x"8150ef08e6d2ee88", x"f64251f88472b349");
            when 21921725 => data <= (x"b675e9788ababe86", x"baddc4df2d13216a", x"9657a876a9cb1cfa", x"0b7b6d9d07583d26", x"7e5636f4970173f8", x"46cb8d90724e413d", x"fcfab6ba3a50521e", x"3ea523f196f29b5f");
            when 9925671 => data <= (x"0bb170d42b3f3412", x"d6a2973b33058d96", x"8f8bd4ee25e0eb26", x"7a37d03a8284487a", x"8a5532869a25e1a5", x"be0daee527b27d10", x"332fb7bc92f01cce", x"2c4d0e71d2490030");
            when 16886339 => data <= (x"b045057c235d9fef", x"ca0f5357635d3598", x"d9e13d01f871f491", x"1b8c03aef69ac3e7", x"3fbbd189ccf6cccb", x"96a90df015ffcfe9", x"c6da2bbc7409b8fc", x"474deb22442a7a6b");
            when 13294291 => data <= (x"215963c1aca93578", x"97b8d6c9f37ba240", x"971c95cf194ae78d", x"d8b5cb2437feaf8b", x"ebb386a9fa31490f", x"629966a39cac9f10", x"ad273d71d7904cf5", x"be0aee79eba3a86d");
            when 10122837 => data <= (x"dc7eb06a2bd7ca71", x"1eafdf3255186c5b", x"1751946328781513", x"77521746ade4a4cc", x"86695e5cc867a9f3", x"ac6e981c52f49101", x"dc75f3e270b754fe", x"fa7c58a5f0ae3d41");
            when 31544496 => data <= (x"7f03bb3995d7c63a", x"d92f97659f6bab36", x"d64732d874ede2d4", x"581c03e2c1b78683", x"eee1ba74c7d95970", x"b4b8ecd1bcf17aec", x"3e0a989f6417fe6b", x"5703a679f5b49424");
            when 10572699 => data <= (x"a555466c3a8c0a18", x"a6fec7b67d91f04c", x"698f7f5a799c7703", x"c48d8d942dc4fae6", x"cdc34769812d8714", x"1b16134656689b3c", x"6dfe56f0db6197fb", x"55f6386fa0806bcb");
            when 11131045 => data <= (x"9cafaeeafd8b16bd", x"a05fb54cd24fa993", x"125e44345270929c", x"1812e19d8945ea1a", x"e75e7cced7dc225e", x"c431d45d0c66342e", x"4f8f5ccef22f74a6", x"b2470c80b5bbd9d6");
            when 565233 => data <= (x"b87a37bc5973bfa2", x"29d0f87abc66273e", x"d10d3120bbab8798", x"0848da65cb5d5318", x"e2403c8f25d8d739", x"2694c930ccc23885", x"1bde957035f810a1", x"30a12d1de871ed81");
            when 9648241 => data <= (x"f6aa35a8d9b71993", x"084e28d7128a8f12", x"61e4c38205bd785e", x"5be08eda2b3d5baf", x"d19a68579557e3d5", x"17180367d4d3cdd2", x"4d8f0e6bd57e483d", x"7de915cd5f5aa01c");
            when 7716345 => data <= (x"a9e516ef6eed9572", x"b6c84d85c6557add", x"9206e96dc9d3d37b", x"5bbbcb424e03a2c8", x"347a5571c9a2f263", x"5dabe25fb166a5e0", x"deee3fd0849f379e", x"22c66b80fa0b80db");
            when 13358103 => data <= (x"ed90d3c016c1cf5b", x"e5b463a434f27cfd", x"b8d05641aa284e85", x"87511a9c4da81b30", x"c79704f1a0afa10a", x"6b589e47007d911b", x"b17b32a161557934", x"72040240cf0d5d79");
            when 30738467 => data <= (x"40cae5315adf3cf5", x"93b19e4a0a1a5281", x"94af43c30ac29c35", x"5293f03e206e0ae3", x"cc2d76333470d84c", x"10d8577b95b88cd0", x"048a93eabbdf19fb", x"b45a411da98108ca");
            when 2797407 => data <= (x"b90dff7a59991b6a", x"169c82eb7edb3465", x"e240101786e1b7c2", x"ef43a732eaf45e34", x"08efddd69c61dabd", x"c584fca44c209c45", x"7cb18588a454a43c", x"0a822604de6178da");
            when 13474351 => data <= (x"05e446293635b0d5", x"fc3d6d546a4bc41f", x"b1b99d6e1e933529", x"7258983266ff2bd5", x"2efeeef9d73d9ab8", x"53b1bd49508699d4", x"9cf5843e1cc0beeb", x"838c71c0ad92f7ad");
            when 22050234 => data <= (x"481fd5c080319581", x"9ee8f6d327a94c76", x"dab8bfde218f69d1", x"ae020cb2f1bf15a2", x"412b8dc96294381c", x"1585394b48cd2919", x"5cecbb8b933c2475", x"f40446528d7495cd");
            when 11360747 => data <= (x"04ef3e0d2837a27f", x"b8fe004805b16d79", x"2ce709a60f214515", x"0fd5597f50d2d9ba", x"7487bae5406d23d6", x"7a66ecc285dfbf55", x"eadc775a2c14afd8", x"b0b0256f020658bf");
            when 23683973 => data <= (x"2fb63623b1bb4d8f", x"f7e8068fb10ae5fb", x"7104845a89110511", x"8c271ba316e861fd", x"f36e0a519024a0da", x"2169457b14e60283", x"abc29d4a7ca11dd9", x"2d3b530bd3cfdd73");
            when 1710934 => data <= (x"19fcd41939e762a7", x"b46daccf8c2d66b7", x"6d0f2cf12d2b492b", x"c8041791cd662f6f", x"7bafe78bd1eaed6e", x"b10e47e83a44f5cc", x"a114d6821884a0a5", x"07e47b572014f651");
            when 13638966 => data <= (x"5d67515f5067de37", x"db326d31a42d6bfe", x"2b83b9dbf0e5fc32", x"52038fa216e4ee2a", x"d230a5ac73bdaebe", x"8399ca11be2f8b26", x"d231ad61c0be6caf", x"b4e9091cfc34fca9");
            when 30459864 => data <= (x"cb51594be5f44c93", x"1df3c07d57b59ec0", x"5008de7dd0f710b0", x"9382e0ad20e0c9f1", x"9205d9622d2771a4", x"5cec3341ba2cbdee", x"2ae13e34000a1c64", x"472ca1f6e5d0600e");
            when 29369102 => data <= (x"c68aa381595c6312", x"62fa7a6a7a6d48ac", x"ff8a76ddbdf512f0", x"9bdb7c2ec6a50418", x"8d255e0469e8271f", x"427f5d162ff062b8", x"a8f6397efee99e8b", x"145dba4628aaa4af");
            when 15922905 => data <= (x"70a19c9a8f4fd844", x"ec827a95cd0a7eee", x"ad050c28ce96dc25", x"fd86aca1e82cd5cd", x"4ab708503b139d7e", x"2673e8d9e717a08d", x"c5573e93ecdbbc4c", x"a7dd9ed9624143fa");
            when 14034502 => data <= (x"f0339881e0ab78a2", x"b3a24b6c81db331e", x"68c65b02fa97d2c1", x"f5fa5adb9407c159", x"dc053b61187cce16", x"131a237ff6eaf286", x"f60c56a81af1e256", x"0724bdfba1a3f89a");
            when 20510818 => data <= (x"9ffc24887ddf2afd", x"a515183a531674e4", x"768a7adc7bc02651", x"6140327492532336", x"3cda83b7f01e2d1b", x"9bcd93b429d40012", x"1ceb54ffe08d8a94", x"454cab972c5fa480");
            when 14655240 => data <= (x"ee5a2d7bb4b7e4b5", x"1188c56507ca2c1a", x"609412cc511f7747", x"ef4a5632a58d84e9", x"b3828b46c352fbcb", x"30821399eb9f787c", x"474602bc4bd7dc38", x"f7cab97c6ef3c9cd");
            when 21623514 => data <= (x"ee7fbdd79ee28c35", x"1581f2093c118324", x"8929e6aa78cb4c07", x"df752a4382b3c4c1", x"84fc007983018f6f", x"e403be03fe56add8", x"235f056f39ce37ac", x"3b407f4993e85d3e");
            when 25535846 => data <= (x"9b2dc5ad4c51828d", x"0952fa1890c462d9", x"7f58411d99fd9006", x"f9fb0672fb12191a", x"8f81f2aa18ad1dfc", x"dd66600c316c8fa6", x"76002d6fa2f44a75", x"9dfefcbc37bacd6b");
            when 21494756 => data <= (x"9078681546fd79c5", x"1c7258019c80cba7", x"c8a4d2297e4246cf", x"5e327d04c97f76c6", x"3c717879f7bbf7fa", x"a98dd6746a6524dc", x"65b78d01dbab454b", x"7d416bf2b63ea92a");
            when 26352110 => data <= (x"73cbb62c565f61be", x"740122f4e1e70d27", x"34bae316d2a36049", x"495c117a28b689a1", x"80b82431c1884ce3", x"694d4b58de18125d", x"36e76db9df45148f", x"a510582ada539c61");
            when 9946123 => data <= (x"dc7634f06d6be2dd", x"475c480ef775ce3f", x"0262d0c8f2e0bbd3", x"f3d4d2d4575bf264", x"4252278a93ffe534", x"2609701601bbe6a8", x"bee37f588ddd2727", x"527c394d6b204d47");
            when 2771101 => data <= (x"e4f710a5bde02dbd", x"edc2a25167e4f06d", x"4379fdb0c0871b28", x"627a27a484489436", x"2b5bb949401f0a1b", x"4d5095acdd94765e", x"f5b10127bd80d797", x"e41fde53ca05fec6");
            when 19159664 => data <= (x"012e9e0b0c41d3ae", x"9f209e06659c5246", x"354c855b69bca366", x"67875cf84635b8dd", x"7d0bb99160974b54", x"fa03a52dbc2185ea", x"1ca88fe24834682e", x"3b643549485b4838");
            when 29747057 => data <= (x"d7e0fbc3e6c1ba00", x"572e5679cb50212f", x"681620a22e551a82", x"cb121790dceaa944", x"fa1d95b2de0fd467", x"4c4425490e64cb28", x"17ef104ab7b7d021", x"6978885a01823617");
            when 25670481 => data <= (x"59b9a2e4e78c0dec", x"65c10db78aa676a9", x"783e8410fbc56072", x"6178a3873b426b8f", x"253c9ef280bb628d", x"38e6aa94d65ffa09", x"5e3914f1f239701f", x"299cdce8735e960f");
            when 2545367 => data <= (x"42d19628f02cd14e", x"98db62e906d43904", x"abf2ab1fc7f2070b", x"5a92290b2338de15", x"cf7a972e3a8dcfbe", x"d85079fa86f49b25", x"0b35e9d78b24eb4c", x"3d65d7efafbcd263");
            when 23533040 => data <= (x"c7953a49d584ceda", x"b32fb65bce2897c3", x"c65f0ff5668583db", x"b31e1e986cf4d0f3", x"f2b2861ebb36f23b", x"ea8154fcf119045f", x"f63dd627523374ab", x"662c5b11b7b3f348");
            when 10923459 => data <= (x"461cbf80eb286713", x"722dbb1553717547", x"ab27c2b3267c5721", x"337d4824864910ca", x"6d1ad07408642336", x"91a10699c35f1f00", x"8c15d82ccc9bc53e", x"bd750be739443b96");
            when 5841203 => data <= (x"ce574f8c307125cf", x"7d71bb63df15237b", x"c7bd94f360492815", x"31bdafefd5b71f55", x"6cedbb2c27039970", x"29581e2a04926579", x"3e509d3308aed0df", x"834479e620e1b839");
            when 13724428 => data <= (x"b010c003b68f256c", x"30099c65dc71f92e", x"193b16551e68298f", x"862c70c069f75c05", x"09550053f9a6afea", x"494bff9dd3c104ad", x"3f17777e4e43d416", x"c4d4359c9659d6b6");
            when 5135677 => data <= (x"15daadaf249f8429", x"1d56165101e346d8", x"44c6bac3f83f43e4", x"5ab87942146ff49b", x"8d4e58d1cdc25170", x"207076522b1f264b", x"3a3d5a9ac54cab17", x"0a3ec6a89fdc4557");
            when 3517448 => data <= (x"90d02222cff47da2", x"72b4c52b9997fb6d", x"75ff1efa5496b3fb", x"c89ee4952e3fdb9d", x"c97e05da5180b7b8", x"35cd458621216829", x"1085c5cfb95c9d3d", x"2318b0fb345c7558");
            when 21114550 => data <= (x"dd72baeba348ea3c", x"30ab5a60e45ed5f0", x"17737ce03aef23cf", x"309658de22d53d95", x"a66ef460b603719d", x"d07c846fe89543c4", x"3e146316b70e5a83", x"1392851d4cb15a3a");
            when 32481151 => data <= (x"8438001899c116ef", x"f686c5bda4b36a86", x"8cd8abfb36070af2", x"8cf98cff4ea3c311", x"2f7e55356518bbc2", x"6bfdfdb795cd3dec", x"516f2cbe240fa5ed", x"4462c1e3cec68c67");
            when 10678544 => data <= (x"6ca548b7dccc8e4c", x"651c24c863e8cc54", x"5cb888d73b427385", x"7e1d5bc82a24a847", x"2060fa79b31b7ac3", x"d8abebb0f144c999", x"86728f4850e71f1d", x"9dded8eef7591e68");
            when 13431698 => data <= (x"69c252183c9698cb", x"04307186425f2f79", x"2c4c747acafa2f8f", x"8f3d8d2b56104e3c", x"4959b3bcd5ee4949", x"93126d842d051a52", x"9feba96110eeb276", x"c2015acbca8c683c");
            when 3603536 => data <= (x"3c7fef30f90c6074", x"316298553afda5f1", x"08e0efadf36ee0e5", x"ba2631c62b7641ea", x"2d370acb0c9f47f3", x"62b7a3a7559d7141", x"4af850a1d38b5b4a", x"aaaaad5a0a372f54");
            when 28833884 => data <= (x"4c07c99902540710", x"6e4ce64d2c8c676d", x"e4d1e3977c5279cd", x"3a41dd8e1f700a8d", x"ff7eb6750c83df65", x"4b5573eeb0375f57", x"096730008a7ea605", x"78f278239874fe2a");
            when 21155946 => data <= (x"6b503da3b6a88eab", x"ce130974fd78c72c", x"f74ac8e7bb8efab2", x"d1cd6f013f714448", x"a2962edc057680d3", x"b1a9e9a29cd6854b", x"08968f8b84a089aa", x"c29a2bb18d347c7e");
            when 18364757 => data <= (x"7f8f8f510a7af8b3", x"631daa4c9b433e17", x"06c6d93902752b2a", x"b8d35cad0aeaef7d", x"14ba90e023a099d1", x"90ce65c4e97024a9", x"b751a9df65b54413", x"e1736eec24030dce");
            when 25992649 => data <= (x"d4f43a88eb4f1556", x"23bda2aa55b347cc", x"d931d8fba591c1cd", x"d23d70e0c35537b8", x"14f4df31b832933a", x"5af7df58f9ed8413", x"770726d1e6b35f06", x"01f03eea54ec38f6");
            when 12892112 => data <= (x"fe08042bd00b85ab", x"068ca8430771e986", x"b0a1f66c3d5bdb79", x"087b99bdfd2e4bf0", x"a4c6c5d7300e8b49", x"8399a04962fe4b11", x"c7bc226addfccfa5", x"536046a4a64a1553");
            when 14778798 => data <= (x"353d87be8c23bd24", x"6d2bdbc408e18079", x"b598478f307554ea", x"d3e533e1fd34935b", x"5d6e1fa897f48020", x"ad3ccf122d2ab0da", x"d376f5af8035b385", x"8dc1ffa693a7f39b");
            when 9276035 => data <= (x"bc517d36e6c1cddb", x"04c38c8f877a344c", x"50e51696bab1a489", x"26fdfeb9c5ffb2a3", x"d9824bf0ddf333a1", x"ed740dd923fb41e6", x"e165d8b964756f80", x"dc9f5d2ebfb2c2d9");
            when 28780141 => data <= (x"d3f14126e7a52f68", x"6baba2ca6f71ced8", x"dd69b391ca3afe30", x"ffec1e87e6cbcf74", x"ad950a0d0bc0eaa5", x"b83dfc632f772391", x"5b977f5a4fb566da", x"9b586792893267d0");
            when 4527039 => data <= (x"b37ef19a182a5808", x"5805f9af9e1c6130", x"22b055e59b94a34d", x"672a452727754e34", x"53d51b8df364aa08", x"898191f3b4142b87", x"b77e5163f1a708bd", x"f1a5c39607749d54");
            when 10129055 => data <= (x"0bb9728999808e3e", x"4de1234823d0eb40", x"777e6f56347fc396", x"dcb3bf2f337fc43d", x"249ea3673a6460b1", x"ed2031e83c71d9ce", x"372a3f36618d6a8e", x"a2bf0ac7847bd80a");
            when 8304706 => data <= (x"89b7fca5c937640d", x"077c11f83b2eb023", x"e9e7efca8615d0f5", x"b395e5e3cbaf867d", x"479150f7207ea4d0", x"b7d0b2e844f1d756", x"ff834039c8091f82", x"b8b40e40e48970f7");
            when 8707945 => data <= (x"1c4adf81fbff8ac5", x"78821295231f48f5", x"0e545e0b27162a60", x"d05cab610cb8929e", x"0ffd3daea734fbd3", x"57eb93883e644d4a", x"fb0459b36665916f", x"86ec66989e585b13");
            when 27150903 => data <= (x"bee283809c94e984", x"97dfcb9dc4c328a5", x"a6748e48adb77d28", x"a08e1f62b5721a49", x"b1c3b217bf79d69c", x"be8def96a306f5b4", x"41bbce2efb083fa0", x"cdb6986a3fc2345e");
            when 9854828 => data <= (x"f46c8623cd5b83a8", x"6b83b277178600d5", x"cc0e8bbad810d01b", x"d5ccfa9444fa9fc2", x"6df110e953a9946b", x"4d79f7ad82dbf787", x"8a50dbd96d8e995d", x"13f5ccf31a5b1eb8");
            when 3433652 => data <= (x"f0833fbda4d0e246", x"01ff518125484c72", x"86a78d06abe2e77f", x"25deda86c9ed9fff", x"3e49d0fcc65767f4", x"cee755feaffeeb1f", x"f8e767def3d882d9", x"cffb9f224ce37541");
            when 20716877 => data <= (x"cbca403192aca4ee", x"6668594a20febf3b", x"766034632d90d150", x"bc78ce913aaa89b7", x"20f6aa30cd7b05db", x"a2ee41947cf01259", x"c7f68385195e6c90", x"01f5daade1a5e223");
            when 26635339 => data <= (x"8fd5e130ce19f7b7", x"4840c9b054d1a1a2", x"50d7886dc2a6b0d1", x"afece473caab4427", x"1aed9492f0d7c5d5", x"c41a226528761ea2", x"dd3d5c7a5c476d0b", x"b206a7ced047b753");
            when 22372253 => data <= (x"07ea46ea3fb4bbf2", x"fc6c6bd136f9576a", x"fdd8ae4ebdc4fe79", x"edbd41eca335461d", x"8034c1e2696171cb", x"530f1fae52506e8c", x"3b5f24a1f215873a", x"b0ad5e77a9f520d0");
            when 6940896 => data <= (x"0234beefb3358a4d", x"77fd5ff1a8dbd883", x"bae0860f579a1ae8", x"014b7caea4914468", x"ceadae60b246646d", x"e6c98ddf13a6c538", x"107b4053dc377e5c", x"04d0150dd844382f");
            when 15467149 => data <= (x"db72a30bb3f78b6f", x"4811e8655c92f2de", x"ecc9ddb948c3db16", x"46ed3c68cc05b6d6", x"2a438d1af57a1f42", x"0865d84193bc2f49", x"55bde52bd0b23246", x"f764309762411945");
            when 10325188 => data <= (x"96c90bcbdd32e0e9", x"679b2d14d8205dc5", x"3a4ccbb4a98dc594", x"5155a5d791e261d1", x"e0bbeae004ea8494", x"64fac41ff16f44ca", x"607a52bed4d6acfe", x"3c23509f3fd04322");
            when 2398061 => data <= (x"6a3fca407ff58f6e", x"9dc95a22eaaa9a66", x"9d63b139fc8ce8d0", x"b839d8275015f6d8", x"07799af04ab88c2a", x"9dae927b26ead920", x"283be8589f7cc07d", x"097a018fd329fd8d");
            when 23533325 => data <= (x"3cfc2644ff5266fc", x"272107fd3998429b", x"5aaf4ea2dc63ef45", x"0ec22dda1297b9ec", x"5cefca3eab697da8", x"05974ac3a912bd91", x"681c25507a83cd75", x"da45142d5501c40f");
            when 12579787 => data <= (x"d340e468e42042b4", x"c511c39fb353f2bd", x"fd9a1e195ae0012f", x"c9ed8891b4c97a4f", x"1b756709fd31f643", x"7b02464d2cf4343c", x"5fdeb230ef46f1e7", x"9f6f6f16a3a1b81b");
            when 23330996 => data <= (x"a69a471e2ad40baf", x"dbf7fe573c9cfafb", x"1a3f3d4067f44600", x"f23303d1701b5a57", x"2b478333f731341f", x"cd8cdef4dc1f71c1", x"cd43b484356f881b", x"3b8265f5a464a6b7");
            when 25543668 => data <= (x"c18d15c773367f93", x"fcfc73b39c38d39d", x"7f108918c5fcea22", x"640f2b8153f6bc02", x"cf3d5f6a533ef074", x"31580f03ef25f1d0", x"1d04ee53f547e5a5", x"2ed310667cbd13b8");
            when 25531749 => data <= (x"ea008f54750ad081", x"bdd928878f9579ca", x"9e8b3904f114c92d", x"20d6b65a608fe23f", x"56fa819c02269edc", x"19f07f11940848cd", x"fe224a561a74ebeb", x"4496731ce7405765");
            when 8171139 => data <= (x"5fafd0d78a8f9e35", x"9daf126625c801f2", x"6e57a0957f5ee31a", x"10addedc10d98022", x"6109485f934fd5ea", x"9dffff95e5a725b9", x"ab97221187799473", x"0b5642b1ce4a1781");
            when 25334499 => data <= (x"a4604358a8f81eb3", x"9ffea00e9b9c3e00", x"992aa641eb55fa54", x"f735da5b15f3676d", x"05ee82f51e1b9e91", x"181d252c7f50b0bd", x"bec32085dd0dd889", x"f5d1ba439ff8c3c1");
            when 27856536 => data <= (x"e7b620afe1016f04", x"eca80fc5259ff5d0", x"92d20b314b7bd7d3", x"5372c0ab292245e0", x"180074aec3bbb998", x"15d2c02c4e80ba2a", x"5ea2d45618b0e2eb", x"28c52cbc753603b4");
            when 13261657 => data <= (x"d40d188c83ee9250", x"511d28f044deee94", x"c6f21b56517afa72", x"821b0821062ee2c1", x"0ae184ab623ce0ff", x"0f49d5b8d3a2145f", x"11ad118093696b79", x"baad32168a06168c");
            when 22188544 => data <= (x"fa3015bf05039245", x"4dd82fddd29fae42", x"7ff5103baf7ce5a3", x"e8b1b9f4bdd23135", x"816ad870d1b9ac1e", x"2fc4ab0dbea53427", x"4c07d6210c4d6ad1", x"ed645469cd6ef016");
            when 6855592 => data <= (x"c76c0c7484c825b0", x"28d2146de42f7402", x"39af0d6811ecad21", x"41a4f63c76163269", x"d959feab9570fd79", x"177ef43598350436", x"875fcab7117adee6", x"78ef61f489066d5d");
            when 5551241 => data <= (x"265fbb07ee99f35f", x"ead2418b0503b6d5", x"dbe4a63502d37bea", x"9f2205ecde080a5c", x"f657719f0501ea06", x"ce9238f13bf5caee", x"90cda499f275552a", x"209a08dcffea01d5");
            when 27211109 => data <= (x"03ac0ba757a57c17", x"a53dcc31e1d31d41", x"6ebdd009b39c1a08", x"c002838123b5ff1c", x"32dd7258384a0024", x"b75c42c33e472c39", x"a90be47792a16365", x"fba836d7531e6a50");
            when 2876806 => data <= (x"f66e0b5f7f069e31", x"ca2f2128fd650eda", x"0192fb8b2666b835", x"d3923f27e9965319", x"993994f56d32c4db", x"d52c6dd10b69f587", x"8cc163e7e8741bc8", x"39d9f18bc8b7e6fc");
            when 20436097 => data <= (x"9468936fc50a969d", x"4eea5056505a242f", x"249dced77e9c9779", x"6e08d0168383aea0", x"d14f0ecdae87a932", x"d9bf6999346740ec", x"cf4b62ccef11c13d", x"6035df9d128423ea");
            when 22667328 => data <= (x"2f9d57d2a647e537", x"e23de4343916dcf3", x"a51097f010ba8a3a", x"0be2795624c09a5f", x"8c90be7e21903eba", x"1a088d89755bc952", x"ab4979c9f179ae4d", x"9dbe233c5c56e34d");
            when 27414028 => data <= (x"ee5db3c556249a22", x"c2e399067c0e1bc4", x"244251138790742a", x"8cf736ed4b9f2a66", x"e5dbd5026d38183c", x"a120f38efe6c638c", x"4045431a1bc54c26", x"e909fe2498908b49");
            when 600931 => data <= (x"9610d9e32ace6bab", x"3787ae17cd1446ad", x"bedf939dc3638cf9", x"31b40fc880eef45d", x"717c37ec10914890", x"0f07025995cf7552", x"c4d9bbabe25dfd91", x"9757993408568bea");
            when 5198461 => data <= (x"1433dd9da11bce9a", x"6a583341a2960aa8", x"84a63ff73fc93640", x"97491ff612c242f7", x"cf9ddc3c0f713551", x"5cab89ee11882f08", x"7a94e2fd4db20636", x"5e3d6712ea013ee0");
            when 5892739 => data <= (x"cea10b2be2113be8", x"19520b708e51e391", x"c19466333b418a14", x"0b9fcaf74342194e", x"32d0f31a5b042e6e", x"0281dafca34fd490", x"7b6f96419c97a38f", x"1a28a2e3f779a617");
            when 15006383 => data <= (x"141fa1967b7b4ee7", x"7a8e7117d36c844a", x"30c5ca724f4e80d0", x"984c14032e19f89b", x"8f304a1741f0e28b", x"8c39f99922bda233", x"2e70503c2ecfcc7c", x"89ee6740fdff9baf");
            when 15663267 => data <= (x"f27b5d6c1bca5e02", x"e53fec8025d5c36d", x"db6ab73bb3efd0de", x"9cc094b7548b63c0", x"213cf905a4fd6417", x"d28c602d4f4fc9a1", x"4d4fbd681ba260df", x"e61c113814e664ba");
            when 31816759 => data <= (x"d85fa8d9ca00b83e", x"6574f0872f71a3d4", x"0ddb0bc6a5f18df5", x"00639fa435c05952", x"31d47f418acfb4f2", x"c8c16d6cc7941250", x"5a435ed552dcc6f5", x"a8caf91ade46cbb7");
            when 1478532 => data <= (x"a77721f73acd5b1f", x"55e1f17831eea6b0", x"0c8a118198cc7da4", x"227de268f838e717", x"55471d2a1df82d9d", x"2a50d009e3df82c2", x"b570c8660a5c7ce5", x"de233f99b6e30d2b");
            when 2494545 => data <= (x"359314c55d76413f", x"f677b13fa4040f28", x"8ec22ef1a492973b", x"740b4eaec3b24d6e", x"41cb65d336731eb3", x"f1997738df065141", x"3a70cf808633635b", x"4a6b64e0778b202e");
            when 20390392 => data <= (x"497e4d5a16ceaf78", x"fb52ed9bae4ff234", x"a341594e8e2ec1d2", x"86f7d06414d60415", x"dec1851daa4593ec", x"f974d3982d03dff8", x"817ad32747629a78", x"72fb4c932128424d");
            when 1985973 => data <= (x"6308cbaff0c61f87", x"57923668d6079e49", x"7b6fd33558410731", x"203543769117f26c", x"27548aaa26f65653", x"b7fab18ff0f29248", x"091ad6a6d4d438c4", x"38aee6a34cb58c9f");
            when 16707420 => data <= (x"085c8cbd8b296396", x"9c0fa268ffc807c0", x"a0e6fcd3a3966787", x"f317b052ba196090", x"c7a6e8fe54900632", x"670dbea711c32949", x"c94b87ba532e5aa9", x"e98b3ed3cf3d5c3f");
            when 19471796 => data <= (x"b3edfb8b2935f143", x"4a82e145c8dca1bb", x"b7a6bf67d52fdc76", x"5aaa4b66d90629c6", x"e202895c8734646e", x"98ada5125497c961", x"62ebcbbe1223b6b3", x"ef1a1c9b39a869df");
            when 20394274 => data <= (x"925d83e123a87c46", x"5486a21418a8e3a9", x"bdd532622a5d9ea8", x"e684bae95b3ee8a3", x"0b58c91e24917a8e", x"0e696cf67b343534", x"3369345dd7ac1d52", x"1a0033f60d6edea5");
            when 14313979 => data <= (x"7080738fedc9463e", x"4674da7cc358e089", x"930e26e01cf81c93", x"189b1d3d234508e3", x"b55270c15942beeb", x"9430de041c5b307f", x"6b70454f5e820ae6", x"5b20a834be06c2f8");
            when 12495514 => data <= (x"4d13fab8ead3bbe2", x"9db01f1cb3123595", x"cceb7012c560e78e", x"68fe063ab59767b4", x"fa8a4fcf394e00e3", x"8f9e68f35d8caa89", x"15332c7b583a1252", x"1fef76938f78ff95");
            when 4677252 => data <= (x"89e9c802f5ab26c5", x"3d96f4192897167b", x"24d04750aa05b16d", x"3182ad7ea0519fff", x"bbc7702a8b923f02", x"41d7117550943df1", x"628954f0aab47eb6", x"ba88f01f5767e97f");
            when 9198150 => data <= (x"2c487a3cbc17c0da", x"cb9a0ae585524782", x"57b1c364bb736c91", x"418d34b8bcfb9217", x"17da22ada387f64b", x"7c29208238efedeb", x"77849e16f887cb28", x"a2ce2bae56018d45");
            when 29029707 => data <= (x"d4871a1b7fd55d0b", x"81b6ad67cb2a1584", x"588c64b8f98d4eb2", x"aae8476c45bbbdef", x"5028b58e28e249ea", x"83d9a1b8bfe9f966", x"c996eba114922abf", x"076799f7148afa00");
            when 28109944 => data <= (x"f9328c5fef1c5eed", x"e032dca669a4885b", x"da3f68b9d7029277", x"b623e03e5b3808df", x"014a8a83f2778c07", x"688ee86184c73395", x"ef5d9e8c2ba86609", x"8c6bd4e384871c09");
            when 3136551 => data <= (x"e55ba437a848847b", x"3383f08baf217674", x"a3772f837bdacf0a", x"8a5faab91a76f568", x"d3c46c52dbfe37fc", x"702e9b5b84d60895", x"029080a5f4d4ddcd", x"4b1b0e54db0c5f72");
            when 31923489 => data <= (x"282114b0d2ccb8b8", x"ad8108db0c33cdbf", x"f104b8b2d38dfde7", x"6fb4b4f8526bfb05", x"adef398b442e4efe", x"9ee0f3c5bf1f19ee", x"d72eac7c45f1aacc", x"380d179ba2b42380");
            when 30215252 => data <= (x"37b354843dfcc9c1", x"0a9f8c80d9a8639e", x"eb4055ad0343f30a", x"e745ca01fb1ea71f", x"f67486367fd1fe95", x"adea290a365b0d8a", x"c65a8443c46b898b", x"952c891336793988");
            when 18643720 => data <= (x"df225f699333bf8f", x"ca4e350c0a3dd1ab", x"32e9bd2f066283ec", x"fe9a7fb907751ceb", x"b4f9eef3b7783ced", x"17fda87ddf7f4d23", x"d0069b356be593bc", x"caf9ea619137a442");
            when 15112499 => data <= (x"21838191bcc9020f", x"7b8c755fd304caf4", x"706089cd6dfbf6ee", x"4684ed7b22d8eb49", x"a43c1472e3bc49d5", x"7c60d39717119e6e", x"82f725c99433f5a6", x"fdbbfb78be2b95c6");
            when 6586426 => data <= (x"233c1cca0b57df54", x"2adc933d2c11da09", x"dd6f86bc98930662", x"85cb56c3e6657888", x"652d82a17681c270", x"9eb83d966cb6a70b", x"7d7f3066ddfc946a", x"093e943d3682e652");
            when 8786704 => data <= (x"4532868a914c8790", x"8d962b415b547420", x"b1a4302a6ae3f05b", x"2a0d76b325207b6e", x"24fb6141f0be30f0", x"9ad0642a642010f5", x"cbf2aab07dd77bec", x"dc248b92aab10ca2");
            when 2422626 => data <= (x"a3bf4df084e6bb8d", x"d333537449b72cfc", x"d216a7a69e9a96f3", x"34007f03ebdc6c81", x"db0dba38f9332c74", x"512231b17b0d8620", x"50cd47a195102cee", x"141fb63083a48765");
            when 14254024 => data <= (x"98201aab94185a48", x"c23ae48e8d57f8a0", x"ed47a2d5d2092a2c", x"8692dd8367123c72", x"be670290809740c6", x"28b4902f4fb49b71", x"0764c7bc067127cd", x"9b827bba2156564e");
            when 29347273 => data <= (x"1d6929cd6c7343e8", x"542233e396f9073e", x"9c05866a23d247fe", x"e2a700e4d769f96d", x"6accf703a2dc6cd6", x"b0a77feb8983999d", x"09265ebffa702080", x"ab2ecd95b4f7ca56");
            when 26196910 => data <= (x"5f9ea2ef49c70839", x"e9756ee767920e96", x"0fcee0b37980802c", x"0c714e09f50b3bca", x"ce8e930fb544ee10", x"948d218c314e7534", x"2f882c620608fb05", x"efa599c6074c9fc9");
            when 34035294 => data <= (x"bbca97340286bd6f", x"a4f4a7a8706851f7", x"e31859f49225e4c1", x"86e8cdfe10c8936b", x"ce563e413fe86bd6", x"0523645d7c4aca5c", x"61eb498f5806d093", x"a4ce8695e28c4101");
            when 8051659 => data <= (x"14c11f99e631c047", x"f32a3e27f90725bd", x"bc23829aa004df37", x"66b435a33afd9d7d", x"f3ac9453d1a775df", x"e68743761293b40f", x"c540a53b2616e334", x"efbd9be80cb15ad9");
            when 1444621 => data <= (x"8f622b6ed5d796c8", x"178b5e984e44b11a", x"b3f8fe06e993bb0d", x"0cb4c1fb79cd4cb1", x"89706f5b079db97f", x"e582ea9cfaa05581", x"1fc68b9348b2478c", x"8a5e78b78f4c4870");
            when 14554136 => data <= (x"135e6758ae8b5285", x"95ac71ed314cdc4f", x"8cfea27237a024c1", x"978ec8104f2db8fd", x"e90c8010eb34ccf9", x"28f275fd540ff880", x"46480409afa3f530", x"ff02ae0736a5a316");
            when 2023804 => data <= (x"83c8cb36b9117a2c", x"58623e55c240868e", x"09f03a2bedd5069e", x"2f3c2682db29bbe2", x"84729fb737ece0fa", x"289bf1680565a6f4", x"7e00ae6336866885", x"f07c330cbb11cb59");
            when 15467316 => data <= (x"7d666ea797ae10cf", x"d5fc65769ece4b35", x"c901fcd49a2c08ec", x"a8719fe72d061b41", x"234035fcffba8d12", x"356212994b356849", x"17fc75338f64896e", x"8f8bfecaf94e676a");
            when 2416993 => data <= (x"48899b43e783024a", x"d2eeb575f53f3788", x"e252327b753dae45", x"616181901256e63b", x"79bde65fe5eb062a", x"9bf65104becd357c", x"8babcc1b4a769570", x"0863299a2417f453");
            when 26679715 => data <= (x"1df20681afb549d4", x"ab9a80b9256283ce", x"de8beab6e610ac7d", x"fe01425f3be0a452", x"2b7a5c26db336c8d", x"1ce787fa6fe57da4", x"09f6588a5c06fca1", x"8c976a11af707659");
            when 20343828 => data <= (x"388ce96df2f23284", x"a27b6deedc34b2c3", x"f54e0044ad8bb3cc", x"aa3dd92b23fb9da2", x"2ed9ef8c31e1d9fa", x"159dcbc2b82403b7", x"8fbbe0e73fc1ba8c", x"df159192adf9d357");
            when 12987229 => data <= (x"361e2a7f1153e3c1", x"e3172369c9524ece", x"57d5b3f81f7f15b2", x"0d90c59afea39440", x"0bdc1dc4fe01bf99", x"4b76def91a649b61", x"17c11234c0ce9839", x"8e18c8c5760ba37b");
            when 3709534 => data <= (x"3672c8cb1a47ae8a", x"74cc18560cf9736b", x"4557ebad32b8987e", x"01db88ef5d7572e1", x"8e921f6d0efe4620", x"2df40be4244993ad", x"bfe438676079a362", x"b075fab932e72d29");
            when 10272022 => data <= (x"b3b308e2ca6e0dee", x"2a1dc2669f53564a", x"63f814050318cec6", x"0f75f176607208de", x"3bbf69d79060595d", x"2e425c72770617e9", x"0a70ce8eed6caf1c", x"361226e8debafc1a");
            when 26752897 => data <= (x"4bd07396e2f06dad", x"67f8a96a7226c68e", x"c46787371c311d32", x"6b8f15f7f4fb1874", x"0bb2154868a85889", x"a65c8e7821b69fd6", x"ffcf89d6e5ded2ff", x"8283b2fbaafe9328");
            when 33177957 => data <= (x"b6ccc2666c106280", x"e338832f63b1269f", x"a8d82edd18695a8f", x"4425a0c5c0fdf258", x"56722db686860ddc", x"50014b389ed4d804", x"83b05fafc1b22ff7", x"0633566bf0c6acef");
            when 13872789 => data <= (x"f20c48a1822c0500", x"17c7eba02da34cd8", x"c296ece8b2dd313e", x"53d247d7788f1da7", x"02461da95294cbda", x"74aab3b55254283e", x"81c2ba0731674612", x"e59ec85c0c099faf");
            when 24671957 => data <= (x"8d0823066e8ed8e9", x"656b3c6cf020c737", x"30d3f681c9cdbd35", x"7c7111c0ed52e980", x"aaf66729caa0f884", x"c68f0c2a38a41cc6", x"43eacb44f7a5b53c", x"c98e0e0a030017c5");
            when 1880347 => data <= (x"6a1b748248cda527", x"77272c3730213d16", x"27527b6c400c31bd", x"da404a9cb73f2bba", x"37b02c43cf3366ff", x"6228b499586e7f60", x"e9a165142e3d2376", x"14ebb302350a29a6");
            when 16266695 => data <= (x"c83514e2aa0341e4", x"5e19fe50aa516071", x"ad8aef0e94db7d88", x"ba961fc564affe5d", x"2b132681a820e8a4", x"719178e572b22e84", x"b0ba3e5dd671a276", x"929733a2e24dfeb8");
            when 19723491 => data <= (x"ebeef58eb145c0e8", x"e9a730afc6b3ba2e", x"cb3781ff4b5216d1", x"e223d1abfd34b2b0", x"294026fa9a274dd4", x"9fa9985d96101c6c", x"7b5628c312b665a2", x"0c02512d24413586");
            when 1331893 => data <= (x"61184ab040ebfcd0", x"8da4caaae41e1f06", x"c4f6b7b14bc9b26f", x"f592ad0f7de5e958", x"8ca567349e3bfc2a", x"9dbc68ff5e52f7f2", x"55b7616087573be9", x"6ed419896d355dc6");
            when 16283471 => data <= (x"9ea2a4f92318bae7", x"e8698db15350c53f", x"cefce72dc6e2932f", x"14e623595f6baffa", x"0a68bbf51d5fa0e1", x"fe536fb192570dfe", x"68776b5b46c6f939", x"359d51e403bbadc9");
            when 28102741 => data <= (x"da2c7eb90b5ef654", x"c6bdd21172f88937", x"3cb5d04a4d5f798d", x"347426ef37c85a0a", x"d483654b4913e90d", x"69f7d7ec97156cc4", x"4c2ea77379f0a09c", x"fa1df116e3894609");
            when 32274719 => data <= (x"07b123773fa5d04e", x"4594e1aebdfac88c", x"a178caf2cdb86b23", x"1b331bf8eba99d6b", x"365e3cd5b5e0975e", x"6fb24c47052efce7", x"1273d173ef97b426", x"7e53003267449b55");
            when 19219058 => data <= (x"98865611a64a28ab", x"475f116292aa3d98", x"5590625633f73135", x"5b499c7f3139829d", x"6285299cb8cfedca", x"f3b10fb944b58867", x"01f7a8607fe0fe1c", x"c471f40ba37161e8");
            when 13607167 => data <= (x"900eb40d8f3a7a50", x"8fefe8672072f1d7", x"4b7acac76ad3afa7", x"0f2579beb6e33fea", x"2bd052342372ad56", x"ff19f807b58ef801", x"9549c7f64d0ccfd4", x"15f9dac2769037dc");
            when 7275354 => data <= (x"b02d42e5a43eb64f", x"166daa6e41be287b", x"697480e9cc921851", x"a8eb7afd7f6ee1f3", x"65ba85e78efaf170", x"e5e4c3beccef77db", x"77016fa42071c566", x"c877060e8c0f8626");
            when 5224442 => data <= (x"8de53d3149cd0c6b", x"3f9d2686f514ecb6", x"fbe0430224ca1c87", x"2ee8a1dd6594217f", x"7f409464db76ca93", x"5e3c3b88cdfc6499", x"ad35e948961073bf", x"fd2224e116334660");
            when 33890655 => data <= (x"483e4c7962a6735a", x"decc055dc511beba", x"13c103fd768f716a", x"71e43f174aa01817", x"154136fa4cac8c03", x"272e98c6b423d424", x"320a4713d0eab498", x"3b6a2175c9384638");
            when 16666072 => data <= (x"f011a7ef2ed6be62", x"62b095beb608cedd", x"f563aa4ef9960650", x"08c1fea977ebeb4e", x"0b7b1f5e8b4ca5d5", x"49b5a90b6377d2e9", x"20802f65e2779af0", x"8e38d64707b953e8");
            when 15781877 => data <= (x"2c7f2e19821e3e54", x"b9b6a5c1fb3ef9f1", x"2f40a3e39421ea71", x"ff9fd986340ac5f4", x"0939ce7c0114637d", x"6cc77561c179ec77", x"37e2385eb7083784", x"193afb78509b9bb4");
            when 12688846 => data <= (x"40e2af412a9e93cb", x"8bc63e86e0dbcad4", x"06e43f87b928e0b9", x"e41da1bac0c68678", x"707ea4fc2be2c5ec", x"701d8a7372ab763c", x"6fbe80eecd26e90d", x"32d6149f847daac0");
            when 22119636 => data <= (x"37dc76a37cf80932", x"9d8da6cdbf458017", x"2ac26af0c5f1f75e", x"97a3e9d8f9a5d898", x"a3efb92f386b7f28", x"061f3ccc8a55903e", x"4e2a185a64a3e66c", x"4de3e8e09962bbfb");
            when 33012225 => data <= (x"3615f8d45151b953", x"ac53cc9fe40095f0", x"89678dfa32396c8d", x"78e5a85fc988c063", x"61716b2ca22d5980", x"d86e24007bdfbee3", x"73b34d24baa0802a", x"27d96a6e7c11bc55");
            when 3843306 => data <= (x"de7bfab8f70c13da", x"9910e49ff2d66540", x"6ef6e432f5871abc", x"7fa3bf28e91e2358", x"e208e505a73847ab", x"6bfdb74934b2dfe9", x"d8c7a7c23e7e876b", x"774b6e63f112ea26");
            when 16344307 => data <= (x"884ce1a7af1c147f", x"96ef3331a75424d2", x"37b1e8d6cbf207aa", x"e9263996530f6482", x"bfda4640de2cc452", x"68d449478425bb89", x"e7db2ed91d81a7e7", x"c73a46b6712d3713");
            when 5387570 => data <= (x"298117878bde4473", x"b2e284f65e16fb86", x"1c19cdcd4ea94a74", x"c7d73710ca7023e7", x"3460f2b0c297d9b0", x"1f5b5f3da49200f8", x"8aa8983cc807e2a9", x"cc5458c3136b5388");
            when 25618269 => data <= (x"86f6645cf7ca8803", x"68bfb06ca1ba2f67", x"5dc7888b049b06af", x"09ff035436714832", x"53047e4a8db09ec1", x"9d2ac399d474e083", x"a11517fbf38002e2", x"c06d0e0c074e95b4");
            when 9295005 => data <= (x"22e91d96430c071e", x"3309672b1db6d18b", x"8cb695d75a8d8533", x"a81d7ca7043276ac", x"adb05f1144b3da30", x"a34b8a55fc7696b5", x"5c34a6d776575dd6", x"14f5bae3376a3394");
            when 5990745 => data <= (x"85c820f39e6876a3", x"883092e6295e3581", x"4ed10a026a2c2268", x"5b25f879ba273105", x"af8b845195a53410", x"aeba02617e71d425", x"92d80b1bb0043a8b", x"7c384368d9ae31a5");
            when 9813548 => data <= (x"213d03e03ace73b8", x"3f0cdbe60c3e7b6d", x"3b13ce5e7a950fe8", x"8754f3456ab35da4", x"617457d5e90195d4", x"6cb145ccc7cf7646", x"3dc29dfff25c2055", x"f9c7971b6d2a20f3");
            when 11310767 => data <= (x"9814b1093c920201", x"ba844edcd9d2394b", x"5cb38e3448db7d5b", x"8a8eb7d82cda4edf", x"258085dc91c7bf6c", x"967c23e9756af997", x"d420b7f5f0d3119d", x"c7eea50266468b5a");
            when 31671999 => data <= (x"10e56d5739be5731", x"547551a55ecef8ce", x"3eecb96f7cb44c89", x"186e83708643cf6e", x"3ee34ce6ef60e119", x"68d07d6035a11ced", x"5e73c567b4aff46a", x"4f4538d7d2ba46dd");
            when 32675294 => data <= (x"ba29d366ba896106", x"ed41bb09ad432305", x"bbb5e9d2f0414958", x"31604b0553954d71", x"b9ea970187321152", x"15a25237977043a4", x"7f80e6e5a9594c19", x"b089c26f200b5ab3");
            when 27954571 => data <= (x"228f7b97750b815c", x"15f5479cc6f56090", x"cf2ff8c67c02bc66", x"bb036ef9373d2db7", x"e09b0efbd91a1b14", x"dd73ef55fd71f592", x"a4388c87f784ba03", x"40c454881c2caa9a");
            when 29950951 => data <= (x"4ab3d9f16ad26c77", x"1198bd312412fb1d", x"5dcfa137bb8906ad", x"3ec0a888a6c3660b", x"9827dc324c365ccc", x"45e26df9c141a8aa", x"5462a2be07281026", x"944415d8d268ce57");
            when 24811201 => data <= (x"3f60dd734fbd0e8d", x"f8ccaa5c5af229bf", x"b2b375528aa9d1e7", x"51ca4ee395bcfd06", x"b6fd25eee0ef74c0", x"c2550488aa90d560", x"5c7e2ae1a539c628", x"42ae27fb22b283f0");
            when 5400236 => data <= (x"f72e914e44299097", x"da563654bfd16c58", x"c13f3216d06c1c30", x"34888bd6f870c1bb", x"179629642816278b", x"ff25b1c658201392", x"7960e85a9dfd331b", x"98efcdf85af4a5f1");
            when 18368535 => data <= (x"b378d655a8b9a86c", x"4b02e457e665b37d", x"1ba45c7837a75b57", x"3f1e21798dbcf1ec", x"3cb23e918d43f2b4", x"b16e7dbaf5768df2", x"9d6cf0b58be18cac", x"44bb86215f11c882");
            when 32838986 => data <= (x"afeee3a11ac70bc4", x"dc969bb633c40403", x"3131572cb6dccc61", x"104e031493e4040a", x"af9ee669bab5215f", x"bfb16ba9ea4a430e", x"5d370dbca935f401", x"6059f4141cf14ab7");
            when 28205735 => data <= (x"7695b1c8e62d3d19", x"90fdafd72fbb149a", x"ecef31db29c2be99", x"1e83b81aa3b89040", x"417b2351c4e00aae", x"a08f02725fee7c1c", x"c25e4112a53ac098", x"af91336b397f53eb");
            when 3205873 => data <= (x"1363953067419c20", x"c88652a87a6d509a", x"b8670ae260eb9e75", x"8eda86e9ef6ad34c", x"bfba4c6549be739c", x"01b732b27b55f443", x"70500047c48e423a", x"34281d0db45a5ad8");
            when 2182235 => data <= (x"375da68f2cf0e8c7", x"273459a9f8e26c14", x"121f9e65cc86b125", x"0c69f74d60bedebd", x"85c8e40f9b8c128e", x"4fd732875e17e1b9", x"c7b8f5848a4cf29f", x"d6b03091db8de73b");
            when 16494879 => data <= (x"762c34645288a67f", x"b1473f5d6514a416", x"0cc26b4754633e7c", x"71a0d26cdb75998f", x"04f4bea61d5aa1b0", x"9f66f4d3dc62980b", x"d456deb8be708aa6", x"174b10394d022cfe");
            when 24498519 => data <= (x"2e76e2681ddd5c62", x"7a885c9254e23b24", x"2279eee5138cb0d6", x"9950e64e25b11be2", x"570f1ab236cc90ce", x"e498a34a762c6d7d", x"611f299e80f72036", x"bbbad635ceba465a");
            when 8280525 => data <= (x"d91cdd30ec21438e", x"c9fae555f90af027", x"7d5f15d8c15435ae", x"4f4fd778d4037975", x"7367d0951a05bb65", x"21c5122ed9e7b1ef", x"a14ad99926f32183", x"9a8ca125ad2b0c68");
            when 17769958 => data <= (x"db7ac2fca114ae79", x"480f4a8198423504", x"4e9564136ed23e15", x"7c9a59e52b35de99", x"dbd7a265ad0efb3b", x"dd98816e196c73f2", x"207a23c3b5ba102d", x"99a09073c25d3480");
            when 15405963 => data <= (x"3cf5c0e4badf5283", x"6263b779fe1aec90", x"c0e1d1aa9f3884d1", x"65bf6f3bb49f07a0", x"50e4b0dca403aac7", x"2a0dc1f605e0b7d3", x"320c1ed36b9118e2", x"3ca44e6885cf26bf");
            when 4159610 => data <= (x"70c85596f7a856bb", x"cf79ec03c8a0f750", x"847a4ce771f76e6c", x"57f8dcca83f9080a", x"c1b8c0a279c9e2bb", x"143ce5e371120d87", x"ba44258b298e7f4e", x"9044e7a2231b64d6");
            when 30994584 => data <= (x"a0fce52c663abf52", x"dc5de189715f9e1e", x"086484e5f0219e34", x"d03571b8c503aeb7", x"4cd1c1fdee5360f1", x"676a554093177908", x"535f2a666eb6a9c2", x"a2ffe351fa580e52");
            when 32850000 => data <= (x"644fdf0a5b139741", x"0de2ba82ff610fc3", x"ef2a07781f038ed0", x"d3c408900f9488b9", x"377bf7a8006fe003", x"5521ec880bde75f8", x"75fe133613d97784", x"8ab2e14539a67345");
            when 15627544 => data <= (x"2f5a6a43b10d019d", x"cc2dcebbda8f81b6", x"0abcd3a9a8b2f056", x"025b0653a494c363", x"8f8b12e1527f98bb", x"21d58f5d286a0a42", x"d6b558acbbde0661", x"2db4d0f44c0471c0");
            when 9279688 => data <= (x"383c02f228e0c076", x"cc490cdb9bab9526", x"4d6386f6c5aa43fe", x"8910e7cbab221d65", x"da303d8b8130e40b", x"43af6a1f46fca225", x"fc708bb297ec6625", x"6aa7ba0b6ac85a8a");
            when 30777793 => data <= (x"19c99e387cf67f87", x"de206eb8cdf9f092", x"6bcd1cfc62ddb4c8", x"d656354eeea02f1e", x"5d383e8efae9843d", x"f6796b24b3d2e972", x"6570562a830c27f2", x"9f79f8467755e52d");
            when 28449047 => data <= (x"273b74223eca7ccd", x"04dc3ea10dcac72a", x"8fe7646512fdeb45", x"7348de35f9447e68", x"2542ad715c1f8832", x"1d9cc0971eefc767", x"a404b91273ddad24", x"841221b10834c107");
            when 17722436 => data <= (x"340e6bfd5c0e825f", x"b66bc2dc0b898ab0", x"7042358849225bf9", x"4e38c824f2ea36c6", x"8ec24b99d913a739", x"ff6a817919426061", x"7eea64c969c699e8", x"fdfada8816ded88a");
            when 25280811 => data <= (x"74640336f9c53f9e", x"d667473d5d27f82c", x"fc31c8f74f8c83fe", x"597676d3c2971d36", x"255cbfb4a11751a2", x"498893ce63c9c66c", x"0986421da0ec6854", x"586bf6497a76777a");
            when 7169411 => data <= (x"79a478446fb5f62c", x"44aeb11b76641621", x"c74bbdd35d0b08e6", x"59ceb260f0da0ecc", x"517736da3aef00d8", x"6cb1d21267bab917", x"636598c3b4f1c386", x"47d98371614d5134");
            when 14340549 => data <= (x"9700fbffe6cb340f", x"8690e97ef3e9bdbb", x"2461ba2a4544caf3", x"70b80c6ec8babcd9", x"36d0196c09c304d9", x"7734cce4455e854e", x"d4206f118eebc514", x"af4e433b875e23a0");
            when 31871990 => data <= (x"0bdaeaf369afb69e", x"5ce5329c4c96e8e4", x"e9e62470b114f21e", x"bb1d8222133fd7d0", x"a68c9def0b6848f2", x"631f61f5a8dbebb3", x"ea926e5c3fbe3251", x"b94bcace89c51206");
            when 17109990 => data <= (x"69d3e0ad63f48379", x"aac27172858576c8", x"3e636728a36758ed", x"8d2a4f696aa05b4f", x"5ce0b10ab0ad8d8c", x"b8a844ecda0d910b", x"9d2616e28b9f16e6", x"5ad68cc604f52426");
            when 32181499 => data <= (x"0072744389255e8d", x"c340178274af588b", x"6dcba39dfaf2f1ac", x"6ede9785ee5fa54c", x"a3243df51f6c7b35", x"537f2de672c6197f", x"0fa536ade276b7a3", x"3f10f320fa3fef36");
            when 6298318 => data <= (x"e56b236528ccbe5d", x"e1e4f3845959af7e", x"4af34a9a8a4c1334", x"1f81ecd7e5b2a339", x"683a978b06f84587", x"c5c0406561818715", x"bae761a32ca47cd1", x"1b6f0b6a534d0241");
            when 10904797 => data <= (x"d2a1bea0a113f90d", x"d2265168371127f8", x"7d7500a62459d851", x"ebf71d9d483545b7", x"f968e649cfe6f394", x"adca8fd374cff6d1", x"7b2b16b1a5f12a33", x"45c87134350ca969");
            when 6595084 => data <= (x"75942af927ceee4a", x"c846765822ec9db8", x"8805c99f1602aa56", x"aa5cad07751332d0", x"b5bbbd31e017b679", x"83ad1517a96eb023", x"62fce868d26977c7", x"603e45989ff5b6b3");
            when 5040003 => data <= (x"07ce5e4b043362c5", x"c03e404000475e02", x"ec657ddbec9e2396", x"462f1bd228b1f1b6", x"84c48fc63b9ab4c0", x"32e38f036ede2c0d", x"295bcd6c51f4e147", x"cbe10e4fbdc81c4c");
            when 3715377 => data <= (x"ddd417bdf73fd103", x"714caa760dea0e6f", x"ba6deec57488ff64", x"a033d62af4a46c61", x"9f5510b628f7f2ca", x"7827e7f42a080426", x"3286b07b9f6e65a3", x"80d9dfc113b888ee");
            when 16555412 => data <= (x"d367032077999d4a", x"37b987266656e774", x"0d1513ae33d39c06", x"8a3eeb917741d94d", x"48145bd13eeb8ee1", x"c1d72449fe126611", x"7fd779245037fa06", x"3cbad5302344fcb5");
            when 8069016 => data <= (x"dbfdd1a91c2975c9", x"7cb7f007bad1b48d", x"1bebe272c595f095", x"27a1089ac5808180", x"626586cf9ab02ab2", x"8cc6940a931319c8", x"4bddd787da42e420", x"045571cd53c19769");
            when 22356897 => data <= (x"a0bd173a4d24a68a", x"745677c00cd42aa8", x"303ee0021331889e", x"311ef7227e22b966", x"681962f83e8ad9e7", x"8c313387e1368c53", x"689282cc0b5aa58d", x"f0179df4161991a4");
            when 19633178 => data <= (x"323fb74fe3847046", x"f432e99803f8bfc8", x"076697aba728b0a8", x"138e620e20f9acb9", x"f83d42fbd2c6285f", x"1c187b4931046510", x"ce80540c769ccb42", x"931a4a603a278951");
            when 33160182 => data <= (x"29e3bc754458d1f8", x"d476fef8195baf55", x"700d49653ee16591", x"7197ea09da67265a", x"b885e7587b143af1", x"afdc8ca070ded90e", x"5d8f29d3ed9b0c34", x"4eb5731134f7c47a");
            when 4004746 => data <= (x"79bf76be14c97cd2", x"73b5c5ef783f6663", x"d3e8e07064f72d6a", x"a41c6fadefc43935", x"0dd0cd335b8ff196", x"7a79483b6f99f4bf", x"be6d59b79dbf3831", x"d843f3bb95b8cd75");
            when 15294612 => data <= (x"b9b18c93f1ef50bb", x"cb203de160d686d8", x"5c1049787435e2f0", x"2ae6eb55ff057a97", x"64e90b6ca86e0315", x"82d384efc2115281", x"be7f8a8510b45177", x"e2883bbe696346f9");
            when 27023675 => data <= (x"47c76f0c0acd09cf", x"e53f8001a2a88856", x"00bdb421489b8b6f", x"88b5d54f0b59f356", x"30400c20839e7e25", x"eb7af1ace3685784", x"f4d4b9ed61296433", x"25860a19b35ea712");
            when 28098802 => data <= (x"5e3dd414a16d2dab", x"15b80e2a5d7b22fd", x"a472ddf524af6e00", x"e0663d8599393abd", x"9f74d2e73d263987", x"804b2eb85d9bff66", x"940d9cb773824429", x"9d0f481632cbdccb");
            when 26824596 => data <= (x"f18e7f3ae1a44c09", x"300ce317b51dd639", x"db359ea1338360df", x"8867c16b44c5814d", x"7b95c793511fadd8", x"e62396b9cb752daa", x"b9b76b9f15445599", x"99f751308b3d2804");
            when 11251842 => data <= (x"86ab326ab5b476df", x"47b1b72792084682", x"f234d623a99d6234", x"e1480b4731a522fd", x"121034da5166b261", x"62580664c1d11715", x"ca40c2b89b486f20", x"a03d65432fe4d415");
            when 2933832 => data <= (x"03db59f0e0e45c1f", x"4f11bc85e3aa68ba", x"fbcd4ff3bfd253d5", x"ad441f4acc1e6e14", x"342e8ec2f6dd5b3a", x"12530cfa00f8779e", x"af8f90d8a6a75a6a", x"85bca008da6e3e58");
            when 29746023 => data <= (x"b60f4f0346ca0c09", x"3d71339e7b77313e", x"e6e4eacfa4d49cdf", x"af23d2eed399a904", x"3f8fd3426df71b70", x"4f6af6905c79bb98", x"a530f04ebf35eb39", x"b964d7bd909795d2");
            when 27478015 => data <= (x"37adce34e915b17b", x"4d0dd824d4ff868e", x"1bd09906b1f61d86", x"45eb7140a21bbb43", x"27662b5b1ecf6550", x"750c33a5c4f12491", x"10ca2d9004481124", x"4b910fd7976a7933");
            when 26119021 => data <= (x"6e84b624e9765e35", x"f73677bc99ef3ec2", x"c2278b908709a574", x"2f055c8946c3e25f", x"517f04d0e0c6ba6b", x"efde2569c7a3f43f", x"c891e31c4348e245", x"d164d57548e3c9bd");
            when 5060827 => data <= (x"45710141652a5ca4", x"54a57fe8263383f0", x"e37d0fa7f834f3cf", x"ad37e5e97c8b9ba5", x"dac13a1e8d62aff1", x"ccaaad3d0229018c", x"d3db4d8bc3e1e135", x"113773316ed507bc");
            when 6728658 => data <= (x"e43d6acbc34d46e2", x"8f3236e65ddc7929", x"04df4cc7d904360a", x"92cedf054773a7dc", x"37a14bcab32a80ff", x"461a7f7a33b98cb0", x"16f06266e36ed0a7", x"5e99326644c56a77");
            when 2781146 => data <= (x"c599f8aa2d9986cb", x"616d55f27cd46823", x"d488782bb2750375", x"7f114462f00eaf9d", x"d92b4f05e2020711", x"8155b021349fbf2a", x"7626d43b05840f83", x"14fdda4c6cc10886");
            when 4044683 => data <= (x"a75392376b96f4bd", x"bb2ba78fb3c23fe1", x"6e98768194e60d88", x"142acaadbf7a4ae2", x"aab5281ff6fe2dad", x"1b935cdc0af4fba5", x"d9fb9b55414bc47d", x"697ef569a5f224d9");
            when 814711 => data <= (x"ae7d931997b38e99", x"ff7a513c02c455fe", x"8869cdc4c8420714", x"2eccde1139c8a4e5", x"3046400d09114a7e", x"df147b085eae6639", x"c9d0b654a0eb54be", x"c455cc02bec7563e");
            when 29471863 => data <= (x"2b30946cad9b976a", x"b1bb51487ba550c1", x"2457ec80e82ef2db", x"efd0233bceb05188", x"8628f51819ef46c9", x"05d3a14da8a4d8ba", x"4fdef9e54c47834d", x"adc653a5f0e51929");
            when 24371765 => data <= (x"51fa980e3aa03548", x"bc76aeffaf45d2a2", x"89ad6bf609224aeb", x"51331d38a95ef61e", x"e442fabd05917de8", x"0e07ec91a5337d60", x"b429c2327f97c985", x"57cc345510161135");
            when 24014201 => data <= (x"48437b35ebb2584a", x"988e45f9f1938a52", x"8a5c41c4c985c799", x"bed98c5fc097d011", x"996c60d619523809", x"2b360d3fc75c4498", x"316528e4fe07f803", x"ce8840bca27960ba");
            when 29526756 => data <= (x"40c5dfa44c1b0b90", x"020a79849cf13efa", x"0c8ca8174a5dee5e", x"67d021870e33f2c8", x"495fe428e0d17d07", x"4b7add7ff674f88e", x"574d482e5669a942", x"57bb1e54c23a1d35");
            when 11035267 => data <= (x"93a7d8542247c1e4", x"140c327f89b3dfb4", x"952564a539059488", x"7b741e79044578f8", x"b2a98aae154a5f40", x"e213b1110e468571", x"f0e301101b25e231", x"d4eb364997e15c65");
            when 25510707 => data <= (x"feae30b393b73b5b", x"893f0096741af12c", x"c7158451e82723ef", x"82cb685714bf3c34", x"8b0315aa390ede83", x"6381cce39c026694", x"ca49810e07324254", x"f84d701b449c5074");
            when 9989287 => data <= (x"61f092fa9c223fe9", x"cef38220d3016cac", x"39c3eabca77051d8", x"30caa81426db0602", x"b0dc407beee73331", x"76c354505cb09d60", x"a4b8f9b50e221d94", x"1f0557b90fecf055");
            when 32648410 => data <= (x"a62a9f521fc0ad22", x"d247619b4a621e33", x"384e9e7dd55a0829", x"8ab32c23bdf08c7d", x"7ebe7aa6a6bff216", x"332e6d28476110f8", x"c53fc2b184d779b9", x"35de5a4bcd03f3f0");
            when 15915074 => data <= (x"05925c5c08303510", x"88b07e07e35825e9", x"08b6fdad3c356eff", x"3c4d317414fc0b6e", x"609bf78a732bbe00", x"e8631af414dd8314", x"4caa4e6b8bb94d58", x"3d263a6d8d106b94");
            when 2473012 => data <= (x"0d3a865cb4c3cb4f", x"65afac912434d365", x"39db155c83d031a1", x"385306f081724a5c", x"a96fa974adb322f9", x"5f45b37540a2a402", x"dca6b7bae1c8f4c3", x"c805f9255350e11a");
            when 9887040 => data <= (x"f236bfc5ed8191cf", x"2f8c3412f2ca3a9b", x"615969f53d0fe2ce", x"25501c4b41057192", x"37b0cd06d90985d9", x"b98b0c21aa84fc2a", x"34d9a2c420f1c713", x"a920aa537abc5919");
            when 33384264 => data <= (x"9d93444bfc2f59cd", x"4305090283c4e653", x"90d0941642e848f0", x"c299765c4746b582", x"4af52016935607dd", x"34ed30e15733c5c5", x"87f591ce9d2a1dcb", x"d74d08834537d50d");
            when 2841107 => data <= (x"f0d823f96e29cf55", x"1d741410d095c1a4", x"258023c4112d256e", x"8c0188cde1ad663d", x"0ccfa2c202606b6c", x"112235f2e603f985", x"317c86eb52d5d3da", x"fac3ab86eda5f072");
            when 6768594 => data <= (x"62ff9496d4d8f8c4", x"a1135575f547e7d6", x"af285aa5ae6eefdc", x"fb0981e67949787c", x"8f006e7395eb7596", x"79e445553b781a62", x"9005521e722f5f17", x"3ad284cf1af29db4");
            when 33377269 => data <= (x"a72d1c89be8ec3f5", x"cf4081a07eafd0a3", x"0ad3af99aa414719", x"f623acd42de06ed8", x"90f988af2ad3f44f", x"6bbbe48796ba18e4", x"329e0f28fc168d7b", x"abfe1f5024d21b80");
            when 6361631 => data <= (x"2e9a4d18012ae768", x"56aa358cfb87336f", x"9410300421c15adf", x"8eefb9330c871457", x"60237b8cba8289e8", x"b8c834b9f5d33154", x"c59508ef62f692b4", x"609e28c94f56afa7");
            when 15303067 => data <= (x"a7fd3c1701e1dab8", x"c21c77c5facd08b6", x"32fdeac02dda902d", x"51885367cbae6ce5", x"911956ca93572269", x"73ba47c6fa89b5bd", x"ced2e2f3ea8e77f4", x"f39dde2a348be6fd");
            when 22993855 => data <= (x"ced7119318d6de57", x"fdec3e330a05935d", x"c099f7b59e2f6296", x"2373fb1426837ed9", x"063c047c987c198c", x"77b8881500658e65", x"a5ffb9545e8ab33a", x"1de0993bdca6a5b6");
            when 28445391 => data <= (x"eff1cc9ed08e04d7", x"6c5e5fe5ec1f7121", x"d7c7611fbab8d6ac", x"a0eee71373b11f58", x"74fb2a9f909c5b62", x"5900593fc0261756", x"2bd9cf842216683b", x"cf1d123b54321c4f");
            when 27503878 => data <= (x"635887bf1b84d828", x"6ddb76fbfb58496b", x"6fd7fda615fff1e9", x"f029c8fb7ebd605b", x"cc5ac7f47df2ac64", x"827311987cbf4b80", x"36267eb51871edee", x"5ecdbe4fbe23633d");
            when 3419050 => data <= (x"89ce73f63a7802d2", x"9f178e9103384127", x"7be829a269655c56", x"0524d2600d853329", x"7eeaa75c5ea50082", x"cc5206b431609005", x"e245932bd1b87bc8", x"21988a5e8640c736");
            when 10565009 => data <= (x"878f93133fb6e094", x"e2fd683550b1b7ab", x"eb91de86871639bf", x"3421ba47a65c640f", x"9389db122d154c02", x"9ba9feee71e403d7", x"5df7c6691cb2c4c0", x"9fa6d3e5898f6ff1");
            when 33506365 => data <= (x"4d272013934fd557", x"f196ef2acd51d6ff", x"b5e5589b45f60be1", x"5ac6685755ac2b68", x"2d99281edff7d2e8", x"878fdc2782c3a07d", x"5cfdc050b589b4dc", x"b9ff2c6f7d71f73e");
            when 16610676 => data <= (x"73b23dc3a2989e16", x"507dfe254af1acc0", x"d67956318eac5c63", x"08306f63d926d9c4", x"071d9ce93af0e519", x"3fc06c278f76b8df", x"abd6eed79b8d7207", x"e91bc88060bb70e9");
            when 33915181 => data <= (x"3057446db3d938b7", x"c0e76741843af5ed", x"d8211e9448de18c1", x"df3c12069ca17499", x"399a715ba94daeec", x"fb8349445c0cadad", x"66c8605efcd5f9fa", x"a318b2bc27b0ad5c");
            when 17599954 => data <= (x"690b5c8d9b671687", x"ed31e27b54c5c7fe", x"00981076c05dcbd1", x"5ff704ded34648d5", x"11818a2aab00cb03", x"a41da5a5991955f3", x"38c663c1f9c8b99c", x"47c915406388f74d");
            when 11133732 => data <= (x"51ac5df84384ee11", x"9e5690a487268cbf", x"1372ad2a1e2a4d85", x"945b9e9953413312", x"b0c1bd534d006650", x"d5a8f377a267b97e", x"2882ddc423e8897a", x"56b45e8698a88e5f");
            when 12025063 => data <= (x"5689ecb4c06e8a5b", x"e935c5c2925702a2", x"fa36142d76e395ca", x"26a29971d80bad5f", x"fe96d057b5f727bc", x"306ef723fe023165", x"bb056d088e9e556c", x"4f591936258fedec");
            when 23888293 => data <= (x"e83ad2816a9319c7", x"986322667827a111", x"6729c9061ac4b899", x"0b506e78f5349600", x"8b411eaa59e9fc5c", x"a4a32972e0ea7567", x"2b3cf78910486089", x"a7b39d039bb28b53");
            when 7099798 => data <= (x"ec0fe49fa4ce1bbb", x"6f2cfc299a53f731", x"2f7b11d8447ebce0", x"e8c0e9dbbd621781", x"1aef7895aff88bae", x"5eea806a3523a28c", x"07b47ae3ae8303c5", x"3151013b00600fdc");
            when 5304463 => data <= (x"2f1b9dada8e5dfd4", x"a3bd21f3b2fb6bfa", x"ddbce18f5442b4ec", x"2173308b7be87c8d", x"ef8783c826e15c6e", x"21df1cc65a1a30d2", x"94f0fe8b89da8c4f", x"815625e318044767");
            when 5275180 => data <= (x"25aaf34879914fa9", x"67237473b96f64ac", x"4f49b7d41766a328", x"20f866fff83c233e", x"4b04811f1804d534", x"51b0d3a6c8628340", x"9da2acb085cbf2f2", x"46f501f99fdb278b");
            when 23375274 => data <= (x"7749c220d330bc37", x"392cc8cc7c075081", x"d12b65612d22cd3f", x"c490303aa6f351c8", x"db77c2eaecd0c626", x"64a8776232007dc5", x"010c846e03171cf9", x"bf99b87a8a78c35a");
            when 33313526 => data <= (x"9a92f2a7664ec027", x"461af20acea21d24", x"2bc4601dfc8e96b0", x"93078e7d406e64e8", x"54434316835f753d", x"07632afd66af8568", x"88aadc1e43e150ee", x"05335bd1d8168196");
            when 13656522 => data <= (x"1d10ed2a42951ca1", x"8a1dbef4cb8023d8", x"56f7cadc74c4472d", x"bac52b3903f323fb", x"0282677e7db72fb2", x"5586e26f15d08554", x"77c84dbf7960db14", x"8b77f8cb103674ac");
            when 6320721 => data <= (x"79c2881e665929de", x"4e8453ad55c2a0f0", x"c0e82aadc4bc0d34", x"b5b4cf93aa94f474", x"031bc14654a0c302", x"2f37761051c9eeda", x"a92c50243d7c7d3f", x"dd74ea10e56493af");
            when 31886797 => data <= (x"3b5fc5a3c8c2b102", x"e615cb003fe86714", x"61a553e9aa5c296c", x"77fd15928837792b", x"8d208d57ec3ae99e", x"9fad202b643f9595", x"72498714251a31c2", x"0a75a60d23acdc7c");
            when 28680228 => data <= (x"b69f94793ca4f491", x"fade26da6d252103", x"a774f8bca1c2bf4e", x"560b5cf1b283bd74", x"c0b72842cf28d8d9", x"3d6caec1dea038dc", x"612250875baea358", x"135023399e2b9d63");
            when 26568913 => data <= (x"ad3aebb0d90920e5", x"53e9f2b7fda10521", x"aec2dbe0eedd9ed3", x"4bc33d481ef97b32", x"fc30171d7d629359", x"ef2f0af00abc94bc", x"711c2097c7c9178e", x"3954cb6d7a6bd31e");
            when 22064595 => data <= (x"ebbe4c29500dfb85", x"4528f5e95de9c3bb", x"358883c30f3ed32d", x"6685eb5317c578aa", x"92b26f437666f51d", x"7b3a5232bf702950", x"3a63cc081a1a249b", x"957d5de6e93801d0");
            when 20437341 => data <= (x"3ee6f25ab7f2aeab", x"f6736934bcdc5922", x"6cbf8fb5abaf4d71", x"81a277c9593b3f37", x"6fd286993660c9ca", x"adcabbaca28db0ff", x"a9c730d659f2226d", x"213f7ff36695355d");
            when 5712628 => data <= (x"727eb11746f840bc", x"4d7948914d349bd5", x"f32ad567f11f4764", x"58e32354429cd5bb", x"83e2339984cc77bc", x"56b001728b9e1679", x"b5672b058785ed72", x"08ad23e0963ca2d2");
            when 7829906 => data <= (x"798f00ed79f13ff7", x"2a2c52a5297b839c", x"a8920baf31b1e696", x"97bb408f2ee51b2d", x"a7c9d4716155d1ed", x"f8fabb838a1511bb", x"cd0d1717006110ee", x"1cfeb48507d2133f");
            when 5079159 => data <= (x"73c502654ed2908e", x"46a4acf9b310af68", x"f981fa215209ac7b", x"b2f995b4d8398561", x"1f92869dad5227fe", x"b840d4c4097d3b9d", x"2e03929c8d16e506", x"02e06e1369821e21");
            when 18383528 => data <= (x"9c88d5f6fd0064eb", x"a899026f33a4f4e2", x"6c925c2cd770e083", x"b46c2c5ab4608578", x"4d34140b34d72f75", x"7f41460ccb1e1aa5", x"079647a238736ab7", x"c6fc17dda9604042");
            when 16165886 => data <= (x"1b8ac01a8f3b2495", x"ccf2ed79df7d9c12", x"39903efa2bff3825", x"2d1b7ea4dc387023", x"a967179c16ca7a03", x"68cea9e69562c962", x"650536b5459d686f", x"ca530ab293068574");
            when 30894208 => data <= (x"6e9071c8cf77e560", x"ff9efe23c63d66be", x"de1148295f9ecd45", x"2e27d9fa88c3b8f1", x"03b3202e83057e35", x"3c6347b488e32e36", x"542ab7027608c31e", x"2453e70d4a870a7e");
            when 31777774 => data <= (x"a0e67936e3c38e0f", x"eac39711d8971379", x"21f356523a47bdc4", x"4bef77af65da948f", x"62e90400d00a0dc3", x"01e85b79d8b78cf2", x"427570deaaa1e948", x"12e45f382ef995bd");
            when 2202680 => data <= (x"e0d01c6c2fef661f", x"1521ee2b39e32b99", x"21ae45570f22ee74", x"2414e972dfb82fe9", x"138c9ae91ffdb752", x"0b9addfac90ce7df", x"a34a0233f708e989", x"d33036f9658b4971");
            when 11180421 => data <= (x"85d7aabc3c78b5bf", x"02312d0ce36ed97b", x"cd7e1dbbe6093e91", x"3cd825910fee4bae", x"68e4fc87d991a08d", x"0eda0c2015e4b8b2", x"dbc2a695dc47ce25", x"009ab87adb9d980a");
            when 12082895 => data <= (x"bbe87faa96de5eae", x"100efa2927160b30", x"b117ba785262d073", x"5154cea9bdc8ba66", x"cb69b70aad768afd", x"55a78ddfb8c9cded", x"ad26e1aaaccfb6aa", x"474ac6c99adc02bc");
            when 12396100 => data <= (x"d9ce8556d98b38c7", x"cffe53c1bd864f9f", x"7bcc3ebbab653e95", x"8f1f14599c120518", x"3f32009c5379642a", x"ccd06e04e669a3c1", x"223c5579d36062ef", x"25f165c246ac267a");
            when 28246784 => data <= (x"3d22318f8496d13e", x"a080f9862da42b90", x"5af364f047ea54e6", x"5bf88ef587a88784", x"1c2722b29124ce96", x"257e944f34667fa1", x"9c7134be86ab1ad0", x"cf9cce2a9d700d40");
            when 16813081 => data <= (x"3bd034e6507fab60", x"410faa79623d07aa", x"46ba7df96c252fe0", x"d88a3f86ad44213c", x"f222830e87259578", x"634132931ef3b9f8", x"854f9dc16aa0df75", x"2ec22009c23e4970");
            when 21466273 => data <= (x"1ec8c13cd81bf1d4", x"4dc172368a6887ec", x"bb9389f6045ff441", x"b467ecb7352f14a0", x"0d1394b330fd9356", x"29679f4c09f1b735", x"6efc09cd464f1898", x"979a87ffb8813fa6");
            when 15124241 => data <= (x"c8150161bb645578", x"4d809f4c33c5a6c4", x"82dcc6863e18984c", x"0096a88b9c502e9e", x"04d0bc4286ef49c3", x"896b31842d072440", x"38b15212ccbcee6e", x"d8ac329ed59d757f");
            when 7816796 => data <= (x"303fb62af7988710", x"76b29265cdbd6492", x"caba76c9fa064fce", x"726b954fcafd7c2e", x"244b953a9fe82305", x"f3383a79b30d9c6c", x"000ad237c7440e25", x"718866b93923c31d");
            when 9485090 => data <= (x"5a5e10792d650d35", x"091180cb04de5ea3", x"cc9623f4f8a63232", x"3c6c491962ec5873", x"febc964a577b2352", x"7447a92304d918ca", x"32fb33252c16c8ab", x"d526706b7591b6af");
            when 9730568 => data <= (x"06e5702e2cafa91b", x"1067b00090b10a41", x"9a5ec2ef304b78f1", x"2e4e2e99d1d4d76d", x"11a9ca0ea98efb12", x"96615bfbe199e8c3", x"3d2797e6bde2bba3", x"c193545574935190");
            when 31954510 => data <= (x"ce79d7d47331c3e0", x"eea8cd9ce26f514c", x"6b88bb90c64381a6", x"eea40afc22fa067d", x"53ed80a166d6cd41", x"3d214dd42b46f72b", x"fda484ca7ea093e2", x"9255466281e0ab72");
            when 33461083 => data <= (x"98fc2965f46d55eb", x"b2ff7a4cb73f8e4d", x"43da4747c66a469d", x"4b85bf7635742f83", x"2e62fbe900d04e80", x"1017c7c0affaa434", x"42690eb5cd00c961", x"2c152a32c091878c");
            when 22407539 => data <= (x"be4d3ae5dc9264dd", x"5d57da3f06642797", x"2f0cde8cae9d49bb", x"8b69487aaa3bd887", x"ac39cc90a39dc029", x"8db59cc0bc6d78a4", x"d966ce229be1b643", x"b66db78188119b1c");
            when 32759460 => data <= (x"ff12c84e5fdd3fe0", x"d93b130e304276e3", x"cc143d6a94821572", x"77fe33a6f2045a73", x"4e5fe8ad4bd8120d", x"8cbc7ee255bee93d", x"a805f5280b3a895a", x"8dd8151140dfa0a8");
            when 21200224 => data <= (x"97c36fe8ee04e965", x"dfa44976fc3a0a2c", x"761ab8752c1d5684", x"711dcf41b8e6576e", x"2c62cd94c4928329", x"6d987a97587a82fd", x"409f2da0dea80a9b", x"639ee7d4f80d7146");
            when 7555889 => data <= (x"ac353571f8fef0ab", x"e29ce5d2d7d420f1", x"0cb72973c4f677c3", x"e984ab1dfebfefdf", x"3351573bd1dea279", x"0a9608971165115b", x"0ed4ad50d95f04b6", x"18378144897abf68");
            when 23189547 => data <= (x"d18997f2fae3a30c", x"43d3b3cbffc0344a", x"ce933c62af74cedc", x"b21b26ee68443517", x"92c5a505338f0557", x"f350020e4c3e1b5f", x"daa5ef18a85fcc54", x"7f624bf807531380");
            when 28011127 => data <= (x"9e9d61a734a4aee8", x"b7f4ba0eef287434", x"95d36a17a28da93a", x"8bca502f60251ca1", x"0dccbcc9a4aeabf9", x"b3bc06d39e80f4cc", x"7eb447381b118cbc", x"482335547c84fe7f");
            when 8544965 => data <= (x"ffb6236bf53405ad", x"db56a925fdd9b955", x"1da904a8e5d4e4e1", x"f9574ec786ad9064", x"dcfd76f947169349", x"d305c374108ed625", x"8571aa2410777ac4", x"8f50ba50bf3941fd");
            when 684596 => data <= (x"c044870829b87cb9", x"925ac806d7aa3ea8", x"a3280a562df1a062", x"7c9034731244dc36", x"42acd2d49261019a", x"3b07faa79037a51f", x"15ef2c283e591864", x"f9e775c51aeff4e7");
            when 29734537 => data <= (x"d3123bf76edbf583", x"2760a46ffe68a02c", x"e83d0a231ff60d09", x"7096fd67fb8c483a", x"b93dd4dc3599f191", x"25213dde125068e5", x"5697630d531184fe", x"7110e7cb93c548bb");
            when 31202477 => data <= (x"8ca464bee177f67f", x"11bc16d110715961", x"49e42010ddec25a4", x"6da3eb11945e78e7", x"51cfa28d1f2b47f5", x"85a68aebd36892fb", x"e463309d0db71a59", x"4efb99295569383c");
            when 31379050 => data <= (x"db50c500b4778f55", x"cb8bdec0bafcd07f", x"66d02caba94400a6", x"da38d2bbdab95b1f", x"2dbdb189629c2b66", x"3388c0b76dd76ed2", x"ca67f1f034a268a2", x"310c1cbff5227404");
            when 804475 => data <= (x"1e226c0facec0a58", x"b98cdd9d791dde9e", x"29e35da21015da9a", x"aa4fe1bf0050c10a", x"fd63019eaed129f6", x"1522e4a890eaa7d7", x"84ef2e79bfe2d578", x"683f254d0cc072d0");
            when 7601224 => data <= (x"db5b9d5118e6d6ad", x"bb63431f9f3f7304", x"4dda4defba4dccc6", x"308cb5a231f85823", x"16ae7af748e4af02", x"fa0b840f4d8194db", x"bd9d5014db9e7e70", x"3f35878d534eb774");
            when 4376951 => data <= (x"58db59db0cf8d967", x"4d220869da5a83ea", x"977937376fd45d68", x"7abe625dea78d323", x"c536f15ea0a99943", x"56ac03ee66f05ae4", x"e21170daa95c13d9", x"d9112f943ee3e0a2");
            when 3765242 => data <= (x"9ba9b125135f4146", x"949b9b5d93f0933d", x"15bf95bd69e52820", x"61923c85cc2b19a7", x"5c8549cef4faeadf", x"2b71e729021e50fc", x"f210c95a331ccdcd", x"721d07e528aa6377");
            when 7954658 => data <= (x"b2f9b1b008b22697", x"b45a6fd90c0ccd10", x"ee5c01fa2aa660da", x"9abfab3753498046", x"96ac25dd695b2412", x"7ca3f3df87967ea6", x"f236219f192d5744", x"50c7438bc113807c");
            when 11846316 => data <= (x"ca46d47b8a1dd463", x"fbf679c16f4ab9e3", x"1fe0708af4c0a790", x"f3effb751f2bdfa5", x"fb153bc57501f776", x"329fb674f3408c52", x"2e7e4e5ba66e65ba", x"42e7f6b8067af3ca");
            when 3140712 => data <= (x"8bf00209e06c4668", x"1b6a124d59734454", x"d1904e908db54a83", x"6af2d87d18f7255a", x"576b9f7efd3b87ab", x"dd2d5d13f5bcd2ae", x"8218a9bc01ce3d42", x"44a651e34cd28c73");
            when 4032580 => data <= (x"8585deb24f88a3e6", x"7e99a06ad1ecacc4", x"091c278374f3389f", x"3c0a46bda9540630", x"94d7fba0778091fc", x"b4d7a8de30ec0ed7", x"bcb23640b382030f", x"f9caf0af0868b695");
            when 31282047 => data <= (x"e6bd826e81ef14ce", x"7caf30e82455a266", x"9d9829f2efb05060", x"2f9e8529a113424d", x"bd8cf9617036eb10", x"07b4e33adc57a2d6", x"8a2ceb217c7fffac", x"f00695116ce76462");
            when 1643066 => data <= (x"07f046e2a71990b5", x"273c8044e408f9c9", x"a6e55b3c9d14998c", x"46e200e83ab1211e", x"3c3c291d0894537b", x"acf7a7389b1b3dd3", x"4fed671740478225", x"66d533295a2d69c0");
            when 24530926 => data <= (x"13313e421477ba43", x"91bf7acd7833b2d9", x"8ef7fadc04cbca37", x"54032fbf00b5900b", x"b76f0fa7cd6736a6", x"c219dff96f6b0d37", x"ea6ff31002298db9", x"4821962a4f512605");
            when 2953295 => data <= (x"003fdbdbf5bf3d94", x"dc20305aabda0d32", x"e762535cfca9ea8c", x"cda030af1e44f6c7", x"ac978c3ed1d735d5", x"e770d7f5a9cdebf1", x"977c724586e3f084", x"5a4399e158f03c6f");
            when 5579085 => data <= (x"d77b2e71f5a6d4d4", x"1d22b891f0411200", x"60e0d679133b0e78", x"c7a7cfabf5b9268c", x"f8f645d76695175e", x"cdf89cbbf022a967", x"29b7988c5c55cfd2", x"3d61ddf38b813cd4");
            when 3702382 => data <= (x"126d8bf87637048f", x"27c672e64c5430c8", x"5655f5e944f639bc", x"a1dca82b0b5e5b14", x"9c21577ae140cc5d", x"d5702ee83fba73e9", x"8a9b68dccf752fad", x"dc23af0bbeb55b44");
            when 17310610 => data <= (x"0ede84c7386c59e2", x"3b5521fd49fad3f4", x"341181549f565feb", x"fdd77d37d16f67c4", x"549378cd856e1d77", x"2c27bf5b5ac8f0a9", x"0b55eef6642bc5d8", x"cd6963e0eb8252e4");
            when 28261543 => data <= (x"d2ef5ebd298492af", x"1fda512b146c6722", x"5bf58a5104837139", x"c48ef51122e2d209", x"ae0e2508146b3b0e", x"3372c93b9629c81d", x"bb87a2308a679a43", x"7996e62c672f1a82");
            when 1512957 => data <= (x"99f76c637c8bdbf2", x"7439498e48ecba3d", x"bb5cb9e098600612", x"12db254efee0cc26", x"69d263b4b74c8e01", x"b2464687fa56765f", x"e51015ff047e6686", x"12cc2ca67c28430e");
            when 25446194 => data <= (x"61eab5a53472654c", x"f0858639e313dafc", x"344e7402346b53dd", x"4bad55794719dd9b", x"4da81b2f69bf84dc", x"cbe81914ea1073ab", x"fd9c242c63658c80", x"7a8625ad091d886e");
            when 33649677 => data <= (x"0f6dc4737b1ddc47", x"c8520b61f7c9f462", x"8f212103ef094424", x"58b1303a9d383c10", x"c84d5d03461cb592", x"2170f91f7b89ccd7", x"4f7b074367e22d19", x"3aeba93211d1aedf");
            when 23213008 => data <= (x"e336e272a6ff00bf", x"6a1d473e4c9dba88", x"30eae5c4f4b5b74f", x"aebaef3ac34ca6e5", x"0e845255b6a9a4c9", x"fc9f653db970aa0d", x"6ab16cdc32b06d21", x"2f224a5f3a326e71");
            when 10481356 => data <= (x"47d2520829bb1db1", x"934db24e6f34f8e4", x"1c2cdf15bd92eee2", x"e95de55fdaa882cc", x"28494278da3f1af9", x"69621e8ddf1356a1", x"5bad3643375f1562", x"5ea31e084cceecb4");
            when 7303955 => data <= (x"88150251a1f60933", x"df4b289b9d688949", x"40382e52e2aad820", x"d1c4b0d7ea4a630b", x"94fc8e30dd55ff0b", x"56ca52d0cdf2d6b3", x"2467a0eb5f7003f7", x"06d63b1d7aec3a84");
            when 9622761 => data <= (x"b83cab17ef2ce78a", x"3b4d341bcf825cef", x"e2cd9774070090ea", x"4333b1ac9f70a25a", x"bf19c50999c0c2e1", x"3d04f32c54e7e421", x"5c01b6fc615749a4", x"a369eee148ac940e");
            when 32354329 => data <= (x"a0099ed3e2e41eb6", x"db3875fe8b57b78c", x"e19023c779f88a74", x"2779dac2fc44aac0", x"d66eaa47f5272008", x"48b2b8324acf3aff", x"432a5338e1f0e199", x"f688a56e5ccae8a1");
            when 4513461 => data <= (x"5d84e8d0cd2fd57b", x"d7964635904414c2", x"7945f12eb0c4593b", x"6c4b8c09078e491b", x"175cdc5df20cb6a7", x"3eb547516b67e24d", x"32d29882fb071d7e", x"fe3d5ec9a7a21f6a");
            when 10935870 => data <= (x"517f5d0ba3c620ad", x"6402688203c7d7d2", x"8d3dd742ca931b06", x"91ef23fc2e568f70", x"89affc9fb15f87d8", x"2f8a63565374620b", x"da325c14773f9947", x"6f883fe023f9b8f3");
            when 23603351 => data <= (x"b0e6a7f908b30f9e", x"0f8e21ff53380668", x"4e5e96f1730dcb05", x"e31408172a264a5d", x"043565292c4a286e", x"06dd5edb51b45c49", x"e15268c09b24a5b0", x"89e1028c04e80137");
            when 25021831 => data <= (x"06a52ed5f7c34de2", x"dedcc29cf0a6a6a8", x"a81e6d4e310e04b9", x"f8aba56102017f96", x"2a5dc03c55bac3c7", x"bf4ba4a2d9f264ab", x"6985365b221daa37", x"d561e65f3bb51706");
            when 24592896 => data <= (x"f82e59205f70bcfb", x"bb29740ec7d737fd", x"6906713fa54d0784", x"e664e130c75ecda3", x"009f3437c8125ea0", x"ece432441560f988", x"54f574cd95b8901c", x"4c502ef74611a595");
            when 16561347 => data <= (x"b558d49af365ee46", x"a4104f1fb314fe8b", x"905fd9a022df64d6", x"9354683d2d68307f", x"470a9c2470f7d3d2", x"9708aa48be3ef0f3", x"2b339789486d4ece", x"5b82175f17bd067b");
            when 32736166 => data <= (x"9c1a73f5e2435b2a", x"70ef0c693bd030b9", x"ab6e2755cc94fde2", x"2f2246657f832094", x"6c26f608c8d197d0", x"976fd947f8d4a724", x"415062f324b44513", x"c2e3a0b530688a29");
            when 14167506 => data <= (x"997c41b0713cfbdb", x"e20231f30eb08aeb", x"9b08ba50a26489f4", x"336f840c16d1b7c7", x"37344a3b2bf9959f", x"e5d17882df72e38f", x"8f22eb10cd5d7281", x"121c4620a0644dcf");
            when 6538319 => data <= (x"27e2a82c9b039697", x"a2d8498c3616473d", x"58125de635b02dfa", x"8b876d491e5959ca", x"66681813fbf7a053", x"62f373ff23a83f47", x"7137ace765ccc433", x"b9fd58c579b053c0");
            when 11769785 => data <= (x"e48d03f8218bf95b", x"31cfd76c8afd3b09", x"457e3c1cf37b00e0", x"25426304ffc89fcd", x"6ce93a79e431c0e9", x"3e168eff731f5ad8", x"e9f94a30a1537268", x"3663feb6942ff730");
            when 31501655 => data <= (x"f06e0389dce9d799", x"d78e579d27499f23", x"843bf8798d8a691b", x"1c5ed9c2af7ada0d", x"ad39f68fb4a52537", x"88eec1168f80dd75", x"31b0e83aa4d089a1", x"80e587c28c34fcc0");
            when 32209325 => data <= (x"5463526c78743453", x"f1c95947e61e59b7", x"fc7c09b9846121cb", x"4cddca0d0eff202b", x"2f42f2351270edc3", x"bf1877c70a426850", x"f665453999b758ad", x"eb039190a58b0acb");
            when 20009968 => data <= (x"25253ff3f345207f", x"acfd00384f73db57", x"00a9ff464deb97a3", x"855f66be85b0423a", x"7e4f3edc85b5319f", x"ce2ca882c62cbe6c", x"d5b16db00185ebee", x"46b7aef41ac58923");
            when 27357062 => data <= (x"664a33d0fc5a6e18", x"017f47397a317341", x"7a5438ed653a2d51", x"967325a0f3b4ba74", x"a8d67952bd919476", x"5858b36b442b8673", x"87b01335b270eb6e", x"41c74fe88b900c34");
            when 2210474 => data <= (x"5914df9422e1da30", x"31d024a238d94185", x"ed726f40934be7b3", x"930a326479339eec", x"d894c13457392269", x"c92698714257f101", x"9cc024f00a5d799d", x"a01e607c32745b74");
            when 19997754 => data <= (x"accd2c6457b2ca1f", x"10195cd182c5062c", x"44072547d49576d8", x"36f5e84d081d8d1c", x"59523bf6e58ef649", x"dc91deb11843b171", x"06139dcaf13a02b4", x"8333415947ce2f88");
            when 17015868 => data <= (x"ee2a036daf012c08", x"32cebd5599991444", x"9a7de3e65ed53a4a", x"6db8da1337221cad", x"284ecaff91b4df1f", x"939ca9334ac4377f", x"510dbf0011952958", x"e574c78a0ea424ff");
            when 17101485 => data <= (x"e393905c18a56c10", x"acabc87a58679644", x"faf49210f9d2a7c9", x"422a4580cc91b9f3", x"0d11ecf8f5a94522", x"cd88f8a6179fa3d5", x"5c96494e83a81611", x"1d450c177182e863");
            when 31379959 => data <= (x"13bd233b24e40504", x"40a4fb08cab555af", x"e2ccbe74b89bdd11", x"a03ba4a6ed915add", x"7e1311ba613624d9", x"85750d14b23d960b", x"4616e0c7a39ef6d1", x"03237e175aa81143");
            when 21063180 => data <= (x"ff8ec4c117f88362", x"d4c88791a5571326", x"6d9747e4eff2482b", x"a6d0a2442efab7d2", x"04210276b3526b1f", x"a9a06341819d3ee8", x"d7db25106f042138", x"65b9521804eb0fb4");
            when 12861979 => data <= (x"3db8d409417e6ede", x"bdab64c1a3708dd5", x"2a6d68d5a49558ca", x"15eb62a701db87d0", x"ed6e1e9bfa4453fb", x"e0cbb44a004f381f", x"609e1df3f2bbe2ef", x"184220147d0d81ac");
            when 27040885 => data <= (x"7f09c6e2f9106ace", x"5e55f37a8da9246f", x"44500dac43325feb", x"7e30bbb0f06936bd", x"adf8cc50317eb7b9", x"d16cc4e60184e215", x"a760926848d8880d", x"6ae1c063a3d2fc9e");
            when 7042128 => data <= (x"3323965803e86c26", x"c7bd102f0bd05e5a", x"bddb5dd5f8fb091f", x"3b06c450f597d093", x"a9d61b53155c8c83", x"0e9c56ffcc521edc", x"16770fba1c12e566", x"9b26fde2e6a2c290");
            when 31486179 => data <= (x"aa402f5be5951cd8", x"92d24c53d9be36c8", x"39483aa1df786590", x"4b90e3172e5dff6d", x"b79c0b39ea6deb9e", x"796cb88ef7224c8c", x"eb95a580c654500e", x"1ac82ad25881a99a");
            when 6201981 => data <= (x"14274674692488be", x"b26f6308ecc23047", x"f9cef080dfee3476", x"de94ac8be0360ef6", x"771982c2c54cbb6c", x"bdf106f78227aabe", x"974b31e023e57cd7", x"35d4c9b84fc10c72");
            when 30195259 => data <= (x"49fa0858570580de", x"a0d7eb8398958d7f", x"407b72b7b3927066", x"9d3dd991be9c0279", x"d26bd367ecfa1cc0", x"74bf815bfa91edf5", x"f899eb087ef4d9f6", x"f5682b51f4908e8e");
            when 31457951 => data <= (x"ad0b9edd8730eb89", x"28b1c259f2f98818", x"bfd4ec232de25f49", x"c4365d237572939b", x"ca911f0050b5bb04", x"3beaa9cfbd8ec33c", x"aae1658a0325186d", x"38e3e8ec3e5c187a");
            when 5516334 => data <= (x"29727acde7dca43b", x"ddd3e30611ce07ef", x"a3c20b0ba1d9fe7c", x"5f31a119e66d8015", x"1234db1d117557d5", x"e60a4f5e28e99015", x"df1f167c56e43cb6", x"8b90ef7a166dd1b4");
            when 33008996 => data <= (x"5b3d22167b0d8997", x"1dd9d12d23d9a273", x"af0c587085d4d115", x"a72957b0720f27ae", x"f76783220293328c", x"1485def1fb51f8bf", x"628d7fceacd0cf20", x"9df9a35695f15ddd");
            when 2135282 => data <= (x"49e1c20a1b1c4b92", x"6e1cf57039d5bb62", x"b82ec0066a4b4d01", x"75d55441e8cce1a6", x"8332312471ffce93", x"2195d1b1895c7eeb", x"4dd43c965de8d36e", x"f4db18c90d96c461");
            when 11436767 => data <= (x"d1262e2c72c9109a", x"b03af69832aa1850", x"625d77d5062a618c", x"15450e8d624e3728", x"2bb85d3f7a7e7ef3", x"e7e289ee4d5c4f2b", x"e0d2d3f6f669e4ef", x"182f7b7534777cfd");
            when 548760 => data <= (x"a6d272f60b28ff6a", x"d231ce5bba0977e6", x"26862beaed7a27b8", x"f4be4e9e47fce57a", x"9b465a2d297ea0ea", x"6f15ff239ac2de36", x"c023fd5be424fafd", x"dd3e37c83e144c3b");
            when 16619641 => data <= (x"d4b348d0ea8ce41a", x"5b721e970d1a8ae2", x"e1c6c33cc13f8a23", x"1a86aab1f2a043c7", x"881aa50873468b92", x"4a7508ee43f13796", x"30d42df1f9ef8abc", x"0511c85e79f63766");
            when 10219024 => data <= (x"6ab6f53f396a7013", x"e3654b438f04f1bd", x"8436e5ac104dce43", x"e4bc7819f9da4968", x"f641485a6211b8cb", x"5f31b87275c4659e", x"a4e5cdb217663109", x"d34a7294e0e34192");
            when 6008935 => data <= (x"e66ed60fa3928c60", x"d71c3270fa67fb5c", x"540808161c992b11", x"7376127fb683ea63", x"44cd9404025fd5a4", x"ad141389de9c7f5a", x"a6d37eb89f8e8add", x"6f8642050d399648");
            when 3403255 => data <= (x"0147a0bc2c9e77e6", x"9d66ae02dfc09746", x"2255105415244eae", x"313bc1c38799691a", x"f66843609fb84bbc", x"e641fe36eb5f4404", x"19982a69676594d7", x"0dbbd3687e26a230");
            when 16820731 => data <= (x"d81b89c04ecceca4", x"37fcc066fe9aff97", x"686f1dc203fd1d3f", x"885a4b011211e0d8", x"c4c35ff5f6800b58", x"3026c7749b749e45", x"aa4fcc64c5cb0ad7", x"de50666acb11fbbd");
            when 21739880 => data <= (x"aa0f8fabc8e40b55", x"fdb3827c081df772", x"0bfa0c466e24f42a", x"a219d80611894226", x"f29b0a75c44dddf2", x"ec098dc3ed9721a0", x"ec56ba306cabdd26", x"f37633be62e9cfed");
            when 30401496 => data <= (x"f8ba76a85270891f", x"a65fe6357486b047", x"5c9ce647011b765c", x"d673600b04ad45c7", x"0ed32c0ac48bdfe6", x"7304208e06ab75a1", x"389417501ea75164", x"565febea1b26c94b");
            when 32744008 => data <= (x"cc90ff93640bed8e", x"2f25f0199a50d7f9", x"5fa70f276a65ae7c", x"23b4c1feb6a8469f", x"40389a7088091836", x"34f7fa1645a5bfc9", x"49d3b4d646f9cc11", x"6ff9015438f36fad");
            when 2709019 => data <= (x"2129d6a7f1729333", x"b4c798a94023b2a4", x"68f0240ab043c1e2", x"70ca935c8f85a808", x"8ffb71fd803cec18", x"266701c89cfb3607", x"2f855ae87753c7d3", x"5ed059b48c8c1f27");
            when 15306186 => data <= (x"9df168a28aa06da2", x"1715b46b15ae8fa5", x"294ecb43f9fbd6ac", x"ecac1d971d6eedae", x"ab929c73b648a4a7", x"1d63dbf1579f73d5", x"770e12056e23a166", x"1b1fa797c6a3a3cc");
            when 10237987 => data <= (x"2286dbcb032c7f3f", x"9d71cd7aed905be3", x"7a6a9bc6465f81ef", x"00f7b8883ea877d5", x"5c508beb7310ac05", x"287c37cc65e8f390", x"3a591ff94fcafe69", x"01d26ddc0b3dd2d8");
            when 20720632 => data <= (x"fe355d2e09d5be9b", x"e1eb7aa719f38c07", x"5004b260fe31aff9", x"081656454c500e31", x"dc89726e923b4e1d", x"7bb9a3da06c65fc7", x"a57313a03da1c563", x"dd9fadeefbb5c415");
            when 6277139 => data <= (x"7f1bf693f91deae0", x"c042979d1996cb4c", x"0afacbe482346dde", x"3243acae3b192d92", x"37b398aa19255cd5", x"17e9c6cbae54605f", x"fffdbfaf5f3972c2", x"fba7e86f79dfd16e");
            when 2465677 => data <= (x"7725cd5b7688a739", x"8528f72d9cb6d474", x"46ef370c6d757a0d", x"baa20d8d43aca07a", x"7fe6281d79c97149", x"a5fbaeb3619b4d2a", x"bc94a931c6e46d9f", x"f55f38b97a764e6b");
            when 12856420 => data <= (x"fd4d3d9e27c3496f", x"d32ac5d1369b4753", x"ae8a5f96a8f3c9c2", x"208659e6193706ab", x"71814116696acbbc", x"63460df67015b075", x"5fe68c8d8437d7f4", x"42f17c7edf233dc9");
            when 20329518 => data <= (x"f3e39281eef8f00d", x"b48d5416b481d1af", x"743f4f5840f8f11a", x"ad8b96aa9c382fba", x"980267a1929c2551", x"99971e7e90644d1e", x"f9651d724d9d7227", x"610f2f1f8ecf6082");
            when 21936241 => data <= (x"58ca45ea60fd1925", x"e59ba9478370bf29", x"9521521cdd704fcd", x"d52c5e5b31915f9b", x"d0150965bc487fd1", x"1ea581c55663ce84", x"c838a4bfdb265e7d", x"e1e280fdbd357396");
            when 9568667 => data <= (x"63dc1cc314c4197d", x"e8040e4cf33b6242", x"7dab3f82402a387a", x"b2e08efd0e817cc7", x"b247757abef28c11", x"f9e5bc093866af4a", x"03f2184f9cb863d3", x"0cebdb7c1dc5ad4d");
            when 29817726 => data <= (x"87fbafe56d3a528f", x"b777583f34e35e70", x"88f32894e66782d4", x"ed76f1839c92baf8", x"a0f0814b22f9db81", x"03e32559d5f7446c", x"f05ba65690996879", x"72d406b3016e0e6c");
            when 11447314 => data <= (x"330136352767669a", x"c79891a5a6c240f9", x"c35004e782e0ceff", x"ac2bf92f8a97044e", x"60cc0b582b1cffd7", x"70a1c994d03faa9a", x"33dd89b2cfeb05d5", x"e58514f3c098b2f4");
            when 2050374 => data <= (x"0b41bd6a94820288", x"52519b1468b0a46d", x"28fad1f8a5e5ea63", x"8af9a20e60b13a45", x"23396121647c887b", x"b55db24f59576211", x"33ea6e2077dcd28c", x"faa596b991b1d222");
            when 14637940 => data <= (x"6eba48ea65d7dc61", x"bbd9daf331cd01b7", x"ef1f84edfd17f813", x"3d8f17398c5ad633", x"592b4251369a5d8b", x"8fc06f6d7bec05ce", x"2860a4565e211203", x"d3723c1c01b7ea9b");
            when 1128366 => data <= (x"fbebd1e7220d795e", x"d24617b88079b48d", x"e2ff360a3d7a71b8", x"866b75dbcbf18769", x"2a2d17eec30e8fe9", x"a23f8044c9f46ffd", x"316dab17ea02ae66", x"d59b6303bb9adc26");
            when 28881679 => data <= (x"8259f2a71f7ccd17", x"e679c6a9bdfc3a3e", x"8e1d4e22f87f5415", x"e7264a16f0c5403e", x"e6e78c9a2b6af2da", x"e2d7d64466c07b27", x"5bc2dc28cea9dcd9", x"734740139987231a");
            when 29462186 => data <= (x"8d16696cc097e88e", x"4025b211f39ce2ee", x"99c80a37ea03529a", x"ae9cfdd5b6de7298", x"d57ec5588738594d", x"2607e860e49f5cf7", x"d9321c1d63346423", x"0fae7d0054499b72");
            when 15309196 => data <= (x"fe24709f5b4debd8", x"e2b6d014c25dabb4", x"56b3ecf036c060a9", x"d32cb363b2d52d30", x"e3fa8d178d0b8106", x"923ebfe2e30c8def", x"e31244543ac2c389", x"1c18820b54066051");
            when 7091682 => data <= (x"344392cc2e3ba1c6", x"90d0e332bee1d66b", x"7113560476ed4ef0", x"7c43c43a920aa602", x"5bbe23fdf9e63573", x"9028566b15b939fd", x"c5572842509fd0df", x"9e4d5c3f88cebecd");
            when 14460312 => data <= (x"ebc6cefaf674da31", x"d7f48b4b6a063c1b", x"f6c2ffcf4a11818a", x"3ba123e0bc548dff", x"67b5fc2bfc7bb592", x"8fa903a4cc5c7600", x"2c3b7967a51a3e27", x"a74137bbd920b1ae");
            when 23034032 => data <= (x"1e416bcb069b31b8", x"24811976df4b2ee5", x"7e634fb6e38d1f01", x"2c989f85df27f3a5", x"d831fc6028b91281", x"d18ccdfe238491f6", x"46042d7de767a821", x"18d197b899ca1491");
            when 14452439 => data <= (x"51fd4cace93c22da", x"494714cc66ef798b", x"15c5e25ce054fa5a", x"046076444191167b", x"3f9433b01205a753", x"056183d4b6c18683", x"1e8f887c1050cafd", x"34f1406762593a40");
            when 4120288 => data <= (x"a3f13d5520d1cb39", x"522d9daf639f35a1", x"8dbf0d05b86b477b", x"b409d6a543b26820", x"144fc4e886ce4a4b", x"ba58a7f620d7a6f9", x"5544f655795e2848", x"a4759917b62ea32c");
            when 14758456 => data <= (x"3d749013d2285db0", x"d990c5a34bc4ec1a", x"09f9b2bb26511e49", x"037196cf2979547d", x"0dfd1009b1a2df76", x"1d3ea45d708c7557", x"7b835ff560a76d13", x"09a3910554235866");
            when 14044379 => data <= (x"cd3ec8d8dd93faf0", x"81c5c1247d99ecc9", x"3ad273172e966ef2", x"457949e9cb70c215", x"db0def1f8ed21c26", x"c8e665914df2eba1", x"5e725f1737a07e7e", x"f7a4dffd564e03a4");
            when 32509555 => data <= (x"93b54476dfce4766", x"f4d1056ea77cf6f7", x"1020cf4a43822f89", x"110559c4b670432c", x"6a40cf68d89733b3", x"d031a4d759cf010c", x"9b3dac7cde9d402c", x"165f8aefd3b63ad6");
            when 29562823 => data <= (x"2a1393061a949483", x"1d337b112c16e200", x"9850146049179806", x"74c589b2c489d67e", x"24110c5d9d963e8a", x"7893f69c44803f44", x"1b3913700abba43f", x"dbf5ec922d6a2dc5");
            when 27564607 => data <= (x"b6790aeabf4c5a2f", x"3980881e02abbd05", x"7e1bad5451697741", x"a902c820ce2816df", x"b7924c63a0e33459", x"b29c32e1be495fa8", x"5f14c9c6db17e4de", x"fcc75edea03c6e99");
            when 13105527 => data <= (x"8024136968f1b91d", x"d704febbb747961b", x"24728bfd2e053825", x"6c256b081050c0ba", x"140d6fce62158c81", x"963086bcb7e061b5", x"2da5d1ccaa7f594f", x"2383d3e93b136447");
            when 9586558 => data <= (x"8f8bb296784bd708", x"c814d37abad591fd", x"0b8fa5c33019e4b2", x"eefd46268e4e9c22", x"5dd2035907e293fb", x"da5e5acd5a15f816", x"bba6a6c2ad605e82", x"80a5a0002aec2ee5");
            when 17213306 => data <= (x"08fdc458fbdeefc7", x"bb6b7deea1dcee1c", x"6a7538ec3950b5a9", x"d9ed7a312f4cd31c", x"cab29c520f8fea42", x"471b70c5e1954c33", x"573f8ec77dd56599", x"4ca6552c3743d47b");
            when 12032836 => data <= (x"35e5e996141dbaf0", x"177c0d26fabf42bc", x"cba8f4bdbb873ef1", x"17b48a820e0c6633", x"6a7b68edb33e3025", x"f2b871cebf3d4f62", x"3c3783bb7b2fe855", x"193e3ef3524d3cc3");
            when 26155399 => data <= (x"590dcc04294d797b", x"4714e233936b4fd1", x"aea672cec5ce28df", x"edb84d0c96b62e43", x"d13bf91e31d10779", x"844ec37c2f644174", x"ff27bda6d27d4ebc", x"9bb4e9e8add64aed");
            when 24888439 => data <= (x"60dec3a10a3468bc", x"b50003e1fbdba4ff", x"0a6149bfc3f6597b", x"f24b504a9260ee94", x"31724cdac39013b0", x"fe80f3c2753d1396", x"18ef1ffce42c0bed", x"f6e872e5eb524b20");
            when 12432472 => data <= (x"2e152bcf121c517d", x"c28b78d5a40f7a5f", x"39156573fbbcb7a3", x"ff8c3dc00058a8da", x"86f74b0a7e81adbf", x"125fd6b9241801cf", x"0061f37bf7fac19d", x"07c069009c0415f0");
            when 788694 => data <= (x"ba1b16c9ced6f7b9", x"b1ef2908d5dec4a5", x"fcebfd4b2a140073", x"cf6e247182ca49aa", x"efef5c689e6eb0c6", x"81e2b550709580e7", x"99cda2a28cb18f2f", x"d6bb2fd1f8561a87");
            when 20525441 => data <= (x"952a96cad894bafd", x"f9b7853a506c0897", x"36f0d4f9c4350e68", x"577589ed2cce3a9b", x"45d795a37775529c", x"192aa5e8a3278859", x"da879c3a4cf3161f", x"211efb3ac0eee4dd");
            when 4269200 => data <= (x"7fdf4653651177da", x"df2a3a6bf44046b3", x"7a9381637fcbb723", x"debf911929e7cb69", x"c4014b5736c7fcdf", x"20e416245e3ff0b7", x"87105ec21d25452d", x"ec501b077b324fce");
            when 24593673 => data <= (x"94d8c4fd8a927cc4", x"d061147016dbfee1", x"5ff5ee15ef3ffe91", x"4006ba5f12a32170", x"437c3b41f50158b1", x"54ae38136cb8e300", x"9dee978d463f4658", x"c047980be7ebdff0");
            when 29654390 => data <= (x"7af9f7886b672d7c", x"59654dd079a50e66", x"b293ed80b9ab1fff", x"83721eb43b3c96b8", x"235c16b01eeb226d", x"3cae2bb0f2bcdc69", x"4505b814585b5190", x"ce5392c5d41171e6");
            when 30568809 => data <= (x"96bc0d0321704d4c", x"efd75f1f50a2d7d9", x"0bad6d02a94307e3", x"0abe00301c87edbd", x"3b7edf10ef6ad92c", x"dcd21412d0d888d0", x"45c9f4454f5bb74e", x"ea5ac74167f289c2");
            when 4390467 => data <= (x"c800628a499130a9", x"8c532f16c96bef41", x"f3ef2930bea96c35", x"7931cca21bbe5daa", x"bc04305738ab1b36", x"e50ead41bebfe098", x"8d1539c6bb199a74", x"4e2c527df7c6f0c4");
            when 4361461 => data <= (x"c0c49e9b99ddf813", x"78dc777e767a4007", x"2d6cafc5273754fe", x"95d4f4327ea9231d", x"83086d7e1c69c4e7", x"3cdd90b687c607ba", x"3aa50a707a6f4d8d", x"3a41068ef1a60e6b");
            when 20656736 => data <= (x"6937c9824b26fb06", x"4c1291160ece4961", x"3c971f04b3b3b827", x"63721a0aec074d61", x"11ae2a55c77e922d", x"4e2fc3dcb42b48ab", x"2e36edc502fe3d89", x"150241064bf5fb84");
            when 7823603 => data <= (x"d55ae8e148b1b7a2", x"9ddd048b956488ce", x"f9bd8d5913ad716b", x"829771fda9c31a9c", x"3a43e5e866711edb", x"9983dfdca3c83bba", x"4919015c4c73c2be", x"e9a850a5c64e64f1");
            when 23367906 => data <= (x"c9c21fa3c0eaec46", x"7c65c0ebd2e37272", x"b29a326fd9243aaf", x"8454dfc4b33e94bc", x"f549322a7095ce6e", x"acc95559374f9661", x"e8e4e358c13168c8", x"85fb69fe62ef94b3");
            when 12002173 => data <= (x"44835ee40e642f9b", x"98f2bc1a235749c7", x"fd3e9f5ccac7294f", x"2121c7350e878067", x"39f626b0af1d7573", x"8b17eb8e0a90d2fd", x"527f5e7e040fe6e6", x"6a44556899a76cc3");
            when 4716794 => data <= (x"5a8f6533d9a1aad9", x"de64c98ad1e33adf", x"89e3e092c67def44", x"7809caee7404c739", x"0e2139be12614a9d", x"9ff41c8323d35133", x"d89e5bc671afd7e5", x"0951391144003e46");
            when 29439137 => data <= (x"eea1f1a1bbf21d5c", x"b9c9e45346d8634d", x"e36ba9a9c01898c3", x"f2e880170502b454", x"e5d835059564af6b", x"f73665f29726ecfb", x"c116a834d5bcbfbc", x"459c9c2dad27392e");
            when 9289752 => data <= (x"4e596dc262a42b00", x"b7ccac4fb9767fe4", x"0bb4a0b0153d8a2b", x"1b3118f929824317", x"5f16c1640c577868", x"ec35ae23a8fdbecb", x"2c9fe303994d7dc3", x"939d2892d45afb7c");
            when 1295634 => data <= (x"a770a4a01f931c35", x"7a1d47b5472d0180", x"fc24d822d4d9175c", x"f3f465c13ce3a772", x"d03d09961e583539", x"f6ad26611182249e", x"42f03ee20f525df9", x"37eacf7262a44371");
            when 21156543 => data <= (x"f4646947f92a48b7", x"7961117555811995", x"bbcf2ba09631dfbd", x"290125b71c5f7953", x"9f12c706f1977f3d", x"c7483615393df72e", x"cdf5fc8805800aef", x"1dd1ba5600168fb8");
            when 31452599 => data <= (x"3f1916eedf9938ec", x"7625b5f3d65f1a15", x"652459e702a30701", x"763bf80cc542755a", x"b7c1973b815dc97f", x"5dc9964585ff43d4", x"9f62c935246b0a72", x"6493e97723cc3831");
            when 21364087 => data <= (x"9bea5ac6aee47646", x"d24939cc8052792d", x"747d656e516da6c5", x"ce9009d33c8f8b90", x"5a41d05c3496dcf9", x"5817041389dc4a01", x"46e6a03e67733c82", x"d3b2eaf492ef59c3");
            when 17897798 => data <= (x"2de18b825d6d28ae", x"0aefc219dc689d18", x"aac42088d2515a73", x"b3d5c7d8da508f23", x"b9bb417d6c960414", x"f4e7cb3d46d43786", x"d13c1e4e6f643f81", x"b2a5ab54d5b33ead");
            when 2679712 => data <= (x"c39a516893c4d57f", x"f99a56b491314f26", x"482ea1e50d354866", x"750842b3b8744b33", x"b618b3213df84c16", x"cbab34e8deec46d2", x"bbc28faf72119560", x"81a9d63c6517c68a");
            when 551156 => data <= (x"961f2ab664fb8418", x"1493d1c849bdce25", x"56f457d825f9c781", x"c9e4e60b075c6f59", x"9e4af128365d2e34", x"c70cf0984caf6804", x"81b6e5a942c38e77", x"b1d1a8bae617c316");
            when 6870409 => data <= (x"f83db4060a3c1419", x"3e25e788f0acc35e", x"95ac43ccd6faddc4", x"7d58055bc772101b", x"0592d422114dfff7", x"ac85d12c34ac61be", x"b8fbf9464bf8ab1f", x"321c73d00a02b12f");
            when 22829441 => data <= (x"becdb3977300c50f", x"25c83b42a6fe8d51", x"9d2716732d51e7d4", x"1e4a8ee7f54fd062", x"fb56fdc47d6476ff", x"b6857f100c8de059", x"dcc4d93cc17db55e", x"398dfa00d0784d28");
            when 13513402 => data <= (x"63f1bed2ac8d9a25", x"405fd97e1fc41998", x"d340e679eedc3979", x"f9fea25c1bcb7be0", x"555aef4346996b9c", x"2f88e8687a90d2dc", x"9ea88d8d8a18e492", x"db15b14117fbf33f");
            when 15833945 => data <= (x"02e1ba696830fddc", x"29c443a57414e820", x"87efa7a8bc29af84", x"f693bed47b23e8b9", x"af75c6cb0032c79f", x"f5259b16a141cbd9", x"d6b2f5fb48cc7a79", x"641738bb9cfe35ec");
            when 31076612 => data <= (x"7e8a1c73b87899dd", x"8a65c2b75fee2e99", x"6e97400f17abdd71", x"a04fde1da9f3a020", x"e045d0ada3827cd7", x"17c70d496cb36fab", x"06457b1a67704ed7", x"c27e317da935b908");
            when 15165795 => data <= (x"4ef7469d9d997170", x"7e7abc482429f7c5", x"33e4b02ebb07bb25", x"219db4a518677664", x"2833f4a4dbd7ac04", x"a52e97635e211f72", x"57de8696b83c21a2", x"4daa09445fe8cb60");
            when 29308165 => data <= (x"d30d7aa3bb2923cf", x"e58c1fe7691441f0", x"4889443fecd99d8a", x"f59f5c6cc86574ef", x"b68f4895a252fad0", x"f33819a63f1d8ef2", x"f4e77ffb6a6d68c3", x"c27d6e9bd048786f");
            when 9157404 => data <= (x"54f7c335ea0f2f8e", x"4d2af4c4a293de65", x"7cbe03e585c46ef6", x"64f5c52325d1f03c", x"c21460c825a109d4", x"5d9f4e171b8fa9a5", x"82c73ff4ef85cb19", x"6dc19fc1b7fba609");
            when 18531904 => data <= (x"0faf13deb52c52ca", x"94c4a66d3c9000c0", x"530f97dfecb1f891", x"19b001020744e683", x"a92a60222ad09367", x"fc1d045e6969a1da", x"7376da9fc84702c0", x"26970b05d2b0e173");
            when 6977401 => data <= (x"dc9f4c1d320d057c", x"f47b826432381bf9", x"827782a76d853887", x"76e858f942889d66", x"a0eb1aff6ed9f359", x"04a0307f8ef46b2e", x"cf9d3d5d87c06ca2", x"4c9cfb2dfe0eca12");
            when 18702967 => data <= (x"935bcb20b1f57b1d", x"15a8cbfe02bccab8", x"d4c3a73a129a212a", x"5be0f1da42a7a0ba", x"71def8217f5ef724", x"6e11efcf6d9519a8", x"89f066a54250560a", x"ca177644b895ae7b");
            when 2462266 => data <= (x"e9d90f323428263b", x"5c021106b84e12e2", x"e074339a3668c564", x"5bd1f158ca2cc41b", x"44b8af45ca5ee166", x"13c4df9f73d64292", x"d701755e5e2ac725", x"33aa2dc67287b6d5");
            when 22872586 => data <= (x"7200e0c0c79f94b3", x"c350e0e208e14228", x"af4209519048fa7c", x"bde7c4c626c91448", x"14c41ca6c1954708", x"e97860e214d23766", x"5d609d8719254c44", x"e0b8609e104d09f1");
            when 19051513 => data <= (x"f98c62aa96451dd9", x"980af2878017dd8c", x"86b629ce579aa31e", x"4598d0fcb6eed7cd", x"cea82d02465b5c4f", x"dbf0c9d921cafe38", x"bc5b1b632b8bf6e7", x"56e842bb035e9fd3");
            when 30967688 => data <= (x"08460ed921b67a74", x"4a552d3dcbeff213", x"7a69040a32cfdd02", x"456281b084afaffb", x"039b13cfaf0b6ed7", x"9fe8b033e5558476", x"8877a2d140fb6a7c", x"6201bfd52d5933b5");
            when 26325024 => data <= (x"801aa3fed512c830", x"3a208603d8e91a55", x"d56131ef6e5ff2d6", x"02b22294b8020520", x"0dbc611d25372467", x"2ac6a90993c0c8e1", x"f96d93c201c0b012", x"22209363dc661293");
            when 14190558 => data <= (x"cf15c5241725533f", x"76e1472cfb1e0e72", x"b08b0bdac4adbc59", x"4066b634fb24cbb4", x"ba3d8cf36b0b0c6d", x"b8b01de6b62567b8", x"2722c5689d467330", x"32e68f8c4f6754a6");
            when 11424503 => data <= (x"758b1dde1de87e90", x"3c71612fa749cc85", x"c6cfb85c27bccadd", x"39ca8bf46eadc2e1", x"7eecd7780afbe9db", x"c204628dc3de71e9", x"05d6434353a39e72", x"931a841d9336af25");
            when 10271511 => data <= (x"2201383e2d4a666d", x"ce0e34ea46ababa4", x"7c737494d180f201", x"20578cd0e79fce6d", x"6ad3051add4a9454", x"646c9a626db5af46", x"1d031574b58cd2c5", x"0989fb309a8b174c");
            when 33729365 => data <= (x"b9f843a3ae79ecec", x"6e24bdb227888965", x"33e286b84d141e8d", x"1e1661a2a40cfb78", x"d1049dc8422c431c", x"43a6ae18dc3b0c7c", x"7e2b488bff1d092e", x"970ae9b0dd4460c0");
            when 32551562 => data <= (x"1c26690956ebc2a7", x"67f2684684a3da5d", x"4d3263480ac13cf3", x"5bfbc652ed93e3a7", x"78909c2c7a352e97", x"5cecbd96cb8bc0f2", x"e975233348c15df1", x"3010f5f902cfffdf");
            when 9634975 => data <= (x"e31cab5ee8e8cb1b", x"8ca415dc8fffd4d8", x"f74a29b6a72593bf", x"858f30f7189f6555", x"503d58a3c3fe207f", x"037921b5099b03d1", x"62bfdf6575cca659", x"93be881efaf6672c");
            when 33738084 => data <= (x"d6128bf75a530760", x"625a7d6eac82f419", x"72ad6a88ff5d5079", x"3e2d0f049eb14bb6", x"8af1b0029a2f0558", x"01bb7b34084a4c8d", x"5827725ce9a32af9", x"1b7892ea48ab7c70");
            when 33655584 => data <= (x"32c27e5f46de258a", x"821fabf94f2d641b", x"beb58793ec1737f8", x"134442af51b1ba11", x"87e0e48e8bec4b9f", x"7093cb403f8048d9", x"ddd54b50b13c9b59", x"61f43d73ead739f1");
            when 31417620 => data <= (x"3ae9606911b12266", x"553e5b9903da655c", x"d660143c51aaa177", x"e22c6fcbed58aaa5", x"00c1692de2a4eb6d", x"187441cfdcdb737e", x"cf7135f44dbd7cb0", x"aa0a42d0f20e1fd5");
            when 25637092 => data <= (x"a250e69d76bc540c", x"23ea533e0f6028c4", x"26d778fac605cf08", x"f866f88e3ba841ab", x"4b368fe888fe5d95", x"1f425ee63c768af8", x"6032824ad8571d9a", x"f19c2fb7771bd177");
            when 11401050 => data <= (x"9e0d8570b7f456c8", x"94aed909ff782840", x"9e64999e69d15743", x"3f19d0fefe79f817", x"46f0e5ab35bea834", x"8be5f267d22d2040", x"23f54c00d76e291b", x"5b95cc145e806182");
            when 9005865 => data <= (x"3fbabbad23057fb2", x"530eb92235aafff0", x"454040b4def633c5", x"fa9cd48ef6f9acb2", x"b2bd9613629faea2", x"369c82cd1449935b", x"e1081f0f5554646e", x"716c9576b980eead");
            when 2971157 => data <= (x"cd9587d09c8c92d9", x"f2be612b599e7d4d", x"0bf051feb141e4f4", x"acacfc342d049201", x"feb9ac0fc1b6ab2c", x"41448f3d856fecfe", x"1b17745ee6061624", x"d9c2ed05504ee3d6");
            when 20045847 => data <= (x"3b154471edb78d69", x"01d63f2945027cdc", x"44c14c8bdc61ff67", x"7729c368cea3bd9c", x"6b520c524e7f6ccc", x"5b645195844bd381", x"d41610f00e6dad47", x"dda5c3a46fb85934");
            when 10829350 => data <= (x"bf9e9f9a42d4371c", x"a0a221286bfbcec6", x"fdd3d488426ebef4", x"6b308589618852b2", x"0b6abb4952d185cb", x"cafb4c3f6fec6554", x"13c41f4bbd74ba54", x"35c4d61242597efc");
            when 18480470 => data <= (x"8d929e58b451dddd", x"b9fe787db40155b5", x"712dd353c6f5b843", x"e1f19e8203c86d12", x"0e52fa62d34a534f", x"7ba97d67d4ba76a4", x"8d5c93784d3f97d9", x"90a841eab448b41a");
            when 16490076 => data <= (x"70fdf92bfc2420ef", x"36b5e2c37656634f", x"ab54ba49a491b527", x"891983840cb8b399", x"73c407effdd9ee55", x"c527f1ca4db9dabe", x"a1a0ef1043d281dc", x"0fdb0c4a293c9744");
            when 1543438 => data <= (x"641556058695cbb6", x"4f1e12a386351cd2", x"99390223bb4be0d1", x"81835ea5048af55c", x"d09cccb9a0a9f7ae", x"613ce003fff8aa9f", x"89db30d636b74cc9", x"b61559adb34bda6f");
            when 34022627 => data <= (x"f9ed1e28a5e3394f", x"539590bf7a48f280", x"6c929803b03e8e9c", x"1efd6c2e9e1683fb", x"c5be8eb0e03165bd", x"a26e6ad5338e07fe", x"5c60abfaa73aecbc", x"bf720363ccfae516");
            when 18024036 => data <= (x"ba79696f69e7a093", x"4cf1fec8fe513658", x"6d150fe0557595c1", x"7a8cac45fa7f76a6", x"cb2690b239ea2a0c", x"b1569cd88127d2ed", x"4992cc90ea8795b5", x"5559fe8cd1bdc14f");
            when 27087949 => data <= (x"b0116f3ccb4ed6ee", x"f48b44242b7c9c03", x"2b2bf29bf629c549", x"a20228d18f17f970", x"dd4690baa8f4cf64", x"cbd1118b1cedde50", x"ade1764b2453338b", x"b4f21e0f416f4213");
            when 27650243 => data <= (x"964d3c38b77d9093", x"22db474a4825951f", x"864f9eb11fb0ee1d", x"4f8fca35b116abe9", x"8d10210a6dc5cbe3", x"b1366069442dc41f", x"2499ff9dd70ec6fa", x"1dd1ccdc42f02887");
            when 22380923 => data <= (x"5ccc935edc234864", x"4e29cfa525c24ed7", x"06a96bd08ebd7c9c", x"d99733e6d9e85355", x"d48f5421eccbe31e", x"725d53dc4e408c63", x"c101934b8c056ffb", x"ec46f15f4d3c34db");
            when 951049 => data <= (x"3ae2e81993601e66", x"4d1ac991bbd776c4", x"11a91f27b2920079", x"c993350e170e3f87", x"25d17c532b46e44b", x"34eeb4588450d035", x"55e6edca863eac0b", x"daf887cd694640ef");
            when 5261576 => data <= (x"1145cfa50d370204", x"0cace14272f0b91b", x"a9c2a22385053102", x"0f331cb240597fcd", x"f714aa0c88a4a577", x"76455a9fc63ef98b", x"520f9ac1fa0669fd", x"390ba24d9e5dde75");
            when 27718034 => data <= (x"25a81dd18c824655", x"9f8f0f0b7bc82517", x"67f7665d66809cfa", x"b2622543f0fd407a", x"36f27be9cf2476de", x"1609bbf270e40004", x"a3d75115c6c6553c", x"41efdc3b55c35cb3");
            when 10606304 => data <= (x"36da06af4effab6a", x"b21cd0480739f8ba", x"f4858f510abcd179", x"ab768b941088e2d7", x"e739116345b3e5b2", x"b77e6498e4219896", x"281b97689205c0a0", x"888cb45c6497aaca");
            when 14007221 => data <= (x"6f4b105aea29a3e9", x"fd15dbc17a7d6d5d", x"cf34aa0e152f32d5", x"95a6b9823ebdb56a", x"6f6093a6dcc093f6", x"796a74d80bfed780", x"1d58200984700eb2", x"3e5027c335427935");
            when 33659410 => data <= (x"b016bd435ab73d51", x"6b8136be85cc9836", x"3aa4a1839122a1d5", x"475160c68eb2c96f", x"73950ab80b5f6b77", x"6ea018920be37b4b", x"9d269fa8e20fa8b2", x"dd585ccd4d13b5fa");
            when 11199095 => data <= (x"97ea8f0afc77fea2", x"a5dae21227e1c1bc", x"bd3d314c84156be1", x"50749c6977d791ea", x"8fb7e4252ebae223", x"4cf1e5bb5c31f0c5", x"a1cf3d150eea4b95", x"5fa1966f28a9828a");
            when 3735038 => data <= (x"4aeed90065d3635b", x"d060837dfb1025ce", x"1c9b17b476275109", x"0645a2cfcaf7ae6f", x"a6db88d43a816b3b", x"711c0a12d0274ba5", x"7c47ad68e3fdfcd3", x"68a9cbf90511c859");
            when 9446162 => data <= (x"9d3e2e8dff632a29", x"1283d4e2348c1fdb", x"4d73a31513faeb25", x"a7fb1da59dc37bb4", x"6d8ec509c03fef35", x"475d1a29267df31a", x"bc36a86c53ff9b11", x"583940c44cec5e34");
            when 7008306 => data <= (x"e95665813dcdcb64", x"74b24d0199d66c32", x"429e1c69ea58c2e1", x"0503a40a8affa96c", x"75e06302bf310fe2", x"c2a0e88153a07b54", x"8e560687e6c791e2", x"93cb800f189cbc94");
            when 14098043 => data <= (x"04d687183620c5cc", x"32c1cb50dacd60d3", x"1c9ebff0145921ca", x"863af17d6dc037ac", x"0c76e6ee431e6d8c", x"d36b9eb6ceedb913", x"8db07a517050454c", x"6c950f6572ddf14c");
            when 23781821 => data <= (x"11fa836dcea9ab87", x"8ad97a4a2c46ca9e", x"64f3caed94d48b8a", x"d09502c2417d838d", x"3b2cc0ae130ec508", x"84184866c302503c", x"f6bc7260aa504dc9", x"b4185e36d3549f5a");
            when 22145944 => data <= (x"a6e9310a78a2e3e3", x"94d9df70df0016b6", x"5cecf176da09fe3d", x"8b991dd5652fc271", x"af7e9b3cb70c96db", x"4d0293182cf69241", x"bde53b88d9415994", x"b883dfad5878225f");
            when 23593361 => data <= (x"3971f75c483a7423", x"3960a748cf25acc0", x"4deb16b75f8b694e", x"0d6eccbb10820a7f", x"e718869f4a19c54d", x"c8965ed2293376d1", x"ad674cd60a792344", x"2fec19835d4ea411");
            when 14438634 => data <= (x"efb5502a54e7eb26", x"c874609159652eae", x"54e8ed7b6e16266b", x"8d0347def11b46c1", x"8b27d6fe106901fd", x"3df82013050706a1", x"a70a8125bb6c5866", x"cf706e2e60a0b9e8");
            when 7981572 => data <= (x"bd5fd79afd569ee7", x"6bc4b4bdd75e0054", x"2736dc80568cf5a2", x"bba34bcce9da19d2", x"e68acb5074a05ecc", x"e2c89256015c433a", x"aede865f3ffda626", x"6677738c0f289f9d");
            when 25706961 => data <= (x"64eca10c2d182b16", x"36c85d848d5a8143", x"2986c97fd97bd233", x"f011f2e3dad14283", x"2f1a11047fb0c0ab", x"6ae19345190cf663", x"6b8c8d61091023b3", x"6b6a44e6b710c720");
            when 18646475 => data <= (x"3d2e36043fe61808", x"b84aca7f25536c66", x"c3c01d4599af3f3a", x"00ca9430d8a2ba72", x"e4b89e0c3c63d7ec", x"11d85f53d83e22b2", x"9175f2f1d11855e0", x"8264f464573a3de1");
            when 8516229 => data <= (x"ae3f532871a1a754", x"10ea38bb4a8ff71a", x"f20e70348d4e81f2", x"cce4dfcbef798985", x"08a07c40a3b97c94", x"8bd45937717fa2c0", x"0520d27e0054a381", x"41c2b1bc46368efa");
            when 16881445 => data <= (x"7ad275b2d1b0959e", x"1b2ce43cd0816cdd", x"24187839cbda1bfd", x"8980b3183aa89f18", x"b29b53205883d30c", x"0d69cb80d831851e", x"94ab1749589ecde8", x"c4a75a2dded55c47");
            when 27665056 => data <= (x"993cec8fcc59876a", x"c8746fbbeedb451d", x"916c2d6f4ac44de5", x"9829f55db8ba0ade", x"25e48a7bbffa0f5a", x"b56d3c1d421e6f9a", x"7e279decf5588942", x"8ded26823d4ff7bd");
            when 27951784 => data <= (x"8ad9036c521ddd44", x"280df8152dfeb75c", x"16e7bfb662e3fc3c", x"54b5a13fe19dc15f", x"b119028c48d29de4", x"726918777ccb988e", x"9f60bfe686e56b11", x"b885c5f15374c098");
            when 15754255 => data <= (x"4b509e16cb905125", x"acc06348a0bab1e1", x"1719e80989a44885", x"757397f31ef4dee5", x"0c2d9b26d365f084", x"cae9abce82afb1a3", x"d45fb62ac145a468", x"7f5814acf5cb3f39");
            when 22723137 => data <= (x"4aab52f2de6e1a2b", x"b8b10155c51085c4", x"f1f0534a917f36ac", x"44c060e01affbd3a", x"b4ec5dd418ea093d", x"d5a0f063cde7a8ae", x"25324936840809cf", x"594095fbac38c1eb");
            when 20950049 => data <= (x"4a55747fae1a6890", x"3994e2b691aa5759", x"6abd0af5eb3aba57", x"3d20a1ccfb2d1ec1", x"094cee8d2fd5a76d", x"4e5611e45e2e6197", x"324b46fc135cc76c", x"60ea1cded6a59b3e");
            when 19355068 => data <= (x"80b1bde2ae6e3c8a", x"67c652bfe2e39ea4", x"85a8943f229ae618", x"1d37efb2925b511a", x"dc2d012e1cd36435", x"ab45fbe22027c92c", x"a0d1f7803cb2f4e0", x"e4964fb8f5b2a85b");
            when 30976215 => data <= (x"3be35c7c1a60933a", x"e0714379301dd143", x"62e409731c14d419", x"376dbe7af5a599ce", x"ce0b2fc17ccecf9a", x"4d2039a859a3e90a", x"063a0d0d59fb05e9", x"b22e7fb6aded194d");
            when 25459519 => data <= (x"635cf882240d0a6f", x"ddf46ecb8fda296c", x"5cdd38742aa3fce7", x"f374a7dee009c266", x"e2047bff8087452b", x"bbe976bc9a98064a", x"e72e20c4077297bc", x"e23febc6cc5fbfbb");
            when 20469593 => data <= (x"a0ae23cebdf2b93a", x"c74c4a19c013d354", x"0abe8ef014e2ee9c", x"a009fff1f2a6a947", x"45be8ffc34d0c68a", x"441b57b1c700fdea", x"f61049c0fc6788b0", x"b8a0982d9e0f75f7");
            when 12959388 => data <= (x"e5da6f0be905ab58", x"ed5cc59c3d72b17b", x"4104bacd8f87f2e6", x"22e11ef1b272acd0", x"e5854d5a1e2b0753", x"09ce6b1d7598610b", x"3fc8608518874ce7", x"9b6d90af479be22d");
            when 27997334 => data <= (x"0018a867ab47b28d", x"6b2c7434cde9fdf3", x"aa60832df5b683a8", x"8a568e75bcd2c2f5", x"1befafb4fee88904", x"e88f3e51ad4ae62a", x"a7ccfe63d99fb17c", x"f8ab8b573748e784");
            when 17312483 => data <= (x"ea0806a6085d96eb", x"3f417d980fe4cb42", x"cb77f222b686942a", x"92c69aad9368834a", x"09974e3b93ddabb8", x"1d82938e66ece735", x"feed8fe9a5c7239c", x"717ce17f59b58ac7");
            when 25488402 => data <= (x"92d0d9880a88838d", x"99edd78c96dbbbe5", x"419482bcc8178e2c", x"05da687bd38c052a", x"d806fa708159c4d8", x"55859bd31b2c5fb5", x"8ccb2c7e30dd42df", x"7ad9a4b37c4583ee");
            when 21210492 => data <= (x"ec63068488b2900c", x"a3becc987a92e2fa", x"c2865893e1456904", x"9c762fc79bd06a88", x"acf643fec7d8606d", x"1bf3f386d183acd8", x"e7a9bc96b7cac295", x"d25f34439dcfa988");
            when 10475769 => data <= (x"8653c87cb35593d9", x"fa39c163fc8e5093", x"13651c4f89687e28", x"9109b5eed6e57259", x"3928fa4802a7ce0b", x"c9e82111bc1a64d8", x"5704b9dae3108c0d", x"0224d70afe3da149");
            when 14709327 => data <= (x"ebf8717a013d317d", x"6fbe247e58e01570", x"ea13f50a9810428b", x"35ffeba30c23e791", x"b94a713bd649cbcd", x"a4abf92b833d07fa", x"e23f219b98896d3e", x"cb14059c68d2b905");
            when 27653882 => data <= (x"f46a46b7f8fec1d2", x"b65540b62eeb93b0", x"1c7b2af4d0ae23e7", x"993456e288ef0db7", x"d252e314cbe327d1", x"d2eb1870ca7bfac8", x"9dad578252fb103b", x"1100e577af612173");
            when 30371228 => data <= (x"d89f471af443e605", x"5994b0ea1a392639", x"c7c25af18412e8d5", x"952c5d1954338f6d", x"865d66eb6320c943", x"5708ee6a7581497f", x"1a95720d471c897a", x"b4f934d8f6ac551f");
            when 5504428 => data <= (x"be0fb2963f8134c5", x"3f1cce2e422e9016", x"bf4c7833bcadc8a1", x"ce4fff34ccafaa08", x"ba30add1d058d9e4", x"a68c6d48e5b63f74", x"04f9af60bcf0f053", x"6ff5e2615b1a21bb");
            when 32413123 => data <= (x"8912423c8e1b28c2", x"62096bb113a5ce0b", x"eb9cf5bddb0fa94b", x"52e72b35e0ce4e79", x"c6ce5069a89b9c0c", x"4c6d42071bacd1b2", x"dce755cefb5f0291", x"661d134978f0c378");
            when 19400514 => data <= (x"1cd801bf67060a7b", x"fcec7890876dce82", x"d08de503dd781912", x"67efcbaa779c20e9", x"377ad7fb7a4c03f2", x"2d13843558e5f6eb", x"a14575ca074b92ef", x"d5f144e97de3bed0");
            when 26908773 => data <= (x"02ce3110263144d7", x"aa91cd0f09ea70ea", x"b20d424e84b4a041", x"7f79f9a3bf3f2f87", x"3d3afca514958f7c", x"cc9cfd35ddacd545", x"c0639f9e057deb5d", x"7b07f149a81e25bc");
            when 30602170 => data <= (x"77da2a6f1f9671a8", x"6361269b48717d4b", x"8a832565738e16b2", x"fef3c8a9eda12de0", x"f74dc64e3810d922", x"b0b70447ed6eab42", x"dd6687739dda1b9e", x"0c216833570d95df");
            when 1337851 => data <= (x"5bc4195c720d75b2", x"386098059df6740d", x"2922f551af4b4997", x"07dec0f8d9a28917", x"68a5e7e39f3d023b", x"fd7f65254523e058", x"b77c75d92de197e5", x"fa8565829f0ab8b6");
            when 21336418 => data <= (x"0c04da6a547a840c", x"9003b9af13cb1724", x"ab09725503aebf17", x"32170ea2630123d6", x"0e52451d5978df1d", x"016b5aa80ae158b4", x"70f5eb101e3fe17c", x"dcd65e83480de5b9");
            when 24244990 => data <= (x"5e6d5de0d7559b9d", x"617ff0e940e1a17d", x"3e407fcdc95d0ca1", x"4beacbcf7209c5ab", x"cf13f676f706d595", x"0a58158983bab4d3", x"eb189a26168c9b83", x"0fbb972ec5ea0c56");
            when 28840206 => data <= (x"921a375e55f4d6b5", x"42493e6989bbc628", x"80d1ca09b9fe064f", x"df32c5b1c0b244b3", x"f5a8ed26999f0272", x"18df19cbdc910a72", x"4f481dedeb00c387", x"dab4454a90c8b2b5");
            when 1159586 => data <= (x"de026786a0798ab2", x"139608f4ac5ef2ba", x"0c77bb02d68d4880", x"c78619fe2e8e43dc", x"617c8813657fbbb8", x"4c955d4584a91d9b", x"8f5fc16a162b1c68", x"c21f687b0a2df3cc");
            when 32465526 => data <= (x"bb5cdb8b3c211bc4", x"c11d914ada92ed86", x"d9d647a080c7fad9", x"7621035c38fc90e4", x"d407c20b0851afa6", x"aa9d8fafb9a8e88c", x"49cb5e5fd60673c1", x"f4256878ad3f3702");
            when 27452501 => data <= (x"4a6229751925e9f2", x"3c1c8b2f50653774", x"e9093b5c6440f397", x"0696d8e27476b5eb", x"8054c139f944e8fa", x"4046e21bcd03aaa2", x"cd79432948f4ab94", x"34727af5018bb74b");
            when 7797297 => data <= (x"8edb46487b452134", x"d2bbe1ce8ac3be2b", x"3559a3d6d73e3ffd", x"dfb76c0dc63fdb6b", x"127525731a8c3e27", x"df8b503c9fdf60f6", x"e0e60fc1ff08b210", x"a9dd0701c482d877");
            when 20203285 => data <= (x"d54935c463fc765a", x"27da218eaa435da3", x"5833e673b34c5781", x"371219ab4d9b181b", x"9622ecca8c50bee4", x"e0f494b6248b079c", x"60cf3f939acd6c27", x"e9fd4a7c3acefa55");
            when 13522208 => data <= (x"62ca2513b8a84571", x"62ccb5a7bb13afea", x"ae802feebc173b23", x"c5923f1ec3ee6e11", x"b83379c7ce62318e", x"be7d58194e6a2634", x"a99cf9555c8cdc18", x"04ce33754fd3c9d9");
            when 10227518 => data <= (x"be89774e6172b93b", x"186a710da429f9b8", x"9eea261c6753918f", x"ad9f88ca0603de25", x"2bd158490dd08415", x"7e49d6084da9d02b", x"1038f43d0c88227f", x"fb59e450d354fa07");
            when 8610988 => data <= (x"c3246931a9473ae8", x"211ce84082380b5f", x"624c9bb115425567", x"b346db489c848768", x"2cbae0706b60672a", x"84e492096a23f919", x"4e34c3307dbdcbee", x"881962cf48d00e6e");
            when 6536971 => data <= (x"c060caac752537e7", x"d09f7bf6d87ca3ec", x"f2105046cc0cf8bf", x"9e2735fbe7e9b64a", x"9647ba3b545be956", x"0434f537daa56d67", x"654da5c787bbcb1f", x"4de610992215ab9c");
            when 33448778 => data <= (x"8b83f8f71518ae47", x"8b97f40ad7c03acf", x"2b2e8673d696d09b", x"4db9f1bbd426eeb5", x"abc80cbf84e74a76", x"1eb31b2984afa75e", x"979ded580baa6001", x"83f9bc26da4af0b2");
            when 18335929 => data <= (x"3073a1137a7bac31", x"b4cb1a399afa81ed", x"837163271d5e0808", x"5043d244799075af", x"37ec669d774c14dd", x"530d6cff6f6b25f9", x"f0d8aff9a19fa780", x"1f83af1a20243eb5");
            when 1902785 => data <= (x"91ba87f8374541f9", x"939c74bf8dbe47e5", x"959aacfb11132d11", x"95a68833ebcf10c6", x"c92d9ff6ec823272", x"033131167eeadde0", x"6c13eaa21b427ec0", x"7c43e7ef1f76f6e6");
            when 1951632 => data <= (x"db5be067809fc897", x"a507b5d10618680b", x"5a9b2f099e260969", x"21c430d0d0c02993", x"e556a5413d5ce746", x"a4e5a11d860f0361", x"b25f9988fbe2f7b0", x"2374bd924f16dd68");
            when 15330188 => data <= (x"4feb44cd663c43a3", x"9167d1aa4e797a18", x"50c7a149a5de5099", x"d52eb907e189848b", x"b7fa819530906805", x"fdca3904388f71fc", x"594ec277d8d81e5b", x"571f7d70ee03a367");
            when 11173150 => data <= (x"dde53b1b0ebbcf07", x"3c204ed4d8490541", x"9f65c37ceae6e7d6", x"11c2006b9ac8f135", x"9458c49a087105aa", x"8bd7d7f23a9acde3", x"19e137b1862657b3", x"c67491bf47e5b718");
            when 32876154 => data <= (x"6163cfcb5988a006", x"4c22fb7e50fc3c62", x"1079d0aa48766154", x"5725542e2115ead9", x"8884898607045bcd", x"eac10ca5690e033d", x"4e1798799201615d", x"90046508fc41f2cd");
            when 28993663 => data <= (x"2ee1a295f87c3764", x"08fdf5c176bec832", x"13d77398b0d22cf5", x"6f09d5e39d82f033", x"8f0859773cff2b93", x"f9c991807e9be5ba", x"af63533f88160109", x"3116b5b4a0881d94");
            when 1961442 => data <= (x"a406768dd0bdad69", x"891bafcb426f1d10", x"4747ef0149fa7853", x"2bb2b9c7cd9e4c96", x"6462bebd71409b6d", x"e5be9d0690983148", x"0045a737b69ac6c7", x"2b73acc32068c303");
            when 667533 => data <= (x"d27dda04eb2193fa", x"40d51200030cfff4", x"2cdc088cb4eccfd4", x"56f518c400e37d8d", x"8ac777ded7efcada", x"cd58dca2502f9980", x"5e53bbb4085943fe", x"2e003c497284f65b");
            when 29989081 => data <= (x"cdfee7c285df37a5", x"ebaf05367923ea58", x"831b3a2a496c0f42", x"6f064202cd47e0f6", x"788da280d9e1825b", x"4e95f0bfbdae623d", x"632f5f3c9ab0252c", x"3a197838b04bc83c");
            when 13710232 => data <= (x"5024533282551d32", x"683dc39a5a78727e", x"1dacc4cd66c1dfdb", x"b0951ff8ae551030", x"2092ea1b407516bd", x"830f28ce6cfcf057", x"dc860327a754f437", x"a210e54685b11709");
            when 6483826 => data <= (x"a138b62bfc26bec6", x"40b1c9ec4d87aeb8", x"e93669650416dfc1", x"c76e18c459642ec4", x"4d313d0b620c3d13", x"d1e0cf06dc3d81b7", x"b9922e6ecf983ae8", x"3b251f0ea93215f5");
            when 22827626 => data <= (x"e37004f43f6cad7e", x"8a52efcefeceedf2", x"f605007bc7a664e7", x"9325679be28a7d7f", x"81a4bc569e346d21", x"99d853095b3d6cd3", x"6cc6b0831e2c647a", x"e9ed49696028110e");
            when 4851046 => data <= (x"89b7ea456d866fe9", x"8f8d2ba931a3cf0d", x"1f70e3efeb3d18a9", x"22b93e4d6c33092f", x"df1b8f6bac9d4249", x"cb70b89ca8751f46", x"6c2a5652bd7c2f33", x"c70913f49c3a6df2");
            when 7196262 => data <= (x"14ebf44f421ef357", x"165f2f97a9dd4d80", x"0b156cab20f9bb24", x"b738214a0fa2cb8e", x"d4e2961c2548391b", x"1ef39feaeb06eeb9", x"b8e019f8ddf7577b", x"451467b0ddc1f120");
            when 4986653 => data <= (x"9d09d80dfe6e56bd", x"ba8006576fb85198", x"67e722210a506ea9", x"b3caec3f6f97924a", x"ef6f15cd8970406f", x"32bc074e9d798902", x"04e0795f3293a6c6", x"70132034f25e488e");
            when 1716194 => data <= (x"231ff70ef6f47562", x"53ef3c1758d81446", x"38aad8cfff5d5dcb", x"47ce0752480b3e84", x"2b79cf01a9929840", x"83e74eed51a8f654", x"5e79c763d060b3bc", x"8744cee9495b6526");
            when 4341011 => data <= (x"6e5fb9d102a2badb", x"8b6aa9148b1b9935", x"6ddb018458312850", x"3703f77cc5426fb3", x"ddf7fdb676d59215", x"89acdfef1e47bdb2", x"732b0aecc627cf05", x"b2c01e81b337228b");
            when 21556193 => data <= (x"f78c4ba43cc76c83", x"a3113e0c47244c63", x"19b13cc0a38da649", x"50621b2248270b1f", x"fefd39af67e35b9d", x"af0b5d710eba552a", x"7b854dba0f98eb9c", x"0af11512544edc6b");
            when 23667249 => data <= (x"d959da7e431bf2cc", x"a4716ec45319b469", x"c6798182ef6f0ab9", x"82f05a8d7eaa54e4", x"54f254dfda4dbdb7", x"041620471b6b5328", x"ac9e225b86d0861a", x"b0114147ed28e44e");
            when 33365930 => data <= (x"e9a5bdcdeb60d7cc", x"cf061e6163119290", x"46185fd2053cab39", x"df9e866a8923cd8f", x"0f79c4ba778a1d2d", x"2d766f748fa955aa", x"b02871fb6eca9417", x"fdd488f173ea7af3");
            when 10459594 => data <= (x"454be89e7080e988", x"3113522f619e8d3c", x"e65c118649b00ce0", x"3129a41e5c165a77", x"4ea81f9929a77180", x"26779b66672b42e4", x"968b9a652cca9e70", x"25c6051e62b71aa6");
            when 6705811 => data <= (x"d77094d83f2c8a6c", x"4ad1593a7b2757f9", x"1bd45f37fa58de42", x"fa005418cdb7f02c", x"cad0693b41f9533e", x"bd715ab5fde4109e", x"e712c34b261e3d3a", x"48d933c15b9949c0");
            when 11865106 => data <= (x"b2c6b4db30e2c125", x"60bcdc374b036d4a", x"f0151e55f454b771", x"17239bdca1177968", x"30f987d0d0692eba", x"e60b19c26df61799", x"3ecbf96cdda656c3", x"f49214d611bea596");
            when 33746458 => data <= (x"fd8ac6b55050d819", x"41915d3ea2aa6b52", x"bf2bb01676bfc21a", x"96dd79bebe447279", x"852f9a6c6886924e", x"3e8544e685cb92d6", x"efd489202be4798c", x"b5a4860387b0ec11");
            when 15815780 => data <= (x"2d6e9d87af00211a", x"aa2c687ee222e9ca", x"0b387a8648a4a845", x"3bec8404da39d638", x"183c3507d258a7b2", x"7ef61a1a67260c8d", x"fb5116e3172dec5f", x"c104bab8f3b95717");
            when 25893676 => data <= (x"281262c01e34e214", x"e1fd51d8cf137937", x"58b4b47603c7e6b9", x"e7a60e04a6c03b08", x"7f55093a37e7c061", x"80a2d457cf4bdfd1", x"d7616702be34ad7d", x"e1cd72094ddccb12");
            when 28797697 => data <= (x"4b3956e00c5abfde", x"3943de5a139729bf", x"dfb78adff7f57e18", x"61e3c4ca9081a366", x"028d54be3f15d754", x"f1a5d744d4fa8ab3", x"b269968975c3e940", x"a4722d801497ba0e");
            when 33598192 => data <= (x"dc6e5cdedea45f04", x"54c4eae09dcb8d62", x"66f1e0a5058f0a47", x"1d48ff46fa2307f7", x"8089474be7ce9bdc", x"f2808baa73a73e2a", x"7e28e19e0dc56307", x"f65f3a0d9de9e700");
            when 28813582 => data <= (x"afe7feb966cdf31e", x"6a296329cb2a3aec", x"cb134997186bea16", x"8a4d17ebc2b7b5fe", x"5ce673a321f0c1d1", x"6f2f0167a8e6294b", x"dbeab96ccce00787", x"77871259768290aa");
            when 8539700 => data <= (x"ff536babc1684f83", x"5da567a8ca2142bf", x"5801c49796c4d600", x"f15c6f014f4bf02a", x"31a0447986c94a24", x"2edee198a0a94e5e", x"b643dcebd676d545", x"99e0182744e61e30");
            when 10158232 => data <= (x"a244fa4e151e6e94", x"8d35e352c1fdb0ad", x"8696a7cae187ae7f", x"951c3472755862ee", x"4edd8a59fd70610a", x"de6feb5b5b2c243b", x"6461c3d8285fe445", x"90bf4f70936a48f1");
            when 6085427 => data <= (x"135a5d9afbf9efa8", x"f8eca8671e3910ea", x"83b2da2b7d24a4ad", x"84115ac02693959e", x"03ebaf673f0f666b", x"fba6f26d5e8e46d2", x"9ae6bc5ecdf64357", x"0de891a697f07952");
            when 14876094 => data <= (x"3bc7cf6d393da20f", x"0e6d738af1492e75", x"76aaef2c1f9c8b03", x"e62312c741ce18e7", x"70cc6f6e5c9cd3b0", x"8eb6d9f396f11531", x"9218289653296c81", x"6e916c2ef047e764");
            when 23964560 => data <= (x"d08357647efd05de", x"79211686b0c26315", x"4b0c4665f8ed6398", x"e283ed94c52ff6fc", x"e90a3437abaae84d", x"70162542544c667d", x"69bac10234a126b9", x"2f36d946616f0697");
            when 24565825 => data <= (x"c79796dd29da275b", x"4a55e1c8eea340c3", x"91c99db325e9fdb1", x"a7788ba540076f97", x"41748b1416e13bc5", x"4082cc0408f7a3bc", x"0abf8d0e76d4e82e", x"1ea2c81716e44f60");
            when 12084924 => data <= (x"c84f85322c0e7adf", x"f7b2e1930c55e704", x"72c33fb0b21c98d1", x"48a960a5c82f5477", x"d781cc2e322725b8", x"9cf89a29a675fc71", x"1835b69b73fc324c", x"b03cb08e27d9100c");
            when 32232175 => data <= (x"bce8559fffa885df", x"48808b5c3ecc615b", x"74644c51780b9679", x"49dff7164a96e66c", x"6ccafc625af7b649", x"01ff6b1069c232cd", x"afb4a7240974f5ea", x"6f225df330190ec5");
            when 4695226 => data <= (x"3a60642fdcf1f8bc", x"b54401edee626ae9", x"c4939cea48341548", x"b4bc48e291972965", x"f563a4d6cd9ad440", x"569f79d83160406d", x"dbbbe595422dcd96", x"afce4203917ed3f1");
            when 4133299 => data <= (x"50cc6b9568af8aef", x"bbee3cd6387ccec9", x"cbc8dd09701dfd95", x"61b4537ff4054ffc", x"c60ed40d8ea1e90d", x"94af75dd41ca5d3d", x"5d9b1cd97fbd10d9", x"c0b7f4176ba29979");
            when 28870348 => data <= (x"29ada92305047a75", x"d2feab25da538d56", x"6ca08512f441e175", x"6d15818e793511c2", x"09e84ea026944c61", x"117257f28db5fb68", x"5533c38294b66c4c", x"695fc54dc4c982df");
            when 33418794 => data <= (x"2a238eb28a5677a8", x"1b42219f82301d3e", x"707cadb56dc80871", x"a31ac104d996975a", x"5f6fd87e119228c0", x"0d96ea617bc99520", x"2dbbcb910eb7fbae", x"999ceacac597ee8a");
            when 28098723 => data <= (x"9d9e7353f3b5980d", x"3483d3c29ed07e86", x"f243973671e9c770", x"6c71ef40afe0fd81", x"d3e2de57e5247f5f", x"dc38540295e9a396", x"9f40bcdfc2ea2584", x"3c6081434155e8d4");
            when 24576341 => data <= (x"112cb111b620caf5", x"21bf824b864af217", x"4325a3f5b782cc9a", x"df082a5223de4886", x"c04032f8877b5004", x"eb1b6b238feba07e", x"5a27691824cc5342", x"7757777d9e878a27");
            when 22459859 => data <= (x"ca61a2b8893c94a8", x"8bc0753dfb214aeb", x"f1eb25c63540af75", x"1459a5260862bd21", x"0122664f27769c24", x"69023c12a35be602", x"8f2ed701cbfc3331", x"728806a0ae96d51c");
            when 20193975 => data <= (x"268086e28ca889c2", x"f6d99fbb3dae5dc2", x"9ada050ee27a6133", x"b98d00ae423ecea7", x"3b4dc5836302b4b9", x"31f57328057b25fe", x"c6ef4155cda19c2c", x"b8cf25468fa6ab24");
            when 28305206 => data <= (x"9ab92d060390530a", x"4fcf79a595fba2a6", x"4ea27223b21641f4", x"4abc0d939ee8cda7", x"33ae376e46220785", x"b906c55fd4d31ac4", x"b4581075e1169374", x"c2bfe155318bd060");
            when 29106350 => data <= (x"fae4f50568dcbec0", x"46bd21f74ce5f290", x"5ea19ac954f7272c", x"269dae2c2acffbc9", x"701a5adfb7594cb1", x"0a878cb36dbf8e21", x"acf17f90b4e600a3", x"f722b810a2a25ace");
            when 18370087 => data <= (x"073314e11c38f5e5", x"6c8bdd0d1d6de6ba", x"6bbe97b8af438251", x"8e4359266a7b9d9c", x"a0f0efec82d85235", x"8871de598ebb861e", x"e3163270a69b95c9", x"3e74ba525d9f7d0d");
            when 16821052 => data <= (x"721ca984a357c773", x"c354e6b6ee775734", x"e4a284d67d5d3801", x"ad48ce63976cd2e0", x"5c0959b9fdfe9b7e", x"c7c46f89696e4c7f", x"f7d180c95fad76c4", x"34b70dc541f6cf92");
            when 12656289 => data <= (x"db825727cb7ac88c", x"41a7d34bfe160a85", x"665a0327e94df709", x"3f2a9237080a3b67", x"0211e097f0e28bf7", x"071216a9076d89ed", x"33d548e262b3d266", x"f8311bc7b27a7c48");
            when 18121613 => data <= (x"8aed1e19d2732a5a", x"6985767413ec4da6", x"835112c499509ee3", x"f935d48a0f1f30b0", x"e1e4f01fb15c10b5", x"d3e40510229486b1", x"50c1483c68b7f28b", x"603c35993961942b");
            when 18790217 => data <= (x"10a8e0edeed4698c", x"7120b1ab095dc7c2", x"89f85c91d73d2b43", x"03b861d504f75a47", x"5faeedaf26942d8a", x"8add725850243918", x"16cc7ffce888a268", x"cae9cdacaf3f9a37");
            when 29108687 => data <= (x"c95256d611a959ca", x"0bffe097cede8d7e", x"c72db3ab5f2d2d84", x"0571d97d16860203", x"4456f57ac63f08e9", x"d5ea8b862ef6ea64", x"89affa2ccda7183c", x"35b9a88bfaec1535");
            when 25328090 => data <= (x"583ef810ef110012", x"0e52facc4c4be025", x"31a97c7b398bf2fd", x"ac5bcfd781444e08", x"54c085ea8884b637", x"bbf8fcd6c101db47", x"a490e7132c6d04d3", x"40283acb0f56261e");
            when 25927209 => data <= (x"81f0e02176483b0e", x"6bb8097d6fae1ab3", x"be96020f71f868e2", x"183e262d02df80e1", x"cd90071c20458f36", x"e2b7179201cc9691", x"2ef9cd86e190f30f", x"458dccec11c423fd");
            when 14797453 => data <= (x"0c3846d126ab7641", x"38328da1eb5c027c", x"554f4ac771cfa61b", x"c39bdf3469d557ba", x"27661b9df0315261", x"451bd78f2042eee7", x"ba153e7acb3c2846", x"d0d3094f182804b2");
            when 16498436 => data <= (x"4df0f96319595145", x"679ec669975f9fb5", x"3bb269ffb44c27e3", x"ca8c5de097d2db56", x"a69394ea335d33a3", x"3ffd9c0c71049e6b", x"f64ba293885ccea6", x"7435a65042d7e163");
            when 20147063 => data <= (x"e679b4c7692b2ce3", x"02391f1ac3817f61", x"6e63ed7642f2b8d8", x"bfd1b09554fd45e1", x"88260bbb429b0f40", x"bce53a6ba8452549", x"b75cafbe185ee514", x"78eb26bfd7884cca");
            when 5779686 => data <= (x"21ca2af05627d2b5", x"ff586d831bd0c548", x"b74be66fc493b6cb", x"d6e5b492ca2f3732", x"799affdb92d72bc4", x"6e9361b0bf948622", x"cd0663a1596b7a68", x"d4141855f641b576");
            when 26042245 => data <= (x"048f4a9543d9897a", x"0837356633be2643", x"ec1e185db40f9626", x"7fd59bcd9217d2a6", x"a87a0927a4b43f67", x"e837ba5ee7607cf0", x"b1f26a43f701bfcf", x"79adccedbc07e590");
            when 12005679 => data <= (x"a77af434183065b4", x"44409ea72b514685", x"8b44d4f230c72cbd", x"37c08b48f22e5d19", x"90b08a380e1333e9", x"97233cc9c03004da", x"0583a0f003635bd4", x"6ddbb55f69509893");
            when 5337899 => data <= (x"8d0811c9b16d6ad3", x"f7900c26bb18b2c0", x"a0b8aca5da5e95aa", x"74f1de21a7f0a3f9", x"4ac96d0f9550b1ae", x"39b30005489db817", x"afb1fe9b7904d101", x"d3d0223ff1ca7f83");
            when 17539468 => data <= (x"4357aa2cb26b1225", x"503a9bcdadeede45", x"216fb86849bde671", x"5f5ee5824be65f88", x"a211cb680fd3d7d5", x"a823ecedbbfb33bb", x"ddd74d8df587f31e", x"655ea5ff52a76e2f");
            when 16309006 => data <= (x"03f07d6a9cb29135", x"ba8742a66478b1fe", x"faf6badd7ea22885", x"b6ed9f9b1f8cbd2b", x"0d56fef24d865ce3", x"377fa61970acb479", x"f6000d8df9f508e9", x"bfe06bffdfb06ce9");
            when 29519409 => data <= (x"e680c26129793c43", x"7d6e06d7a1fceb69", x"c4ae5533b13deb87", x"3748b9e43f03c919", x"4961b6a5101c439e", x"c3a207e8f592bf96", x"473f6898eb36b28b", x"e1bda620ec1bc9be");
            when 14172017 => data <= (x"5e3999e3f4f45704", x"4168af5b631358c8", x"93cc3f2c0f403274", x"eb4b4fd43d85d911", x"26c3046a5379fff3", x"f9a561d977f864d3", x"2aafbdee47743d42", x"c59d41d0610ae18f");
            when 20376989 => data <= (x"e35516b1c5b96fb9", x"079f97664d1b94d1", x"b6de458c9880207c", x"ab74e9f81402d0d3", x"983a19d42651dfc5", x"72645a5213b97519", x"fc90e3cb4d560ce2", x"f7d4be13d0b86f3c");
            when 20885932 => data <= (x"7f608213daa9b9f3", x"790baa5369df3692", x"10dfaa55e20df51a", x"a5bcf34ab4be87a5", x"441cf81892bd80ad", x"7d7b6beb02acc2e4", x"24ec3a9ffcb3d62f", x"afe77496e5c7e2ae");
            when 17217932 => data <= (x"fc597957c2b5f302", x"aa98160bec4f68df", x"0996b88c24fc88fb", x"b1c3e8c435707b6c", x"a4aa7f1b16da6814", x"b9cc332fc917996e", x"0b7bd4bcefccdc1d", x"3bd241c60f061b5c");
            when 19386466 => data <= (x"999c2a4e8b8035a2", x"8f3beef066fc21b4", x"53e30446d58cd6c2", x"2ed6ce1517b5f93c", x"35d2725a4d6eadb6", x"f816741336e9d5bb", x"127a387cc706991c", x"5fc814d2774e480b");
            when 19819000 => data <= (x"c599457d5ab65b8c", x"bcd451a70edf4932", x"1e0af40880b5e2ba", x"36c7c5dc7f185169", x"b6cdc3737b841e82", x"88744b5f9f06253c", x"5bc16ffd2f3a69ce", x"2530e6e475efa571");
            when 14642441 => data <= (x"f4960e2e7373f35c", x"6be8134925a99666", x"50106c836bba73b6", x"3fa577c2131734b0", x"712e3dfb6d13f8df", x"e102513edd58cc02", x"293e5b8657ba1490", x"4a99142d8a396d69");
            when 29512557 => data <= (x"c875fe2e5698620b", x"b4f9e59227051ab0", x"e5b6d9217578e8f9", x"62e22c07d4dcce5f", x"edc7cf21b4a36cad", x"e9005ab42b09fd40", x"7a73234ce46c8471", x"217102da4ed35b7d");
            when 10401145 => data <= (x"9f45a5d96c927cbb", x"81fc89181e799f52", x"4f1062a00095f992", x"8c15f5a05f2a7377", x"c1eeb6311bd8a07b", x"918a479958d4bc06", x"c9858fe2cdf04d11", x"f67bb4ea8251092d");
            when 9747545 => data <= (x"c8d65f9c36797821", x"ff45eb27b83d2f7e", x"ce2843b318b46bd6", x"95109dfef11f35fd", x"e38060088b8ba9d0", x"97a677ad6e0832c4", x"201fdd186e4001ec", x"9f56514ed3338942");
            when 3145349 => data <= (x"927437e23d3d5968", x"50a57aa31da77c18", x"7cabeec0633e7eec", x"a82a87401fefb408", x"f557243fa506cde9", x"525e37a0bbb26de9", x"98d3f02437385d05", x"e7cb954f9f95b51b");
            when 5743082 => data <= (x"0edac375fc626ed6", x"66f5cd948e9dd9af", x"2378c2e0c737d415", x"899d3c09dc95bbba", x"061e10303a8bfc33", x"de8d037d5a51ad1e", x"d7d99ccc3fb5e15a", x"5d9df00857bd14f3");
            when 23772670 => data <= (x"2990afbf62f704f0", x"c94879dc5025bcf5", x"3c38f40de17264a3", x"23702b655ce3a357", x"d2f6ee9269059fbc", x"95e3a2ced7c47b02", x"37588109fda8f548", x"430b9306bc0c8b88");
            when 17702693 => data <= (x"97ad35bcf24efba6", x"de8952ab1381c434", x"7ae9fa5ae668a166", x"d2c7ac793594805b", x"1f84945142f9d85d", x"7cb34ea0e2ab6d45", x"6d113bd9c17cd26e", x"df7c98ce86a2caeb");
            when 6758021 => data <= (x"71e5fbd559841771", x"30b46f84118f0e2b", x"f696d9a08f386ded", x"0a72d1fa3281e1df", x"c279482277fc104b", x"eab74705009a588c", x"8695a08f90ec5632", x"83606d0a260eb7dc");
            when 24865349 => data <= (x"b1d816b4886b4ec6", x"b424133ea663ca0e", x"9a7650a13fcfe7e2", x"a7840e4abbac3e7b", x"d637959b7f6c4e2d", x"9183a9106235e7ce", x"dd5e25cc8fd9199d", x"89a6122f4c17415c");
            when 1711731 => data <= (x"c9d5fbcf3e45d85a", x"5f0a289d52674dec", x"d4497caa002fa5f4", x"9dbbfeaa8ca93144", x"07b211c3f94345f8", x"50e4c5e101d9002d", x"700701fefad64606", x"551db1fba51dd663");
            when 10065762 => data <= (x"c1fa5326c7bd6a19", x"56803554b640ecf0", x"29a25cb2d0b496a4", x"fc0ee94bfd2ad8fb", x"351fc101516b04d2", x"4a8680e6b5abb43c", x"fb9758d3cd478361", x"8eef0281438bddea");
            when 22117431 => data <= (x"110ea0ac859b8442", x"7c347cb5b9b2965f", x"04c2ebf8d397df4e", x"2e7d17194f40bb17", x"55f7e5ddee52d89b", x"6b35b2d32ef2924f", x"746ffa4825ba9d6e", x"fa9f7b2adb22546b");
            when 30876189 => data <= (x"7c00872f55f34151", x"c18f5b3f844a348e", x"0e0e223f184de9ce", x"6bf03e4241cbfae2", x"949683c1fddec290", x"1a01b5896d25d33e", x"5335847a8677be07", x"8cb555b234d5005f");
            when 19708392 => data <= (x"d9e177eb0ba87f7b", x"e37d0156abf80a21", x"39a491c8b9382fc3", x"2fa83836376b902b", x"5a8f1fd96ff5d99d", x"8a40594712012652", x"5a0a80c8d1928cb2", x"72b82b028e4eec48");
            when 24504848 => data <= (x"7d98573011050ccd", x"8fd131f169eb8a3d", x"747fd1c6d1a50d01", x"e2fa09fbc46823dd", x"0e22cb94294640c9", x"9b375c0f30b6e18b", x"b4b0419b3b74a612", x"a0135965deadee31");
            when 13451210 => data <= (x"8e12810932287ac1", x"adee816838766019", x"b0458e3996539103", x"69a757c3f7fb61d6", x"dd18c3a35f7ebc47", x"23c54d2049500336", x"612d5186267768bc", x"aedd06bff383f5bb");
            when 1191910 => data <= (x"51d391c5a29a2a19", x"13133e1e5e1271b5", x"6ae77b0d520ce84a", x"535071ed6b1977a1", x"88adcd820216fb81", x"2434214d9e73eae8", x"ca2a05755619cb4e", x"8e290132950d63c9");
            when 17496619 => data <= (x"557a25a72d30633e", x"efad5a46179ec32d", x"5235d1230be42b99", x"64191a8cc9b56e54", x"30a8b73331fd9004", x"a10a7fe7063c1833", x"f1056e5e9f7dd298", x"bbf29e6d584585ab");
            when 12555989 => data <= (x"8cf71697fd0a4198", x"cbc4b54055419066", x"21fa641d2fca5756", x"e2e75f86ab88a314", x"62cce13299978044", x"841446dd03c892a0", x"b92390f85bd02ee0", x"34fc1c8a8584658d");
            when 23720836 => data <= (x"e9508b0914bef336", x"de3c6cfd3580fe6c", x"3d1dcbb2d451eeb3", x"cf822f8251c5392f", x"a3b1f18c8a13ab2c", x"eb0476eba64bd542", x"6ecdbff3a069f616", x"44c69f90b2455e41");
            when 29522286 => data <= (x"1cdfd2c5aceb8d97", x"2d757965e4a65828", x"a7ba3e564166d6d0", x"ef16f425b19e0fc3", x"bde5e41e32efe2e0", x"dcf966f1230f45bb", x"4c2436115609179b", x"ff7ba32de0cdd361");
            when 15303102 => data <= (x"3a80838e497600ea", x"38b654c3e6a1424a", x"4bc43efb641ce13e", x"286e01c9f2716b5d", x"e34c26fb7a336669", x"5798833de8e0a456", x"a91a9c88b34ed346", x"66ad9983f7877854");
            when 29659030 => data <= (x"bc3e0f1917fb6b3d", x"55fa670998b0e170", x"5482e606c2662ee8", x"542cc87e1aa1134d", x"69a816367cca89e9", x"50b291d978db60bf", x"b6bdafb96d5d98c3", x"6d5318fa0c8c617f");
            when 19223851 => data <= (x"ecebd237f6c02672", x"2fe2f015f32c4042", x"65559b45dc1cfe45", x"afd01cdcc276b659", x"6a9da86c849bd375", x"418aa2cdd8266d1c", x"a5b1adb7e834c560", x"1e63f8f130872176");
            when 11055610 => data <= (x"3fdea4d6b2aa35b0", x"0262baf24f9a2f51", x"1b879344cd8a7dd0", x"84680ed225cc3bd0", x"79c66ced4a013233", x"8790d08ca0f76c33", x"9e6a374ac1ce47ef", x"f6ab17f5281a39b7");
            when 902290 => data <= (x"7b1ce9db3451c842", x"f3c69e962fecb9bf", x"6f70ab77b4464cd7", x"3921d7752f6908fb", x"3f61a8266a54f278", x"6caaa0a2cfc96a44", x"69d6d4630ddb6daf", x"298d6221633bc964");
            when 12119121 => data <= (x"4e978e5393093c0a", x"fa32e8e91e0f421c", x"3cafc838f0d566c0", x"ac6f080f6f8f3677", x"71e1dd859f7b9b04", x"107766350a7b54bf", x"ac49aab9f3cb1db3", x"47e32adbf3252da8");
            when 11361111 => data <= (x"25c5abac306a510f", x"a151215ad5426390", x"98bfd7ef29fe0b3d", x"6b884d3719fe987a", x"79fb2c6abf5700bb", x"7d387f17ea625160", x"cd9ec49e77e32608", x"f43637fe3b4d69bb");
            when 20190576 => data <= (x"599adb00c77f2d6f", x"9002f49da27f714e", x"824f34974d66245f", x"a4991d35663cce61", x"a6ce56280ec7a485", x"7d1f5fce6372f632", x"e34698ae6bb424cd", x"9df24f317f20c917");
            when 18375600 => data <= (x"41155f346ff29ce2", x"40588b76ef5e4f25", x"986514dd8a9df487", x"1181f509820006ee", x"83f0ea60a74ae706", x"6b1e02bd852cb2ba", x"b60a13f8395b75b8", x"a3c00a4034694a65");
            when 20230410 => data <= (x"a061b58af51bf3b9", x"39261bba53277a04", x"3fe78382b9c90fe6", x"b28fc3d4eaaf7f30", x"b3932f9c87eac42a", x"0c39b4ec0f37e725", x"f05f328430fb8338", x"dbca6da007445ce7");
            when 20642480 => data <= (x"008064475dee6b73", x"e7663d5b3458be8b", x"c8c3f19c602e192b", x"16a9c6e60d6f3662", x"237d1b7fc395d16c", x"d4aab47b66d75122", x"d64a5793cb8c95d9", x"d20e87efaedef61f");
            when 22056223 => data <= (x"3def57f33a0fc741", x"77d2522e9864098a", x"84c6afd619307a08", x"0d1c09f1a24888a5", x"7ecb132d1f3cb703", x"fefee06bed4a4c17", x"b69cf13403409234", x"718a898a612f4cf5");
            when 17860368 => data <= (x"c47e6903b0e12cfd", x"7f5ae0f01bc600e7", x"a7ec9013829f622f", x"f2ea7ee58551d11d", x"6dd0aac5bd7032af", x"3afc76f00906e39d", x"ee76139b05955fa4", x"3621b9963a8fb68d");
            when 12045161 => data <= (x"92d81a1f29725806", x"409d741ba86089b2", x"0f4987435db078ea", x"08d5c429859e81bd", x"bb5e1b76429f377a", x"7cedf34f45357ab5", x"39a7491853bfccbf", x"332f85f29fe672f8");
            when 16415214 => data <= (x"efd8e35e5e39859a", x"bebb3fa90c208ef3", x"9c4c27e178c90348", x"fe8620f09f7281ca", x"53c134e22a95ca8b", x"0613ff32f31c3776", x"1dc49f1d08e0ca25", x"a3795df2b74f6e2c");
            when 19713599 => data <= (x"9c07fd04e8df0b82", x"3c60c708b51ae8ad", x"c931757f7d778f19", x"586adf8ef5ced85a", x"c30737ff57de3530", x"2b7a345d9b3f0e20", x"af832d5b0ce04faa", x"4414915a47e2d24c");
            when 10766472 => data <= (x"f90a589db5bcf646", x"22708e03c95627b3", x"792c6e50800d8ab7", x"9b3de9a0129528ad", x"ad9febb754a9c941", x"d2f9ded8e15e498b", x"c988823e23741266", x"15caf8ab4b9df215");
            when 7908143 => data <= (x"890b35a196f34f95", x"f5a150f4e6248f18", x"b02facae428394fe", x"b9372868ef8fc50d", x"0e1fa67539016ab7", x"ccd4478231302c2f", x"f3a49666a37cecfd", x"a6f77c3ec58a26a6");
            when 26941095 => data <= (x"b80b7f4be02c5ac3", x"c6a4649fa5af464c", x"b05a710afd767ae6", x"4d196b1c9ea6822c", x"8688881fcc7a41ba", x"60f94474adc35978", x"e70dac1e5ab89dc7", x"ed0bdfae8c72795e");
            when 15413376 => data <= (x"bd49c27f4b64f08a", x"a371bdcb668cad63", x"5e267c704bd53a85", x"1ca430f223d13c85", x"f8764d905625f03c", x"73a80342efe0e3e9", x"f5deb53942651614", x"e5f555989974305b");
            when 1690193 => data <= (x"00753e076db11073", x"c583b08ef1890935", x"5646d87ab442c9c4", x"e463a1299d147ed0", x"67ae1dc4875fb07e", x"30f909e1480daa3e", x"53eb77abd657b96b", x"9fbf513c44423f04");
            when 17373155 => data <= (x"6cf75c75f8c09077", x"891b88902a5734e9", x"98c7b9269d64431d", x"4afee087a3f1a663", x"6b502801d97a37a1", x"03cd8a232436351e", x"4dd0696293a254be", x"972c784507cc0340");
            when 3181167 => data <= (x"8e0a98a119e45be7", x"f581529bde6653a2", x"f68732150216d5ec", x"ddc6b96226a1ff17", x"ad8350efed7bd548", x"205cfb5970119557", x"6b3bab061c830565", x"adc7097d23192a1f");
            when 16175425 => data <= (x"b71fa9e4246b46e8", x"d232e3e491b8167b", x"bcea95aa8f0fb0a9", x"fa5045d8efe862a6", x"6283705ac8f8386e", x"64235143e19255d1", x"1f19b5a70f04028f", x"43660f07c20f4d48");
            when 18609610 => data <= (x"72881ca0d31db08c", x"5d3dd23dba3e4047", x"30e1c9f7d434622e", x"7cb7bed92e7a405f", x"89ef79698f27c47d", x"b1d3b2e991e37317", x"69b04b1716c7e7d7", x"d8fd3c2bbf9365ae");
            when 19084760 => data <= (x"10e5cc442d94d76d", x"241ee26fe194e5df", x"202e2174aab4d662", x"40631e72bd53637f", x"769d628e31b66fa3", x"c8a37ccb40582a76", x"16e624d4a51cf874", x"e3d5363e5e4aba9e");
            when 9009900 => data <= (x"61283926f0ac1dbd", x"090acc7288d782f9", x"35a6d2431523c656", x"8eb3e45180517a44", x"9cc4f95238b65d1b", x"311d3d0f816a29ea", x"ad2bedc5b289629e", x"5158e99247998483");
            when 18810409 => data <= (x"4986113b1f3c8cd2", x"c16abae54b10e7d0", x"f9ed3ecf92fca2c2", x"357031cae935014d", x"263cad966cc68683", x"13471d4aa9e08cbf", x"f6fbad08610e42ab", x"bb9f9cd088dd8bb8");
            when 20284621 => data <= (x"e7938da4304806af", x"24d6fbbc290a0412", x"7064fe710ba3ec32", x"d1ba32ef3d40121c", x"cb7f4c5ab304a29b", x"34ade0aac08b75e7", x"6386c3d81c15f4e1", x"7b9ed7fb13f2b4a5");
            when 32137026 => data <= (x"8d02bb087a019810", x"518a191606c82fa7", x"dd7d200730a553ca", x"1699f06f94a1e2bc", x"9759ad8b3f4e2abc", x"1658fa4f00bf6d31", x"468db1640fb4daa2", x"dc51eac82657a127");
            when 24696343 => data <= (x"3d563848dca43645", x"36191b24b88b0fa4", x"d36e7c9d05f2801b", x"2c7c8aa8ff7e9df7", x"e3834ad8b19e3285", x"ba2c109e00bec97b", x"f3372093f480c96d", x"01afc1644ae4b4d5");
            when 25371491 => data <= (x"8966f215a8a3dacb", x"4a8a0c46e4cc1fb0", x"7ffc37f9b2086e0f", x"bde61131dc098f95", x"8dfd31bab6664dd5", x"e3711a7be3d3c1b8", x"496a23e87aa6ea49", x"cb37d761918ba112");
            when 28059147 => data <= (x"7f8557f7cc38c6e5", x"faa6bf7b7fb65a02", x"efaac12e873096fb", x"37145f0936e0d7df", x"28a84e933d6b6b93", x"f81cfd4a89943a6f", x"e8250a9c956ff2aa", x"206a857ace962025");
            when 23096529 => data <= (x"663a62c2ab9de84d", x"a7793270973b2ce2", x"022809f517ce2dcf", x"9ffed456631b5058", x"267110bb9085676b", x"3d085443c77906b0", x"708400be6035d0e8", x"1756a1579af78839");
            when 15211200 => data <= (x"8ac5c962754dd32a", x"7551eb841d2ef6d8", x"5379d7c99a8ac5dd", x"d7e798babdbfd517", x"24d9faaf6a2dd593", x"6d7b8b5d67d30265", x"d24422c9d24f567c", x"ad497f624bef699a");
            when 1174681 => data <= (x"ad8129d35332f3d9", x"b51349f6c6accb75", x"41dc3dd30205a1bd", x"22daf98abcc59795", x"0431e152822b3a56", x"f23c4fa2cfb8b854", x"d439093d2734c007", x"db0d8c36b0016dd0");
            when 4068948 => data <= (x"a7e2b23ea342fad1", x"ced298024a0d51b6", x"582b34489f7d0ea2", x"9187749e004e1e85", x"b1d8cb255ecafb97", x"a07273d5560116cf", x"7dd14825452a0771", x"17f18201e7e096d7");
            when 30191445 => data <= (x"0f2fd3e94fcf9185", x"a23ef5efc02c228c", x"130a93256992624c", x"575ef2c45c68980a", x"9fbe491c7d3b1de9", x"8b34dcf28cdc7df2", x"7d7e759a8b723ac8", x"9ecda770b49fa22f");
            when 30078796 => data <= (x"396a59a5bb619929", x"af32bbcab832c83d", x"6c8c5c02894338bf", x"6076673c432ef645", x"7ec86a2959c1d54d", x"e17304364350b971", x"94baf0bb878c6f55", x"1f305eedc38c46fd");
            when 29450985 => data <= (x"9ed91d90a264302c", x"8c21dc289f676645", x"8f53402513cc28fc", x"1867f1f299347d06", x"4b4e5624879d4482", x"036051be1737ee5f", x"f960374529526f6f", x"4011cc8eb1ef3323");
            when 19885054 => data <= (x"5566d7148998094b", x"517bfc96ceb14c2d", x"8b709892886c0265", x"e34b5b952a676ddb", x"b0a05164bb17a5ee", x"a9cc714796371300", x"7c12eccaa75ab3cd", x"1545597333ab007a");
            when 892126 => data <= (x"caad55e06f97eba2", x"f8eafac32045397c", x"9665413394360284", x"d461a4ff7fa5fcd1", x"b5352111b651cd7d", x"5e8738c22cf4abdd", x"1431a375197ddd3e", x"b99536317d54be88");
            when 23361549 => data <= (x"183ee4f0598e1c59", x"721f6ab01920ffce", x"4662cb6ffbb32c72", x"3abc5df0693c2983", x"1bf938d062ebfa8a", x"1b7c50dd10f8f214", x"84c23b8970ab731e", x"4173e5561c636f91");
            when 30814891 => data <= (x"92174dc306a7d3a6", x"cb4a18922f80b9d3", x"97de87203c16c0d7", x"24aeb7e8f15d7e0e", x"2fb3761b2d03d745", x"5722dce6025bc22e", x"d27ce639b7717c10", x"1d88243080146055");
            when 16986478 => data <= (x"42dc36845d4293ef", x"c235c8fb8dc810fb", x"0dd7695eda217f17", x"9a4dd4310c6c735e", x"18cd0f3800b6b4fb", x"33d8addcb9530bc6", x"24e8bf2bf9b53564", x"cc56f0e931d4b66b");
            when 13453353 => data <= (x"2248732552e36f26", x"7bb154cd2e7ddecc", x"f341f75a64894bdf", x"31d50d909de17a90", x"ba2bdc29984c179b", x"eba9a258dcbec8a6", x"f13c1e6badcfa100", x"d270b8ba3e93fd08");
            when 1240274 => data <= (x"917c6173c3a3848b", x"18b97f5fa378de89", x"2abf883b5e20de9f", x"8822635db71438d4", x"7a6d5845d4709df0", x"76d1941a4faca4db", x"cad43d417a18ea37", x"be8bceb66ed29201");
            when 33358693 => data <= (x"e93d354b8c4db01e", x"823d3b0a316e166e", x"da83961d1d71d3ea", x"bf9f0c8154b0de5d", x"7ac50134b9e49393", x"45411970615d1925", x"3d2fd395a0184ab1", x"e90ceea527c0b0b7");
            when 14510882 => data <= (x"181c643acc31eaac", x"58b5c0ad3e74939b", x"ce8879f58f0e4694", x"35c086336ea16d57", x"c9cf9d37879dd2cc", x"92591deea42ee789", x"9caba9c12764f3e8", x"a7a15fa0e2907731");
            when 13513937 => data <= (x"7d3ebaa94ac49631", x"21f3278a7f1ef2e9", x"10e60ff834ae3b6d", x"c6b82bbc8196d32a", x"afc003e8cfa84c83", x"8b82db48d021bb85", x"58a5677c78531a47", x"3bab48c5058d04fa");
            when 11211739 => data <= (x"531c9d847b09c19b", x"70ec8d31a3de5484", x"6b172adb19c01919", x"332037c0ac2cde75", x"1e59fb454aaf1bde", x"1fa38cbd202656b6", x"e1a42ce171d2fddd", x"8c06b4d9dd18b895");
            when 546150 => data <= (x"3f3ad7cfd9558a63", x"345a2a6ada4484c1", x"6ace825e09d242ac", x"7518639f6ec1b18c", x"e8b22d9181dca1f3", x"9f1c81dd3d26fd3e", x"d8fc25f983a43bda", x"957155c0f484bfe1");
            when 31664087 => data <= (x"f7b662abeb377c6d", x"d2d829467822813a", x"afbb5f7183da15c0", x"64e4a9c6b84ae1d5", x"911ee554aa767d58", x"9d67293e3c737c00", x"c4649a91b34cbc29", x"a37cf6195916aa4d");
            when 15577171 => data <= (x"0f31a271dffebfd9", x"bfdb5e5d9c8db6f9", x"cc38d1210448db80", x"c75074b8716e41a1", x"73c1dacf74e5c0bc", x"ce45bf9aa03038aa", x"ea52d31d3f0fb65a", x"71d39bb83e9c5fc9");
            when 28106454 => data <= (x"57f6a7443c86809d", x"c10c9e1b70529276", x"5b47acd74de796db", x"35583723c87bef7d", x"2c1014eb7be38e6e", x"7950594cb8ab420e", x"fce583e78289a609", x"91a5237746b7095d");
            when 19666015 => data <= (x"de5d08c42cf7b80d", x"b9f6a9f00f11aabb", x"a041d89643cfeaed", x"a057ed512c6e61f7", x"b674c9d933dbad98", x"c2a317dc888e2946", x"2c99ccaf5b9d9dff", x"0ea81dd1bec20586");
            when 16175643 => data <= (x"1294507468bcaad8", x"174b9057b946268e", x"26eda63750bf4adb", x"531290cb716cfb5d", x"21980066d817fdd2", x"f8548fc082efc800", x"101dd2d73e97969e", x"8fa186d4712dcfb8");
            when 32217771 => data <= (x"4ad816b12e8b3065", x"10e875ea8e1502b4", x"ad9f56b6ac9b8a74", x"0ddb944865f08ef1", x"d5941882ea5c53c7", x"3fada02392bb559b", x"b6430f88a0efa1bb", x"bdc76ef18176d70f");
            when 3110578 => data <= (x"3bc1a742f70b07f7", x"ca29bd7c13105169", x"db0ff23c42dfab2e", x"64efb3966ef9ac80", x"5e7af90981f07e18", x"188d9b0d2818e288", x"a73235b9d2ef71d7", x"b7ce8fb797f0a730");
            when 32706986 => data <= (x"240c1a0597c6cbaa", x"701c82c49b14eea6", x"69e62c96e8bf3dce", x"91bdd35152680cdd", x"1d8c267bcdf6e746", x"38fb58de8513f489", x"1cbf15b1c33150a9", x"8c570bd134e17855");
            when 4607237 => data <= (x"3836311d5312c8a0", x"1d587c61b614ee34", x"75b76c0aa596a2bc", x"a08e5d9729c55c92", x"9d7a53e7ec9a31be", x"045c1735affebd0a", x"1a5541d2b37f4108", x"f9a692c8d87ed3a2");
            when 31004835 => data <= (x"836e3651da155b21", x"fd8fd5be41dc5ef6", x"89e5b5cf6105292d", x"05ec1272933d1289", x"4a9572f3e0ef2db1", x"4731b1a3186d3261", x"8d5df8462819b7cb", x"a2373387350619c3");
            when 25711625 => data <= (x"0a6f3b936e8526a9", x"dfeedcfd40082bd7", x"f079eb6458691a04", x"168d9bcc9a8d1a3d", x"c6bbac8a9f833fb7", x"e2af3959514fb0aa", x"04e60ccd1b00aaad", x"bc1a83ac1bba7908");
            when 11590016 => data <= (x"33986a82f6307f51", x"2291e2cab4afdcf9", x"d981eb8998618f01", x"f4a2b91a970ca6e6", x"d5afc2708e38546a", x"15c002d56c2cd8a5", x"6d0861a6eb9b5a49", x"7433ad1c4746a5da");
            when 19558665 => data <= (x"099eb1506f1b4cef", x"4efa5e2bf8de1d0a", x"b20f0a0b6563c9fe", x"21c447e95913dc1d", x"10f8ebf617b28a4c", x"1f487acb4e67363b", x"3df5ff001a3233d6", x"f3eb22bacec6a191");
            when 32965259 => data <= (x"77998c8e28baab55", x"27c35408b0fe6f94", x"cc39b1b011920add", x"bc2d7a68b655620c", x"228a023dddf64ffa", x"c15b70821e2d3bc8", x"998dd98ce81ebb86", x"f688dae1537b2bff");
            when 17252901 => data <= (x"c9fe96ae061e7bc8", x"d432ccba70aae0f7", x"382cbce36401040d", x"762f368af6bc5ba2", x"0df0e2243b314922", x"6653c767ccfce520", x"4d064d6d492d9f82", x"64e1412130037dc6");
            when 9061187 => data <= (x"82221e0bde82c109", x"b05a3dfd98f48de8", x"f19ef03e9a179678", x"673210d7a49153ba", x"d581e44c9f78c8cc", x"c563c73cd9f3fffd", x"7f8eeb93e73c7c9d", x"f394d536bcf1e647");
            when 932103 => data <= (x"0f27138e00d0d763", x"fa50da9095584ef7", x"493d46026b508070", x"2a6d9e895d7961f8", x"1197f1eace637fe8", x"a3d1c14c7e82eafb", x"40d3652e7bd8d6cc", x"39701520db352036");
            when 15257743 => data <= (x"7fa75e76f4892fc5", x"7f92c6cce5f0292b", x"fe7e6c249e7f98a1", x"6f37c1032c8f0f17", x"743ccefefe5199ff", x"d64ac75255dcfdc7", x"e100cfc0cffaff3f", x"ef1539d7430e1948");
            when 12501702 => data <= (x"f70237af9fef4109", x"7940a824779faf59", x"7382fbe42f25d717", x"7ab4e26d200c2abb", x"465972b372c9ade4", x"b3a36d9837dfdb7f", x"dfb53c7a614423de", x"68d441428fde6c52");
            when 10783872 => data <= (x"d62c9ca1dd3eb7d0", x"4345429d81ea96b5", x"38be821475cd14cb", x"9adea0ab47100211", x"2f61baccf002a14a", x"a599d7e60e5e2dfc", x"f80a3b0f978432ad", x"3213b6d44f2668e2");
            when 31551848 => data <= (x"cfa5d6821bff890c", x"f2ef864eee8378b3", x"f920adde76364146", x"76579b866181fafb", x"f971ee5599ca2fc2", x"7bda826140457837", x"33cfedb1d55d322e", x"fb61ecda6cf3968f");
            when 22132274 => data <= (x"eff07905b1149df6", x"55137ea802d7ef03", x"acbc58122d03bf51", x"c284c6856b0ef5bf", x"fd2b5482f394c3d6", x"fa14c81134d31bfc", x"9078bc2b12a89854", x"7f57a3089253d616");
            when 29938126 => data <= (x"f4216e0d8842cb5d", x"77cbe7c8c8dd8d2d", x"13b0cce2dc87391e", x"0bd974711ef9d407", x"7b3f5eb9e1ad2dda", x"1b783f4c369af4fc", x"4582b43ecff55f29", x"4d692944abc808a8");
            when 1104675 => data <= (x"3dc1013961b14feb", x"7bb7c04d2b723c60", x"ee03b88b92c7653f", x"2bc0d94ad32625bd", x"9123510b33f4c5ee", x"7a2ab3640362698e", x"b1e2ae8a53f961ea", x"890fdcf6c2699223");
            when 15528012 => data <= (x"0a48e50c296f9eb2", x"9bc50a22d6c073c0", x"65cf6f74802d9e23", x"b3ed45a636eed94b", x"975caa9a13572ddf", x"c568ae1f93971a72", x"86f7fe65e4a4cbcc", x"23c137c38e0b6c54");
            when 17202435 => data <= (x"3fccaf1e3e5a9ecc", x"54ba16ddb6d86973", x"0cc920cf5d72cafb", x"0ab18656d13758f3", x"6f8ed6a6f1666c2d", x"411654f6cefa74c2", x"0d069abaacdf5a9a", x"01506edd4b496c89");
            when 11965233 => data <= (x"8c44f839dd77f605", x"43179da08b75c05e", x"576d9d7a7d2e3056", x"54c0e97fd72c5ffd", x"25010a3862375440", x"33e923c8e7302828", x"c26afb16ebd94d29", x"87353336957fd895");
            when 33712046 => data <= (x"8e808063e94e457c", x"ab8c36d262223354", x"18a5df9184de74f7", x"ca1d502e962b06b9", x"5773bfc000cc7f69", x"802157bdfa122514", x"6617fc580cea9849", x"f74dd5210e6ef5ab");
            when 22106870 => data <= (x"d2443f98315a857d", x"25b587646a77cc95", x"cbe23d54124632ff", x"fd3b3467519a3bf9", x"892e1da7798eabaa", x"18d06dd3f881f363", x"a0f17e79144b62a2", x"41244467a9651edc");
            when 13472762 => data <= (x"f21b2c159732beb1", x"5e483032ca93aa09", x"748c76ce77e62044", x"3e64b6e030510ba6", x"d4142bcee9932f06", x"bdc42d29c77a20bc", x"efedbadd1faa379a", x"886a0c69803537cf");
            when 7434734 => data <= (x"b2e5b321686730ce", x"2eecf8b36142fb34", x"fd1465a78e366fa4", x"58ea1a4efa1aa39c", x"afc9af2b346a2312", x"e56d51b7d7117a7a", x"0cc67fdf1f20c2da", x"c2d0d3128434f43b");
            when 19012150 => data <= (x"bf1969a2d0545ed2", x"3a46913411e8aa1e", x"36acfa5a3b3ea8b3", x"baa11ecd84ad75f3", x"485617421b84710c", x"5ccf0ca5f9dd6d72", x"06f39a4bdc58b790", x"3e922dfea8d55249");
            when 24012487 => data <= (x"158c1b376a028735", x"d7d51593022d3b83", x"5e50b6ce5c790535", x"25279cecf866836f", x"2882b6c60b65aa9b", x"c34577f1012536f4", x"a81967e467a31578", x"f24afbc358e3ba41");
            when 30752654 => data <= (x"7c6f7a569902a1e9", x"65ff33fdb69f6361", x"2943667387bb4b52", x"5349905f83ac575e", x"07253669cb88cefa", x"d7adfa7984386b69", x"3a20bc78ec5948bd", x"af9ba0cdd62d0c0e");
            when 20627776 => data <= (x"8a4f27b19f3b5a14", x"bf89d9af1543098b", x"f0f2a2147ec96283", x"d16f56d71cf07df3", x"1b96768715f62374", x"3a5e07aa9d3b8333", x"44b07d6613a531da", x"ade4378064ed602a");
            when 22479726 => data <= (x"1c8171fdf326fb65", x"c510f4345653c8e2", x"fd4eb15763109964", x"e56bb230b7c322f5", x"1709f3225cf0d8ea", x"0644a72baf546ab2", x"48bb988617e1ed77", x"0e9878e187fdd6c3");
            when 9514014 => data <= (x"88993257a59a2801", x"457d210a36b69aff", x"b09d7af53af4b664", x"442ad746acf71169", x"11aedd65b8871d3e", x"dde7e7cf4c7c39a6", x"4a5276999ba410bf", x"77cacc4abab268c0");
            when 5959507 => data <= (x"fc14bb8d5c8eeaff", x"37357642d1f73f5a", x"735a07cb2cb5da02", x"25d3f622133c4e04", x"de36b71540d92815", x"f54701b87ec9e70b", x"6ce9454fa05db904", x"2c51235886d9badd");
            when 18013482 => data <= (x"55811f6b6b68b651", x"35c04bd2108fc9ad", x"e9447178d4ead54d", x"c94920013bd40af0", x"b692e198cf88678d", x"1d5c6dcd458a6996", x"c5d96fc9d9e606f7", x"73606cd84dbefa2f");
            when 21716513 => data <= (x"f9c5811720a0f309", x"522748f37081bf5d", x"7624ef04b7d8f24a", x"7d2e07a592e38ba1", x"6c440b4af6b24c99", x"d4178c55bd103c3c", x"b2f124659a15902e", x"b8d2873ca3765d73");
            when 23581747 => data <= (x"c05f09d8de09c494", x"a5d010c0fed1a6f2", x"70c10b2f2d0d9f5f", x"3cf5c26c3ccb6a1b", x"ed45d86bbd457f99", x"a45b632f700515d1", x"de286ef7548e3aa3", x"80948217489c5da9");
            when 32977308 => data <= (x"2c9ba55d0304f516", x"87bb1d9111b5b354", x"2e544c63e23cb5f9", x"a66f8f399b60377a", x"f5995ef8be7d66de", x"552ff1d8295b79d3", x"a5dff9f379748a1b", x"723a870858712f3a");
            when 26562047 => data <= (x"d02f74caa5998e2f", x"20093fb7d3efcc6d", x"a0bb6185c4c37bf6", x"54ea148f55c8e47b", x"a7d74d0860de8329", x"321d1918a1c1db7d", x"cc0a7665b46b4120", x"c5e12bcd13ffa419");
            when 15625646 => data <= (x"48995fc7388ca604", x"d1e98f7d02a4acd6", x"05b12b1fe25d9731", x"b7dd060dc4cd1f6a", x"95031e45a8909f71", x"242c5c955f0dc6b2", x"4079621e31bc5bed", x"20255ca244737859");
            when 12218492 => data <= (x"f3d6ced687b49264", x"404a77a3592579ad", x"b1efe97eb9da2d51", x"801e56e9f1ab73e9", x"439e6b0cbedd92b8", x"0c1bca66a7d11a91", x"fa0fc16fd640121a", x"f55b056860809537");
            when 23315073 => data <= (x"6f22d901269c86f6", x"4a988da1a1e5f639", x"7566eb7c72785d00", x"a236ca76629e4f24", x"8eea98834da2225d", x"8505ce6c14100ed0", x"2522a1c48e2c0de2", x"cfe9e72b9cd2730d");
            when 16033549 => data <= (x"b401798753142d70", x"05c106bde28b3fe0", x"a213a7446b720e1a", x"27d9c4c6421d9213", x"0f0b16d2b40e9c15", x"5a24cddbafe92932", x"618e76c532999bf3", x"4e99b4cb9c3dc772");
            when 22500889 => data <= (x"2cc056e92e3dbc67", x"b8f703d05a89d384", x"0835cecb26db9893", x"8b77dba9a501b41e", x"180af750541f6f5c", x"42a2971e4ce75e66", x"6158736c1ee71ed8", x"8e7730328acf6078");
            when 17091598 => data <= (x"0ceea9229fbda4d1", x"1116a3977bbcef85", x"fb67cc9e308ecae1", x"13644e01dc279fbd", x"45d6fc4c58c3b4fd", x"803d6742fbcb8d33", x"96f6b26212879db5", x"109ad01b1788bc36");
            when 6340592 => data <= (x"e09a288d10f2d092", x"c9b7f26f61f651ff", x"9aa2d2a6900c41a0", x"6296083a6c86019e", x"4bbb3d34118d7a0a", x"b02b44b130b5787d", x"37938b47fa3ccf3a", x"a5160596a181b33a");
            when 32254807 => data <= (x"e06ef7332b4b1087", x"0ee521ff197a312a", x"54a5dfa45125fc55", x"b57fe628a3edd690", x"d18db2e3eb3ef568", x"e8ca548eb51f477b", x"0daedfe0d32f8ede", x"267562e55c4ccfc8");
            when 24356155 => data <= (x"059f5475d7ce23b2", x"80454dacd3076871", x"c17e590f7be4e023", x"fd75fd585ac99545", x"86e21d233f91b529", x"697c33fee2aaf75e", x"106f9ad93bdb69aa", x"9f8899904a4144b2");
            when 19503989 => data <= (x"5e0bdd80e247efba", x"74b8eb2c524042b4", x"a3efa3ebbc7494fa", x"779d86760f332d53", x"adde7501eb2895fa", x"a5e6701d82c8e607", x"c70aa79f17883c7b", x"8ec91cce7cf7dc27");
            when 837024 => data <= (x"366645ba89d119d5", x"1cf872d5723c1d1d", x"fb8d83955f03a137", x"48a223ab3b62dbb2", x"b720604d9cddd080", x"b90074fbd4b3d03d", x"f67876139ee62ba7", x"56a558b7b776f83a");
            when 19898698 => data <= (x"5dee4af6deb88ea6", x"880dea30b746b5f2", x"b1002826a6930e8d", x"b949a5291e04c0a0", x"82fbd18deeac11e9", x"e2618887f2f247f4", x"4a9bfab254cd1419", x"d051a49987ff6fb1");
            when 28498827 => data <= (x"abcec51f287f44a2", x"63c08db3577b1482", x"371be1a4a2e8d6cc", x"ebb4dd4c57ca7118", x"e48eca3609fede73", x"3b486afd9f51347e", x"ef2d7e82e2495dc7", x"7bb0b8ef7c0ecdba");
            when 27757877 => data <= (x"742e634a7bdf3449", x"56eabeb294d7d255", x"1d60429aff793dc8", x"afcbd24209003b6d", x"f3deb2015f8bc6c3", x"5f2fbcf70daa93e8", x"3c39d8421adc64a6", x"3585b0a491664970");
            when 31989217 => data <= (x"fbe5a0aaa3d01d3b", x"963e2ba1dbcb1055", x"674fadc044a0d11a", x"499257877cefc73f", x"dd9c52ba0615869d", x"f9361588c7857070", x"decd22888a4bf32a", x"61452162d6125c7b");
            when 25107053 => data <= (x"14ffbda7309b029f", x"d4ed335bafcf20b1", x"09321b1a33f5367d", x"8ba28cdb7db0afcd", x"b730b00d3e3980ec", x"7445c4544eeb8b7b", x"5304dd7470eab9da", x"e1811503565ec57b");
            when 17499986 => data <= (x"1b1dd6e17d3058a1", x"1afbf2a2488a8c1d", x"7c483d22edd1f1e0", x"607a0b3aa6a19e2e", x"8c15a0823ef6f233", x"c8c7fa39de9779fb", x"7cfa0a246377f83d", x"90e3d4837911e197");
            when 32933187 => data <= (x"2be89bb68705ab21", x"143a1339ad603621", x"130319b8aa043cb7", x"0f3984a39457c985", x"b5e8b1c51090d7f9", x"64d6f3e3e209c844", x"ec7d6600af5fa1f7", x"63e8441b802eca94");
            when 24318385 => data <= (x"c1deda0fa55f3c92", x"5e1c172288be0c05", x"a5b085cf35bdb059", x"d238bdffb50e6d8f", x"05c15ec98a299787", x"6a5f07c247d023ae", x"cdd39f3fc82d4ddd", x"d1b51b93475b9549");
            when 33740746 => data <= (x"52a0267c26486d8d", x"6dcd12e2c6c71ad4", x"bb7eb3f56b7229f1", x"83b4115502c3908b", x"696fd80f25cae026", x"e19bd07d64561278", x"18d215c9bd960c59", x"c12920490f88bc1d");
            when 7964412 => data <= (x"c36bd159394be523", x"d4b6f14b3854c88d", x"f9c4a6b054e3a70a", x"d9a65e62916803cd", x"93f350178c012235", x"f8e61e44829b0f97", x"14fa20664b3a303b", x"2d2aa389d9c8ea55");
            when 10901483 => data <= (x"fcfdeacc7cb14feb", x"712ae0770c79f70d", x"8e79d7fdf8911da2", x"7aafa910488214d3", x"4c3ca6976eaa32c8", x"4823136f8d4d25e4", x"5932eda11c169c5d", x"33f8ccee4a4f0d1d");
            when 10138709 => data <= (x"3fda2da7e7c1b02f", x"c85e4730eb444cac", x"0fde9c4f221c2cdc", x"886d9485eddab096", x"78d65fb2f990fc18", x"d580084e6f85feeb", x"912041de3c5fb95d", x"7c591363d1d636df");
            when 18055325 => data <= (x"a1b5f8c25e7cfa37", x"e917f4afcc33584c", x"96ca2eb65bccda62", x"c87128f78de952ed", x"f9911a100fa971ed", x"4bace63c6af7dd23", x"afd88c4b8610dd6a", x"ebd9593ddfb97596");
            when 15754873 => data <= (x"96ca83b7c6dfef77", x"11cfd3a23927deb1", x"758a63446ddd308a", x"35dc1b22c0a6566e", x"b1a43dad84f7ef0d", x"6cc863d4df5dca7e", x"3a44776cb97a7472", x"3657a9408384065c");
            when 18366722 => data <= (x"af34bc8959142c4c", x"98205750f8203b77", x"f955e51dda06c061", x"ceb08b50134bf31c", x"01cafbf0289c3886", x"15a293157348b875", x"139372cbba0c2466", x"2a6e4a96a7d6697a");
            when 17215709 => data <= (x"eb90339910924665", x"3d8593496bcc0d0c", x"0a17e120aebcea0f", x"0c4005c528be29bf", x"86cb8f7d5b631192", x"740f1c9f95b02188", x"e409a21d5ccd86c9", x"be5b4984735ca8ca");
            when 23156324 => data <= (x"aff2df141e6edf8e", x"1472a63f114cc6e6", x"92cb7570cf9c057a", x"b20ddaa4f13dcfa4", x"783a78e79fad5c3e", x"b9661b1693ccf04a", x"b3e0a3d0197342f5", x"2dc6cd59ea5430ad");
            when 32511118 => data <= (x"55441ec3a9e1fb5c", x"2a47ed629fa3897c", x"6840d381e69bf5ac", x"a63e651064dc831a", x"ca646a5b290244e5", x"397ce4d28c4024a2", x"07c3199fb0bdc2fd", x"6f3b44b07b96102b");
            when 28313870 => data <= (x"8ee67c7f4a40658a", x"e155fe7cfd6d5c02", x"0f40210379c33da7", x"b7b11dd5ae5de3ea", x"ce02bee8500a2320", x"0ea2e8d7d2f170c6", x"63a2cbded0d5ead0", x"7c41caa2aef7ac43");
            when 3251163 => data <= (x"72a8b66f68a03ffe", x"8b841eb3b770da71", x"32c92536d8947dfa", x"5bb191832f28a079", x"fc2de2ebb699c965", x"98f283de7a799c9b", x"7026d7faf374afb0", x"f4ee2ebeb93714e2");
            when 29243210 => data <= (x"a578bda7b1a667af", x"706f62faf209e280", x"6d03669e17599ca9", x"deb1037db16e27d9", x"ba21780171c0f6f0", x"402e996e7c2304e6", x"228696fc25495c2c", x"dee757d33c47ffd0");
            when 2978403 => data <= (x"f65081a88c4d2b6d", x"7a897b55a35b4745", x"012d38aaf85ded7d", x"46b295622ba48b21", x"8d0fa6595c3e8d7e", x"ba7c1cd075a25243", x"56cfa02aca3b11c6", x"5f68e31313326a3d");
            when 1239844 => data <= (x"0c0cb3548d127322", x"d046619a0a381437", x"4eab8f618918d027", x"424526fc59bf5268", x"033b1176b05672f2", x"526d7cf610b05940", x"345e0c2a3f4e6ef7", x"25b0436db8c3899f");
            when 5927793 => data <= (x"ee006e0af690d566", x"3c545fa89ad0c478", x"d57ff241b7d22077", x"04c45fa8ba09f273", x"00ea068532023f63", x"3bd8600196fb423f", x"cb405e13cc379065", x"8f816d82d7713972");
            when 12855353 => data <= (x"2916ccccae69ab33", x"2c54b7a453ed1055", x"435704fcb47c2018", x"874b901215debb8d", x"a38b7dd7055961b7", x"e1c979ac9dcdf12c", x"6681bba134390872", x"9940dcfe9bf35ceb");
            when 8039413 => data <= (x"cc296ae1f9df5af0", x"93d95f57e10510d0", x"8ac1ca47629e7c07", x"c7a85c2cd665f12a", x"016c48d7c950edea", x"c6682124b2eed141", x"26b67a681fd25e2f", x"5f0048f5ceca24b6");
            when 31768718 => data <= (x"d4378db923769bca", x"fab83337d9e3ccfb", x"e960f392d929ebfd", x"06579301d531b34d", x"1b474dba1a8530d4", x"268fa339227b4038", x"8837ca58b63b481a", x"7009867d33b13a0b");
            when 28784136 => data <= (x"e5e1ad6b7281ab4f", x"d6635cfb5468005f", x"75d5934d161e35ae", x"153977c71bff9794", x"718994569decea1e", x"bbd87b1148c3b770", x"91ffcadf9f17c715", x"6ffdecdc8e6a62b9");
            when 30228127 => data <= (x"38e4fe02eb4d5ab5", x"d70a78420d7198df", x"2e9c2598d775d2ce", x"49dded3f07b6195c", x"29b494b78478d42e", x"e5763c87174c2eab", x"8f54e4ee07c22953", x"03928106ab12f7db");
            when 7305516 => data <= (x"70a93053b92371d7", x"f176f3a31df94fc2", x"9b31bf79cf469c67", x"7b0fb146b28c30a0", x"17abcfbb835ed1d5", x"412d17fb7f3b97f8", x"f8c6409b556636ab", x"26ee26da272d954c");
            when 30384953 => data <= (x"31dcf5e511c84ecf", x"5a6d31861b6fe563", x"60df388e3e01bb71", x"42e487ebed33ca58", x"0c9ad2188121d02e", x"855f3cc6d1332602", x"d5c64084b1da6a7d", x"2ced131476a35ff9");
            when 19206899 => data <= (x"4bff73e5e24cc6de", x"6f4a0f563289bb4d", x"72c63a907b06042d", x"2c8ac22457cca131", x"05847d627dbdc9d0", x"6c47f24585307975", x"0decc33b418df812", x"e784be21328b9890");
            when 29392171 => data <= (x"1bd9796d8bad0d62", x"31f57088dc40f9a4", x"218fe00613ca9a5c", x"c44a9b4b0e0127ee", x"91002638abd42842", x"10827371a77dd7cd", x"9199306ca6ba3010", x"c84eeea54a660a38");
            when 4485901 => data <= (x"d5b6edba219e4b8d", x"1ac19b586f379b07", x"8e7b89a73f0840c0", x"0a0b8bc73366f0d2", x"feed29af2abab019", x"9c253bda815118e8", x"e51080ffbbf33ed0", x"d165fc0044f3f846");
            when 4498159 => data <= (x"641174810ea790e9", x"41d0a46ab615a5b6", x"ec6aea530ec906da", x"2f48050779b8ec81", x"e53afe543226710c", x"5477b4a824cf78f6", x"8e9730429454813f", x"11f5f6ab07c92069");
            when 10369464 => data <= (x"63793f0fbda03ff5", x"e5a25ee6c8273aec", x"bd50a76724e78e25", x"596133b5bf8e047c", x"2a1922e6dc96da27", x"59f6483ca5f60a6e", x"1d9f7a74aa14af3f", x"8e9283b05542883a");
            when 26886830 => data <= (x"8773ad015c8e4920", x"7faa412ae88abf15", x"f2933978c9cc2747", x"f4d5dadfed1c575d", x"b482288721200ff5", x"9a323828365aa3f1", x"5502b051f8f7eb20", x"ebd9a74abd2e68a4");
            when 9668226 => data <= (x"65009735e8ed239e", x"3d7ed2d9c12ca8d4", x"58e852403409c125", x"04f1458e5f131a5b", x"74f73856748159d1", x"8116bbcf83142bee", x"904df1aae461677f", x"df7770201ba3c536");
            when 6507579 => data <= (x"d4db30952787e715", x"050867b5bada4cc1", x"d4586dcd07000ba3", x"e7f41d0a3c02dfc4", x"96021341844bdbe6", x"200c44e003bcbbb4", x"0d980d8a561ccf33", x"358635fcc3d313ce");
            when 15334767 => data <= (x"e51887625e8106e4", x"58896b44379636b4", x"b2bf6ad31c1e1592", x"b617d8d75d812883", x"1a5bf69c7eca84fa", x"9afa33e1ac60c98f", x"3b737f8465fbdd7a", x"6eb094a737d6619f");
            when 30588051 => data <= (x"200ad7c78bab21e3", x"b696146d28c7c3a9", x"ba6e65b57dd30f9d", x"a8b527761836c7ee", x"cce5a1505361e0fb", x"2c284b07153cce1b", x"cf9dc2fb55dc8250", x"c4cd0baf30b8925c");
            when 9424258 => data <= (x"85e798bd9e11b630", x"12c377c5cebf604b", x"88f938869e8d6809", x"9f8c26a79b5c1813", x"2d0f3fcfaf92490c", x"f66fe1a48e3b8035", x"03210d264e7ef62e", x"e69c7f3f469eaaa9");
            when 10326449 => data <= (x"a495bca345761c98", x"4a98f33cb142870a", x"bb5afd9398f6d326", x"a03673ae64c19138", x"0823e777a936507b", x"a15b85413c42cc38", x"f17e193c98a0ae11", x"e5d8e1c77ad49070");
            when 6572185 => data <= (x"2cc0b39a5f86e0eb", x"32b1d89f4711eeeb", x"7dd8ad09d42e1017", x"6d8c431e7e5295d5", x"a5de33ed457821c7", x"34c7b5e7205544cd", x"c6941986af4d9d3b", x"8564490e2c9fa403");
            when 16402000 => data <= (x"287cefff464450fb", x"e9700eff9383efe6", x"eeb3cf0f424d6387", x"41c1c83076a94986", x"524dd977f8eb4fc4", x"77e040e36e002f18", x"685bac8b43177764", x"d6bacb8b4beb1284");
            when 30253977 => data <= (x"53718abc7e3329dd", x"2d993b0f11112233", x"c288bd3809e7dac5", x"1b1d8f53a5fdc005", x"cb5da06b8230896b", x"23dcd378eca4324f", x"17f50347a2728806", x"590c7a053b0acc79");
            when 12222523 => data <= (x"fee82731e98dcaab", x"fce1b8d20714f38e", x"0cdb6b77849d6cfa", x"0802662ed8f9cacc", x"4981c10a97798bcc", x"ad2cde93da0774e9", x"6c27663947fd5bbe", x"6bb9277d6afd858b");
            when 17938332 => data <= (x"80df92a504dadc9f", x"5d55f01f21b104c6", x"435ac9e115a1fed0", x"1b096b736a3c5460", x"e8ec88b163a95834", x"e01941acb63a6f8f", x"72152426f4b616f1", x"f1ee999d86ea606b");
            when 13726963 => data <= (x"efb1b5dcdab639da", x"a0927c1681b21359", x"25761d816cf05c3a", x"8f4e2a81a74f697f", x"05feded68ce357d3", x"5765ad4794b1c39e", x"3f1f8b8195316987", x"b57a4e3a433e3cab");
            when 10137899 => data <= (x"375fa2bd1a89f17d", x"ab1a3e8cd14fc7ff", x"6093f62b1962f59b", x"466c8bde23c1401d", x"71706bd20ee09258", x"b5101af9b33b1373", x"d202b690cd3a761f", x"a137feb184519f22");
            when 19757255 => data <= (x"877d4a7a328b64ab", x"785c429220feb3e3", x"0e0dc6161c6b665d", x"9031db7b497c1528", x"af7988d4e1bc0494", x"ad89091999356efe", x"5ef19d532ad69979", x"dbf5e2132a3e3f47");
            when 1311363 => data <= (x"f2bd17bd477ec2bd", x"539ada532217678c", x"657b95a5f8d51233", x"feb535b5f3d0bb3c", x"df382541e9fdd4b3", x"15dd036b39000683", x"dd0f5f9cc23013e6", x"8eaca2f89b08e149");
            when 17346105 => data <= (x"0aae47bc7cc2bfd6", x"2b52e61599358783", x"cb76616b51f3dc9a", x"684a1e3b39f481d5", x"a3d99f2647cea3dd", x"10ea1cd3d26d7ff6", x"3480973bd86ccd1a", x"276aefadb259728d");
            when 23384700 => data <= (x"2c7334ee7e78df1d", x"bf052e4f1660b762", x"faba95432728588d", x"6b0509bb12e6255d", x"7853817cbe6fc2a4", x"935d401edcc2ba08", x"5b1591d269e75daa", x"058ed16b0e1230de");
            when 33915040 => data <= (x"73258015ab73b30a", x"aa62cf4c3319a459", x"d3f5e7a4fde648b8", x"7cd26a7c1779395e", x"7e7409e8b3773113", x"b0a890ffbe549d7a", x"42b433d5a5469666", x"224639250d83517d");
            when 14065916 => data <= (x"74d5d574ad283a27", x"587a0a25dda83a41", x"525f3af80d8337f9", x"d74aa709afff4128", x"30fed0e99a17abcf", x"bc10a4c195186cf0", x"e224020324ba3dc7", x"cc766cc0cdf6bf31");
            when 30775775 => data <= (x"016ee3d897417eaf", x"44802434b8faba47", x"e04daa4c1226d5bf", x"206c3e38027e0073", x"4f580852c156a398", x"13c10f43ebcc8dbd", x"a3de96d9cccbf710", x"26e03fcd9d5e965c");
            when 7476347 => data <= (x"51b3fdda19882158", x"14a825cdac17b043", x"f5c754021b58c761", x"d38f13342738abaf", x"9bd576eeb5581f65", x"7ff10ea5449f87ec", x"e2b58a1f2bba2ab0", x"0905d30be9cbc170");
            when 22321286 => data <= (x"eeabb5a6652aaffc", x"8aacb6286c315640", x"85053cca6528378a", x"3c615969949a4865", x"53ec97ca6e8b5a25", x"bcccb19557e0dcc5", x"d85a30e0c52e9126", x"49cab92ea4612109");
            when 23494480 => data <= (x"b5e29ff9016fe4ce", x"75de16807d1c1b36", x"b08135ee62b243d2", x"a2e016f3ad8dc21e", x"bb249a70db37d8d2", x"e31529c662829fde", x"0371485090e4b590", x"8093cbf444f23747");
            when 1062415 => data <= (x"2a6e622b3ef84fa2", x"b178b3f8007994b5", x"12a03f826cd320e0", x"2b217150a6bffb6f", x"b042e5ece161c575", x"41ff1a7e933de63d", x"bb7e0b8f48b2ab00", x"7f17c805ce4ad1fb");
            when 10236817 => data <= (x"7d88077b2f5f58ae", x"b1cec5d7a9083148", x"be6a54c63f6d2ab6", x"5279db8805b05009", x"4b6af62d160f465c", x"ef13205ad1dbf649", x"fd6e352c048d4a25", x"898961361dd78a60");
            when 18071783 => data <= (x"8c352c589b773e8b", x"85844b0b25e49334", x"188f28592b05a1e6", x"930e61e3fe7e86ec", x"20e2b487300c0ca5", x"13085bd2fcaba11a", x"7711deca83a6eab6", x"095d4467c8dc9f71");
            when 2823686 => data <= (x"bbc80af2a8961dad", x"efdbdace8a09289b", x"26c658aef18ce5fc", x"2f06ca3d6d13862b", x"7a51e5842bc31b66", x"e9a6763734792cba", x"84589899f26d50e9", x"111683eb94d508a1");
            when 9618388 => data <= (x"e0e8a4f842270306", x"500019b88cb0edff", x"05dc91a6a84ccf7e", x"b18d772f1b74eb18", x"ecdb9bff20807ac7", x"9bf6fe609e3ca852", x"e68376ab17a245bd", x"f410157ab7a367df");
            when 21069570 => data <= (x"15c8f84a736f235a", x"b782f8e98e30e8c2", x"e9f4f25643a82c0b", x"3e67024c12fb5282", x"d88d67a4645f83ff", x"98dd995343ca5e88", x"581a29b3b4b54615", x"b431c1500c50006f");
            when 24771086 => data <= (x"eb5977e04d426abe", x"9ac10839b1233db3", x"cac8bf96747b5890", x"eeaf93c2d8b52d6b", x"403181c4444314bb", x"fb015be91e55e9ba", x"51a4158c923fb4f3", x"0ce24d0acaa7a8b2");
            when 1309268 => data <= (x"8e1497c7b35103f2", x"fa441ee36dbcce13", x"c440c42f4f207760", x"a7e2a471e9d13f2c", x"8495ee51bbf84651", x"a66cabf7d96691ca", x"30d244acd897092d", x"6382bf6d5b768d1d");
            when 8349137 => data <= (x"b289814db0fae7f1", x"f658b5070e8f576d", x"b659794c91a9193c", x"9106d798e847a55d", x"f73a05ce254388d5", x"1de5b9a77300953d", x"818c3cb998eb10f1", x"a18d65b56a0e1b39");
            when 14897840 => data <= (x"9748decfd78a6f3f", x"b00136cd225e1c28", x"31fd883b7175a676", x"bf379d7e2056a0c6", x"91fe70e70326861a", x"5b82691050fce5a3", x"7eaa6126ad0345c2", x"ea7a3c02c36600a0");
            when 22985022 => data <= (x"8b739ce50ff53208", x"8b5e512f9c7842ba", x"181b8e915a9f3b8e", x"7231e9cbd83f93be", x"e395472cf000e6cf", x"191c8f02c0f43263", x"57479d29446692cf", x"99754baf78ea0daa");
            when 8771251 => data <= (x"47d2a3f67dc09a0e", x"65b1db30c5e63e93", x"6984edd535a8c42f", x"6e18fefb6308d25c", x"9201d029e4629d8d", x"5da5c884642772c2", x"a105b58273690f51", x"c2d2dd573c89b6be");
            when 21440038 => data <= (x"224aad14e5f217e3", x"a08ac3a99f319cf1", x"b03d2b618c2ab0e8", x"56f75a611f3a2bd0", x"f624ba87bd5ce3a8", x"3a834e5f3cdebb1b", x"47d3971d541aca90", x"75354ceba2e88107");
            when 4040421 => data <= (x"ba964300678017e5", x"b988b449656811f6", x"8ec500cded617c85", x"18eb3a68bf411535", x"060fbddf3a62e375", x"85a269dd075b0b15", x"2ceb1015eac303f0", x"e877570ce8f9c252");
            when 9157633 => data <= (x"7d326849513bc078", x"abbaae00c9228c7c", x"04d609a43fa70561", x"0bab0c7b8877ac7e", x"7538b6fa6499644c", x"5338a04f29ecf48a", x"f9479f42d9ce159c", x"0a6690572154a4b5");
            when 3552762 => data <= (x"52dc3cd4db4fc574", x"b0817dc70152a02c", x"c640f1bbdc53e46e", x"33bdd12816b67045", x"59b813a99148efec", x"069aa116b1ab5d1b", x"c77d92698fd49d48", x"a41057bc56e47e06");
            when 17296325 => data <= (x"85bba3cf5a070f20", x"15a9c2eb1513a226", x"14203b68dbc16cc1", x"e240ce6a66d0ed1c", x"dfc035efa5994165", x"c2d90ca982433abd", x"4b1af989059d9683", x"5ad6c5eed90081f5");
            when 20429289 => data <= (x"e079072272596247", x"37fb356641bbde3e", x"6dd5b7f6ff34f637", x"3ccf5a49a156e0fa", x"0e1c3d81d3794e8b", x"e68aa104afd851e5", x"68780e8b2ae4ed5d", x"c49e7ac531e9a777");
            when 20510680 => data <= (x"6de4230d092fac01", x"0b851dda092cab5a", x"e02034d0ef991611", x"f14bca8093059a8a", x"29e189a7340335a2", x"9360fdd8440214ca", x"d143f6c291d6d0c0", x"3cbe412e828d07b5");
            when 11959379 => data <= (x"8eebc7607cc32019", x"c09f3624345995f8", x"6ca4ae90bd725435", x"3cb80d689be57818", x"7d7ba1c61fa0ec2b", x"f28335e5f7e63e21", x"b091e3ec81ee462b", x"6c825db2e457a65d");
            when 3153714 => data <= (x"360e4c0de18ab018", x"c99debc4d48b5cac", x"287d68b38dec72a3", x"18332a47fe2869fe", x"b3252e19416411b0", x"cf7b5d548db79a8d", x"bb89c82b72b17e57", x"7aec231e88bc1d44");
            when 31440128 => data <= (x"e7b133a33f3ddbb0", x"fdd1c78d37619d3c", x"a4ad42c826fb1cf6", x"b422e4f9261d65b2", x"db2b6d143e41c5b4", x"b113f32c61ebc777", x"529733c5c2c4c2e7", x"a9db402896d41c17");
            when 24090942 => data <= (x"ef845d236a1aaab8", x"4e0563ba877d6151", x"12f0ff01c0503d3a", x"9cfac4fd95288268", x"d5c3a4bef61b3194", x"bdbcb80b5261487f", x"05a6545dff18b016", x"ed8979fa10196733");
            when 5865361 => data <= (x"ec619b3a986a6522", x"46b39256f05e351a", x"414d5b9a0f984c7e", x"07a853454d5b2d03", x"327ac93952c5b969", x"6d594ae378177a2c", x"7d81d75bb593ef79", x"2b2cad2e427e1a83");
            when 17736241 => data <= (x"1c184748a637ac9a", x"0d1841180ca33538", x"1f3864240ffb7bdb", x"9bbc4c12c224a3b1", x"90e2b73a9174e572", x"9a3a6f3e13d7ef0b", x"cb843025dd06056d", x"a94e9f95e2662652");
            when 27267364 => data <= (x"ec5ef0ab8f2783c9", x"61ac6244eaf22edf", x"4abb3e14b10243a9", x"f9aeb93519ebfe16", x"5b3100ac3258bad2", x"4f4885dc78482a83", x"488d047c6d3bf71b", x"5dd9bd7ec65c095a");
            when 1595868 => data <= (x"0aa883b250e184d2", x"bcbdc6daaa4c0ea0", x"89ff41eab02f16db", x"8fbf8e52c8282c47", x"d33dd468bb053edf", x"b9b06e319809addd", x"b0dfe56866ccaf10", x"9677b9c8289508ea");
            when 15164769 => data <= (x"2b6446759416b01c", x"d4518d9e9ac26e96", x"0617b594440fe39d", x"95d45d0d90f44d80", x"7b6b608ff95a054a", x"c9d8ae49a6240938", x"b51a6c3bf1f80ac5", x"cfd04c40b42c9d5d");
            when 13116000 => data <= (x"22a61fb352a3612f", x"1590af4d4bdfc0c3", x"95c6c9eea3fc3572", x"e70af752fb848bb2", x"85beb8227bf575d6", x"ddd54ea319df4404", x"2d2024204b461aae", x"90e2570a0b9171ad");
            when 32650830 => data <= (x"05e1a3a328f0949e", x"9feebe14b7aa1f38", x"f2a786f770802e16", x"c8c7f325e3532e09", x"56858fac9196faf7", x"379dd44419b4cdb3", x"f9044537aea1b956", x"7415419f3655fad5");
            when 22048101 => data <= (x"7788fef7b72023d5", x"95db2031d51bcf8d", x"00f7c870113b8ee5", x"0d3ef693b12c7341", x"08b46185aa6691f6", x"b7fcbf3ba535375e", x"0cf8c4ae8309a84f", x"e85f0addcd981d47");
            when 30227820 => data <= (x"072d77daaefe3f7c", x"bd76175ced5ca02b", x"84afb2910f9c55cc", x"889e7653a7c90c47", x"efeb0304d3f8a833", x"0f8764f64801038f", x"5550fa6a11caba11", x"1195646bfdc5c58d");
            when 18363494 => data <= (x"5690c44b039359d4", x"87039b617f39b66a", x"5e1d7f26e93dba83", x"54e18881f2f6e654", x"3f9e9ece67a5008d", x"d4d80a610204e594", x"7850007582715d2d", x"a6fcdebfee374c71");
            when 18550594 => data <= (x"82f84409d8f87c50", x"6a1a86821deb6cdb", x"9af7af75c5f40650", x"0b4fe5fbd10b108a", x"7983c310d23baf56", x"7f4ba11919ce235d", x"4cb75f9ae31258d7", x"3003c69c973812a7");
            when 23714512 => data <= (x"700c21860476fb56", x"894db9d84ecd9ec7", x"7635400925fe3610", x"86c28b54b2e31f04", x"2f2a855a8734294a", x"67e826eebc0901db", x"205208c3be312a45", x"d8142297c7bdf6e9");
            when 30967082 => data <= (x"ec0d56bf688df361", x"fb9fb36247ea7bea", x"00fb312e1a99530f", x"6d48c2a37ec0ebc7", x"31468e290a32bc80", x"bd5cea83909d070b", x"8c5abdd469530414", x"bc299a7e6e8b9755");
            when 8528236 => data <= (x"f1b4b9ee1bf482d1", x"e541a1863b3361a7", x"aa7b135ddf9d21b0", x"32491cb9a245bda6", x"58f3d093cc785f57", x"28f869bf166a3fa3", x"7bcc5e7ae5545b2f", x"ab90b99c629659bf");
            when 5000304 => data <= (x"1f7aeee6caa8b290", x"51f867ead5162969", x"4d2c027bfe6cdaee", x"34b337bf153c98b5", x"1ffecb02a4327c06", x"4b2262cd0e3634b0", x"02616463e1a1fd5d", x"3fa294c8c39524d0");
            when 16575567 => data <= (x"69a14e8ef9efab1e", x"10983f9cfc0060e6", x"a8d84d21e7bc943a", x"0e9cbca9ff093b30", x"b06377af94e8eb20", x"f1c449bedd3ce228", x"7639202adba82c0b", x"ea563b72aa0512be");
            when 28804509 => data <= (x"e0f2d3c27f8e9b9c", x"c2830d3e79b586de", x"a3cf7d5ceb94b83b", x"35a53f28ea84ed89", x"f966e6d0bde9bc84", x"834bb21bbf812799", x"9816e62585e4a496", x"629d1353551a1d5c");
            when 11794344 => data <= (x"c707a83aa11686fc", x"5ac7478da72beb03", x"0d533e7af31e5e6f", x"6a570ece22229f32", x"3557e9ccdf0e327a", x"c3638c6100d4bf39", x"fc8dace1ecf0fb53", x"cc96b4df4dbe2ec5");
            when 30941261 => data <= (x"9c3c0b2451326a38", x"9e7f9c025c51e7d8", x"7eb540ef82e4e1eb", x"2dc0c569ca12f9e0", x"152e84c8b48de08f", x"34bc9c033c235d8c", x"d88a0c245cdaa725", x"58b67b60e429c68e");
            when 25283773 => data <= (x"0ed8c2b2997a00de", x"13b3bddccf6b7103", x"314e17b6d8725ab7", x"60a33abe3e008459", x"e2dcded2b5468cbb", x"c85bf2c27438411e", x"3918027a45e90898", x"4cd3deabafd2b00d");
            when 3152113 => data <= (x"fde6680c24323445", x"6dd98ba1fee4e909", x"4a4c81dc7d3c613b", x"545bc594bd556da4", x"4cf70e4910374618", x"659e7b9c28e02f68", x"af230165fea1feb9", x"9544bfe8a4fbf010");
            when 25346238 => data <= (x"629a096aa0c467d5", x"b8ad0f497268eb65", x"e74148e3e235d5bd", x"d3d484c4b5a96eac", x"c9d6531f2990bbb0", x"49d5dbd01c8f9596", x"d597445155e6df5f", x"dd7d452a9ecd4315");
            when 8657188 => data <= (x"ebae492cf91d7236", x"54f64c72408def4f", x"6046c1a7cbd3f48d", x"e18b193f6ff66f5f", x"793594e95f7b7c4c", x"10722dc92f5f8161", x"307ff3f7ac6473a7", x"9e7c53415cbaff44");
            when 9397108 => data <= (x"783495df51256be0", x"78edbef5b4e3c4f8", x"4c50e2d4c724187d", x"0b67207592a16257", x"377ce580cd0b7c06", x"361d56eec7ed767e", x"1d756835669d5c70", x"afc9741410bbb12e");
            when 13950954 => data <= (x"18ddce9c7a1d223d", x"3895bdb013c28cd2", x"ee4537bc72203d6d", x"61f25127ad17c49f", x"e6568f9d14553ea1", x"62ca1f178920c1ff", x"ba851118b1c2880f", x"250cf325a2d2a5b6");
            when 5383966 => data <= (x"c17fa38a1f4443d0", x"25e0a15720a0630f", x"70f7dc3139e73acd", x"cc515fe10764c46a", x"c24d5162e0ca3f8f", x"bedfdb07008a967f", x"4a99d363a472ac5e", x"002052a4f088a8a5");
            when 33180165 => data <= (x"4052e3ee7023275a", x"e4442810cfbe999b", x"b3c43dd585002205", x"f6b376b418c57e36", x"51cbde9ac81ff73e", x"f5403f1f392870cc", x"cf5db41fc45f66c4", x"61a9a8a1dd7007a6");
            when 31495589 => data <= (x"87d5eca6b5405445", x"df54c99db9e50b4c", x"44ad3b9a6a177cdf", x"9047de3abdd30efa", x"ce0dc5ecc452f83f", x"73c6135b0bc7c732", x"7dd7e547b041ae95", x"07946c9363c2c91d");
            when 16999605 => data <= (x"310757bd60ffdb54", x"09f60b4eca942040", x"85f8628203902f67", x"ad21af355bb3a663", x"07be9eb1949be077", x"d743daceaa930f62", x"a7e03af1798874fe", x"00e07fd73ea27634");
            when 33492990 => data <= (x"503bfd6bf6e3fd2d", x"d70a0f81a4c27a66", x"38569471379dfdbd", x"139f265983096fcf", x"0a388aa20b702609", x"3e6e4044cb6f6099", x"95d547281180fdd9", x"c74ed53d727645aa");
            when 20152233 => data <= (x"a89c706b88ac332f", x"6f53cf039e6634cc", x"2e18f4ec924a9d8f", x"3c8cabf70c49de1f", x"00aabe47a5b6a13c", x"cb0c70ee9f9675ac", x"e3a2157169d41b02", x"2eb5d414b480150f");
            when 31264824 => data <= (x"1abf998d5488315a", x"d572b3eaa0db8936", x"f45f04aa0fc8473e", x"36f729999ed66bdf", x"1283c85c2d94bbdd", x"493e83117e780fe8", x"98ee130952fe67b5", x"19a8e3d865a38197");
            when 1930151 => data <= (x"aef1f6fd8ff691fe", x"b4d8e06b550ffb07", x"dafed4ecc0fcb643", x"fa2b1ea95707500a", x"08e29d38e006e51e", x"b72428c7d412d6ee", x"0ab152f94941df50", x"4ad550890532d92c");
            when 30181763 => data <= (x"c9defd1da9aa3b0a", x"4ffeee0b344b7ef6", x"474b52c7fa5c9b3f", x"418f0244fb74a9c6", x"abf42421ff8e85a4", x"c7613ea130fe6ec8", x"5f95bcc55c9191ec", x"1b310459ec119d38");
            when 21496466 => data <= (x"e36bad6acfd01037", x"9407d5eb65e54ed6", x"000b6aa73c899c96", x"3aa458a8d4a50fa6", x"1c5ded6167d4112c", x"fdc6e42b7cdb2206", x"24a71d471b999223", x"4df2e6df50e52278");
            when 2620782 => data <= (x"26faa3c8aa77f411", x"c515fb99f5c48c2a", x"7210f12a82139268", x"d5c2673ad19fa8e8", x"99a38ece23d223be", x"2eb57db68c2f039e", x"e58a68894631c031", x"9b9b0e056064bd08");
            when 16788284 => data <= (x"a67e37787ed886fc", x"eedb1ac0b1248790", x"1ac69dadbb7fc400", x"2e8342d345a703f0", x"8502467e70699471", x"077a767d9f02377d", x"dc42c777c201f184", x"e3f9d99a089a26ba");
            when 5992343 => data <= (x"fd29fc9979091eaa", x"63cc020a46fbf256", x"1767acef81c856bc", x"67bd255e9b26627c", x"db6464954d1874f0", x"e7f15ae905969bc3", x"9e3ee253045803dc", x"3e97c5342c22d5ec");
            when 31866755 => data <= (x"a18f3c470f6d1705", x"65529d0211cc0c3a", x"e5f305ef9ca253ce", x"14cf666009ed5a0e", x"06e52e0e9bc97266", x"776b5e68ee56c653", x"8de47a4fa140de13", x"8740d840872c0d15");
            when 28717281 => data <= (x"9325872e386c1f6d", x"d8912419fb5a9ba4", x"99229b9f67248d6c", x"f065fc0e5fdc9422", x"e03374f845cc48a3", x"cd426130a0d0ed03", x"da21424a431961aa", x"1588ed7e5765b097");
            when 19945323 => data <= (x"e74edf6c6d6f4356", x"4aec69ab8a18e30e", x"de30cf1497345d9a", x"43ed86620a40e1b5", x"2ce7a19ba63a8214", x"e58cce169344fb5b", x"1f09ec17811efc2a", x"39812d1a089cda6b");
            when 23866769 => data <= (x"95917ae576d9009e", x"95459fa3f1310b81", x"a12bf0e5bb22a100", x"ad78fdc6f3e90e3b", x"cc05f1d98ccbf8b3", x"d50cea9376030018", x"acde3f5bd655f24a", x"b3c146a80d9bcb00");
            when 33658634 => data <= (x"5bb4277c5a418fa4", x"e0b82b6c1a14f09e", x"cfb3faf569d7e2f2", x"4e29cba5e0fd8a4e", x"01f0c39fb5af0e54", x"781f16520994002b", x"068603754ec6e3bc", x"61385953ecfc9c6e");
            when 3074756 => data <= (x"7d03f8f2b707c4c5", x"9bacbae5750b9c14", x"b9d6084a6af9a12f", x"15be56f73f8c716a", x"1fbd11f608fd1984", x"51e1c6fe4a4ae207", x"e5ed99c49b557c92", x"c8008030c11c1cb3");
            when 14177820 => data <= (x"d690f76862f39f49", x"99e7f28f26239af1", x"068e806657e92799", x"f26def05bcd447cd", x"8bd33adcfb8c22a1", x"07c6164aa42ec373", x"34b916989234a8a3", x"9e6359c1b6abf497");
            when 33404776 => data <= (x"107ec6edd1a85592", x"634dae5b0e222cb3", x"45b8c4ea9337c935", x"cbad70a6f5298280", x"8b6a726b8a89c5f7", x"818c8b175f74a059", x"b43126873f19a16c", x"9e75957d70244f78");
            when 10024149 => data <= (x"abb2b142464e05b1", x"ddad9cb4a2d98113", x"932a03293b9a0d42", x"a99346c3940c951a", x"1630cbbde28889d8", x"1cb50cfeaa6e0ad0", x"134a65d65163d4dd", x"c44f62e848244927");
            when 20174534 => data <= (x"9631f60f20624521", x"3b9e5d093632523f", x"2a9c997a0a9a3e01", x"dafde90e891ec12c", x"658fd1bc8972965e", x"46889b9885a53315", x"0c5074ba678e49d0", x"392435a5306950fa");
            when 26325676 => data <= (x"38be674f6290b130", x"269b03dd97232d92", x"b4a9d79673a28679", x"f0c8adf8be563dbd", x"3487c742019a0eb1", x"649daab2916bbdcc", x"2bb9304c6279d714", x"827a3ead6ff77e52");
            when 25150824 => data <= (x"6f3965cdeb8d2986", x"e2ccc2d7225753a2", x"b454df90fb7da504", x"84d164583ab72df2", x"449df2d1a69262b7", x"96063b3cf34fd5a1", x"14687d8210d3dfaa", x"674506933f58f54f");
            when 1459025 => data <= (x"b775c0393c71fb62", x"cfd38c91ba76196c", x"d0e63acd74708e5b", x"f8f3baf65db9273b", x"e3e8e54796c79370", x"6f1ce65dfee571ca", x"9dac3429b3c2a56f", x"cc52785abd18161b");
            when 25156749 => data <= (x"ef68443ca67f738d", x"81a60b264580c812", x"9e65213377662c45", x"6c5f943ee457a153", x"f2da1b8f221b2103", x"5ffce24025f98aff", x"d7df2244d8624771", x"ab3d3df4d1a2a866");
            when 29018369 => data <= (x"73fc05de679fe13e", x"be369f953bea99f7", x"3b9616e9642fd79c", x"a3993690573dae68", x"216334293e0d53de", x"02c5237b9eed700d", x"a82b9a007bc09ccc", x"c86c52b0cf965cfd");
            when 18678645 => data <= (x"ea177907888271af", x"864064092125ac4a", x"b5a6e3b6f77c0a39", x"b71c0aecb7c8ecd2", x"dc1300277a4477db", x"dd127216fe8f0cd2", x"35c649a181555db6", x"d0f92ec9990db444");
            when 19170358 => data <= (x"0471ebaa1f455fb6", x"db9d71573ba297db", x"6046d5f2301bbde4", x"29cfae5171ab3b9b", x"c2ce66cbfb26a1c7", x"139f7f8f1e36e0d8", x"4f02392966478155", x"423d92d77c509299");
            when 3991041 => data <= (x"f41c22905798edb9", x"add39e8cc4ec9de4", x"1417096b125ccce3", x"2e7949f184bdff11", x"67bc92f78e351feb", x"8acbc906b49979fb", x"71e1e33cf3f9b2a6", x"0b37c38d1418a039");
            when 11548237 => data <= (x"89582a56e2f523e8", x"1b44bea8dddad6e0", x"1e744d9052c62275", x"7ebb7713075a3538", x"437acb8387a614e9", x"0d8af1cff777536b", x"2c4930cbf4b3faa1", x"a1dd5d84765f61ac");
            when 19144511 => data <= (x"d5c2cbe262ef2f30", x"f706554cf45fa0c7", x"a287778c2fcfe69d", x"cb96cb19941a5955", x"5792af3c045a4cb0", x"d991b76b37438e3d", x"cd22a7f14c99d0b6", x"bef6e2da2cb22b44");
            when 17460052 => data <= (x"a490685de1faaac4", x"0f67a9b21198db2f", x"207660c1adeaa79f", x"21afebce5d3da8fa", x"8b7616846d3dec90", x"fb15ca7ee60b9c78", x"bf686cbc8d0c7259", x"437af577db5f52c2");
            when 28286121 => data <= (x"bef51f33f52ccf34", x"73883f389a51309b", x"57a21bde4873fad1", x"0031b7fda41b8e93", x"0b8f6670f274d342", x"b183596dd34f7f2c", x"cb029d6042425ee1", x"1563b753d35b3759");
            when 27251065 => data <= (x"aa817234bc3d42b4", x"c6394a7eba25bd62", x"0e23243e8923c361", x"c7d034cfbeeb91f4", x"db4d51a869e39e69", x"39bb836b3b634641", x"d14458df207932ef", x"0c2f9d72aaa13c8c");
            when 23193170 => data <= (x"d655c66a3d9ab66d", x"c3436b58977239e8", x"2628c86bdad668ad", x"67eab23d4b9b8683", x"52a6a840e4dcce63", x"b2253cead5343265", x"f51b330dc0ee67a9", x"277edc9c93264b69");
            when 25202224 => data <= (x"92bf4767bd85ef5d", x"9a13a859d6a647ef", x"4074497e7b6a918f", x"6551fbc7e0fa5b5d", x"c26e927c0d737e97", x"a2207f0f73aebbab", x"a8ff392d5ee65a9c", x"b6ce166901382076");
            when 32015209 => data <= (x"f600aa811f8a8808", x"c77d7395d850e4a6", x"333f5d7247776243", x"596358791f5dafde", x"e5ab43b5bd15b169", x"9968654f145a38a5", x"da3241294bc0333f", x"782e8ed623ff2ab9");
            when 5000641 => data <= (x"604ce6f8fddeec71", x"6de8d1aa02561967", x"bd6ddfe894cac8d6", x"ceb9d894561295d8", x"9f26e8d34c7c980f", x"635fc4d56def9831", x"82ac9adc9b2925db", x"a5bddf501004bd86");
            when 8979880 => data <= (x"9491ca1d13ae3a46", x"4702283376136033", x"88607892173b09be", x"606e86dcfcd78627", x"20e2ece74dda70ac", x"67c8f7eceb3bf911", x"a40847bbf8646bd9", x"4945edcc668eb834");
            when 12831880 => data <= (x"d3272a2c7f3d2aba", x"9e7e5728cfd221c5", x"9470c9ffbf686a38", x"e4123222aa1954d1", x"2963d2fb880a2a44", x"3b012f06449ffdfb", x"f26f520a198d663d", x"39ba172aceee5da2");
            when 31504630 => data <= (x"398aebced66dd050", x"2460c945509c3fe6", x"77cbab64812320cd", x"fcc9edf38e7547fb", x"0aac64bfc905d170", x"3f573b0a5710337c", x"766b69453518248b", x"274b7a39d51eb123");
            when 2480194 => data <= (x"ffba59412cca6fc9", x"2ac4f29bc13252ae", x"49c095bcec7c6791", x"961d8bc7c0109044", x"e86eea1151301db2", x"179c6b7b16871133", x"db7ae754f36c6905", x"37eb3ff0436c373a");
            when 24026974 => data <= (x"1ad064041ed16c85", x"d3f32c7836ebedff", x"e53f8ff6cd0bbda4", x"3161702dba024b09", x"338b102aaa0fcc17", x"96f25b402e166471", x"533afab2f84bbd04", x"fb17bd27a6541289");
            when 5307368 => data <= (x"529afbcfc97d9480", x"f598ab38ca2821ab", x"ff37311490aedde1", x"8d98604a0d7087b5", x"fbdd9df49c77e256", x"bcf7d2d07e5d2710", x"61f7fd1d00c83af3", x"53731d556e5229d8");
            when 8981734 => data <= (x"cf35c5e88178559b", x"169994c2eb00ffad", x"ad1e87b2b2ddacd4", x"c3a658f9de4bbbb8", x"605db48bd0d0f486", x"4f7dbdd15c21a6ad", x"df9e8526e44fbde8", x"953a191a0dfa4389");
            when 3267692 => data <= (x"e52d65950c334a9a", x"3c8ed37c6203f9ff", x"f8df4b3ac0897578", x"295e8e83112d36cd", x"82e96ac88028196f", x"bf7358fbdfcd0e16", x"e4e90927c2ef1db1", x"b53f8fde6ca68333");
            when 19045659 => data <= (x"3c3344c2f2528ad7", x"aa8d059f9849b686", x"4c4074e2db276053", x"eb4266e7999cfde6", x"1049a8f61bc055ef", x"c53c86b496ae21fc", x"6c75f57799ab29a0", x"f0fa4009359ab622");
            when 8774824 => data <= (x"c4b8b4bd4e3bf0b7", x"722c432e64374364", x"94a2f590a719c73b", x"a651e8a6e67eec49", x"0e371768f02c7d6d", x"58e0ce694bc6d6d6", x"92c2c7d9347de66c", x"f88d389d4250ea95");
            when 33694373 => data <= (x"5fe0e9c59e362a12", x"c1d22d207ca30a30", x"4ddf79467e730f25", x"811b53c04fe22dc0", x"cb57ea8ffbf05309", x"7d9a1df834e25ad2", x"3520571c0951f639", x"7c4e57e6d279c55a");
            when 28734644 => data <= (x"fa8bd9b58f9a200c", x"aa00c437e30acd86", x"0ba223c77bcbb9ae", x"707c0b132800b9a8", x"839b4ae0b46d5157", x"cfc299c735ee28b7", x"e18d965978e61114", x"562de7c58191fac8");
            when 11814773 => data <= (x"9e0bb08b45d49ba6", x"f3a47ed68fa487ad", x"24796cf38a3a5d98", x"0014297dc95ddc42", x"6ddb7f4de8e71535", x"2e8100ea3a2a204c", x"f5d024269e383b49", x"e7fe7736cb161c6a");
            when 14022334 => data <= (x"d4f409b27c1efd6d", x"541702c710db3fa8", x"442e9f708c56d9bd", x"4b95dd327032939f", x"1c70da0c2d4bb70e", x"134cce9ff5ed2483", x"8de4ddee54899c75", x"bb25234a65b690a4");
            when 11621075 => data <= (x"92a9aa306609203b", x"eee406e5f2407686", x"f7409de1cec6e16e", x"ce9737f183c3c461", x"154cab4106016efc", x"3ee8e75f5df72b45", x"70bc18ab6732a5df", x"2aab906b5309682d");
            when 9311510 => data <= (x"1a7def93b8ab3f3f", x"d8d371b4549e3e4e", x"36f1112ca949c648", x"3c1cb7039b1caa0e", x"8a64b2d73b4b408a", x"4f29e6cc92c8823c", x"7ab95a8dd9050275", x"c147cd5cfbc9ab5f");
            when 20196473 => data <= (x"981a33e2178f82fa", x"28871079e0ecfea2", x"c962be26daf3f1ff", x"01a9016be01b1bc3", x"06862be073ce85a7", x"fb5c158089cb8e4d", x"ec814a0275117913", x"7e42456b3737855b");
            when 19261382 => data <= (x"5c19f246551ee088", x"99f9eea6c55aca48", x"59b5ca6b34116f31", x"bbc58d7819bdc2e8", x"471beda14a342bb4", x"ad007566f06953f5", x"0acbf8fc56617b23", x"884170af4cf0bd61");
            when 8577314 => data <= (x"4eca45843bd3c475", x"4dc77a79836b2e4c", x"ff1ace9d5068572d", x"7854e0afc044785e", x"4beb2e430bb777ac", x"3c5c5fa101e3ed92", x"57c94ba9b2d43f89", x"7498594228bc2bcc");
            when 33283216 => data <= (x"acdab15d19e07ace", x"f837b5d7827cc49c", x"7f43203f54fb2c7d", x"b741f00dafdfa325", x"74cce59784e3c630", x"4a873599e460a536", x"5e752f7e0f73f05c", x"3603ec353cee9105");
            when 8646633 => data <= (x"f7323c92f35c7b57", x"9f217936f126eec2", x"005c327e26e9cd58", x"8498f79519dee218", x"7d3086089722b960", x"09ef95e251a0a132", x"31567588ad5f8860", x"06b8c539f0f2c5f1");
            when 6051270 => data <= (x"a6d40e875959c10e", x"dbb99d1c4b69c527", x"361b970b49d51d98", x"c1a314fd6bae6759", x"d0deeec2e10a3216", x"fe648daef633f643", x"882da25cf68819d2", x"33ca98189547ea37");
            when 6598457 => data <= (x"968ec26f1ef46952", x"e37264466e15b130", x"655f2fd4557a7e34", x"2756de05cff9042b", x"b727968f46b09e6d", x"e77a355b7481ba0c", x"7b1d7a4fc5037298", x"55c83a5b7d30231c");
            when 33213262 => data <= (x"db58d0db506eb528", x"14b7a9ddec47521c", x"824a65489b5b6d78", x"9b0ab78bc296f914", x"5809a5328353fc5f", x"2439b0a87d554cc2", x"9eb3c7c034a2d405", x"4480a3636b4440a3");
            when 11597534 => data <= (x"c46b774d3921e00f", x"bef732041236e3f1", x"f93a5eae1d4c5de2", x"72eb5b6da5d49b49", x"691ce5578b714810", x"80489148666d7d80", x"3072a3fa351aad45", x"4d0093f92528b680");
            when 10563259 => data <= (x"8329063f7bfbce80", x"6d4fa8530f1bfad2", x"5931ff8540c3da7f", x"c93be13896c7ab91", x"5966355c4c9d5bbb", x"4e4ac5828583c3ce", x"7fe7d80dee260999", x"829236d1abc20048");
            when 4983223 => data <= (x"0acc33f8d7981c16", x"6610654751570f77", x"d99b73cc06055e43", x"8ea781dbe6da950a", x"d5149052bd5978a3", x"9aef053fa1db897b", x"e114ab1d4a7e4101", x"a10f65a3cde8108a");
            when 27865962 => data <= (x"305e7b23415504df", x"c00e5c489408272d", x"1a58e112f3c3d6e5", x"5e3bfe5536c623f0", x"2ffcda35138542cd", x"3648e34f43b10ca2", x"b4fc1d078ad340e7", x"e4c8cc2ce69368ec");
            when 8165081 => data <= (x"9abd5e71fc413105", x"2bd930e85569c48d", x"39abbb515fedb6c5", x"8c182e1f59cc3668", x"37cb84a3f72ace29", x"1b11ddc70718257c", x"6c0c0f6977d1fb36", x"34ad17f71abb67b5");
            when 11748494 => data <= (x"b0fc0101ba06c070", x"f52dadcdc25b0361", x"1bf50ea32bae0bb7", x"58e40341b149d0fd", x"9af3c58ae708d803", x"bfc6ac94b96db87e", x"015cfdce7addb976", x"85121266953fbfd7");
            when 26046522 => data <= (x"c7291a8579d0d121", x"28612b51a15fffc7", x"8cb24a7755cb8ad2", x"f8a970f28c68e70c", x"62939475780c8ecd", x"a0b70814d0550545", x"0e4126ec792cbdc1", x"b58bdd1c37313337");
            when 4142608 => data <= (x"77adb377cd064c20", x"4849e1f891bee306", x"c833e31c01f065d9", x"3d9ffa0ad524bab7", x"494f74f93a4219b9", x"b7af62fd17289283", x"dceba013fb1b3898", x"319ae95f62e25d75");
            when 3500873 => data <= (x"e31ec3e9f2458de5", x"2513dcda97822c4b", x"1f8aed36f9a48c99", x"ca906a2d01ec19d8", x"949f7839e0d508b2", x"4f5a59664465a4e6", x"58c62115c380a242", x"5925a1c324e0f4ec");
            when 5336778 => data <= (x"6616520c85ea0c5d", x"3b7e3edcd9473db5", x"a3a8b5d5c0621c25", x"5c90945598524ec0", x"121c5c1507d2bbe6", x"16320374f6501cd9", x"ae3ddf5a62886d92", x"c1567f566f02b9c7");
            when 29586842 => data <= (x"50403e24fca4c33c", x"48ae2398e0331580", x"734b0d5dc88bf113", x"048373e21b0191fb", x"dacd63139d62009e", x"8e594e485cb9174a", x"e2968eb0ff780ee8", x"9ec652c5db6014c0");
            when 7747280 => data <= (x"de49b0865396c757", x"c513a078b49f6556", x"83fa6d987581f8c2", x"5520e77c9d20ac9a", x"a5fa39bdeeb8fab3", x"554506fcc64dd244", x"2778fe3c75eadc84", x"30e471b8eea0945a");
            when 5067973 => data <= (x"491546fb5eb9ca6a", x"f008df0ffe69f45e", x"c6c415134e9396cd", x"e29f2ac4b5a33e2d", x"83cc9753233e6065", x"7888d3110d4331d9", x"679204fd43bd69e1", x"26038d0a4dfa5fbc");
            when 20101974 => data <= (x"5c9b343fe16a84c6", x"1020a05730988514", x"0269adba82f976bb", x"7980143e4081fd96", x"798a0323d05ae696", x"61ce208e765d7108", x"e3298ddd0700b14b", x"f9b3aa94bf8a00ef");
            when 14061424 => data <= (x"9ad36a8b49ac7565", x"6075fee6984d4244", x"79319f6d86cee727", x"a5835d34087badfb", x"ad0bba18cb1c0bf0", x"a1eef6fdc2e16bd6", x"f22a6d73676d3d5c", x"6fea741ed5d96ec5");
            when 30164527 => data <= (x"305f58da84121863", x"89ca13c6597f5c80", x"5c2911be4ade3395", x"e88cdfdac54b6094", x"9b424a38dd5dcc87", x"c95f71eae5fa9dc3", x"39b1c7b01293d177", x"6a0f5da8000a64d4");
            when 33478049 => data <= (x"14e146ad0ef38179", x"627936f6557242a2", x"8fd632436ceb093e", x"70dbf60ce8e0949e", x"60855c5069409c1d", x"29812589e53222e9", x"807b02c7d2f8d354", x"6838d5bea33586c8");
            when 23602364 => data <= (x"1d4a1fd3a6c1bbe3", x"70946bd1965c16d6", x"15c733d1f4e1b6d1", x"16b74e772ee6cc18", x"21e3af6eee088338", x"fc7064d692e1e3c6", x"00ad0836f8ec07c7", x"60f74f6e165f7e8f");
            when 4488307 => data <= (x"3780c04b8e995473", x"2f1636f394fdf894", x"7e78d79e4f23fc71", x"8665a106125e3de0", x"c387202df3bf3b3b", x"44eacfeb01aa4e1c", x"1e01425972baafba", x"431ec391a37d72c8");
            when 3958282 => data <= (x"de8aa9ef048eceb7", x"4ece358d4eed2916", x"14def747559efea5", x"51aaa13f8d60df36", x"1306de9127f87df4", x"ea3710971847c76e", x"6a87ad6490d44c45", x"7dd35480ec627a2b");
            when 11011632 => data <= (x"32c351ee17729a1d", x"3e2194fd128cc177", x"c512507eac31b59f", x"a8b0e0bbe88ab442", x"5896167171d414a3", x"9e4282c8bea23569", x"2aba15f6fbc359f8", x"64bd4e1c1bd22600");
            when 2091616 => data <= (x"de0b4b71df27ed1a", x"2937e0d075d9ce46", x"30798c6fcd84fb68", x"3962b1a096aecde7", x"bd82430e36352f11", x"457a6d7f34240d1b", x"a9f58d09f0b38ff3", x"7a8172727d64ae30");
            when 32228870 => data <= (x"aa06fd82d2bb3765", x"333aadbc541d1444", x"c454e43e939da9fe", x"ed678967935c03c2", x"3884213939cf50dd", x"b5e9749a03bc2355", x"11f54d606c8b4049", x"573f3bd2768b72af");
            when 31176430 => data <= (x"ce402f6fe57ee810", x"d9acbf1700f4077a", x"f709856b51e02705", x"28b69d8331f66a8d", x"8cf4d6275cc59a0e", x"4df3e01f39346bae", x"8ff2e84c75def292", x"ab95f18e6bc054e1");
            when 15444913 => data <= (x"e649df53f4e3e41d", x"e75fc931e662be9c", x"e14ef70d56447977", x"ab46ed6ae702113c", x"1c003aab370076b9", x"69868a592bb50b11", x"de685695f07139d8", x"c08edbb2eb48d1cf");
            when 32404185 => data <= (x"b7d40257de4cf107", x"fe00b4fb9d152711", x"089229fbd6485b1a", x"29507433de2cc5e2", x"26eb378ec8a4ed9e", x"ee42c4c4c2ccaebe", x"3b90cfe600a5b50e", x"9b10856a57213c0b");
            when 27260820 => data <= (x"526c4df65282a66f", x"682c37c5547b4cf9", x"87677862e65f9038", x"b3ab48c63281438e", x"aed7ae03e498173d", x"66b3a7d91158f0a7", x"a0c9152a9d0f4a3e", x"ebd7d7ed439a604e");
            when 27830853 => data <= (x"4a441941b5d57c7c", x"590287ce810cd6ad", x"fbdf850f086ede66", x"4730630757868fa3", x"91cdfc92300cf965", x"515f6d8be5d24493", x"802626952ed1324f", x"6b49ae3e131f1f77");
            when 17432196 => data <= (x"56d6912ce2cee987", x"dab0492133f92eba", x"58340df8b9bd72b8", x"5adbc3b4b572b857", x"ad0a62941d996a9d", x"c18395f7303fa055", x"4697389f00f80382", x"d86741404b4be603");
            when 1269323 => data <= (x"d8315771cda92925", x"86c29c6154943707", x"a8197f8cf22afc93", x"8ae195eee443c991", x"61be34ab79475a86", x"ea2ef2b0dc3e8d8b", x"5266a1b3281b066a", x"e8e8ddb02c39677e");
            when 14436397 => data <= (x"841c192f810a19ea", x"232383f5781d0a73", x"e91ed377f79ad5e0", x"eb2d63ff323ba471", x"8ee909c8fe629619", x"0518e4e6eb89a633", x"4b67cfc8fd1cf2f5", x"cbfc69d30b2a090e");
            when 14869308 => data <= (x"2970823476579ffb", x"6e061de1c9edf713", x"0992aceffba72593", x"bf813abf2da6fa88", x"cdd2d3964077b2ff", x"2fbf0589f13c6c62", x"da0e49e0d23c148a", x"7db076de0065b989");
            when 3177139 => data <= (x"2b24bd1e59903225", x"b3f18beed191b94a", x"951048b78bfee499", x"dafd3dd25583b7d5", x"bfafe1b71e69d3da", x"71b06b8ece041bde", x"bf556d568861c1fa", x"74b5d22eaa1651d4");
            when 16116697 => data <= (x"e5a02119465338aa", x"8362109da39af4d8", x"f85f7b43c78e882a", x"fb0b562d9d66fb19", x"2085460b155082cc", x"39bcdba07d0b74b6", x"2f7c3e1874b80108", x"3295d754c56823fb");
            when 7821756 => data <= (x"145dbf5437431f55", x"b5f3226bad5f82ff", x"be0ad9994b15fabd", x"87a797266725c467", x"49a790f8f9fe59ef", x"dd3d46d1857c242b", x"68904d80e4aca6d9", x"40de337a18cbf3c9");
            when 11378021 => data <= (x"eda556138825904c", x"71f916139a621f83", x"cf1b0c706e663903", x"6e4837d4c77c2c87", x"a0f20ee8f9965115", x"54cc04fc60573705", x"667633577e55274b", x"5199877eeb6bc3db");
            when 9537049 => data <= (x"5ab353d4f4e039a8", x"53b32b62b3daf274", x"9cdef176702852af", x"c65c204121e87c31", x"1b879dddabec4917", x"5051c40bf1228378", x"0ab7908ccef5cff2", x"574415db6c51deb9");
            when 17086092 => data <= (x"06921d4b287ec23b", x"100e9d0c4e78733a", x"b179f6e102da801d", x"b08b210adbe333a1", x"c6d52c1d953fc714", x"495f8657b8b18eef", x"a70b28133375c81f", x"9ffe2675467d0c55");
            when 19993180 => data <= (x"d13141d030739ab7", x"6e40e03c3b3248c1", x"6d78b2374b1457d9", x"c2bc79fca86d9740", x"5f92b566d0350ef9", x"b98557a7907a5bda", x"94880f4e9323dd1c", x"db7943c94bc7705d");
            when 31615573 => data <= (x"f46bc1ce95d2e684", x"d227ebab9ccd3f81", x"ddd3e8efad83282b", x"690c956b1bda822d", x"d3e37a42bfba6786", x"35ab8fb0c7c8262c", x"85a301e00c70e386", x"9484e40febc70b52");
            when 8633566 => data <= (x"b887f231473c5ed2", x"6dcfed8660c288df", x"7e37ca4d73206512", x"efd4964792229a22", x"6c67be64f9cb096f", x"82dbcff659f6de15", x"f045a0290c4a1500", x"1ff5f908cfa52926");
            when 12996642 => data <= (x"8ed8e90765d34168", x"527958dc9a07b01f", x"eb110576cc991dde", x"13f27fc593547608", x"6dbe151ac4322051", x"b70d417d2bdf525c", x"ca1f575cf7ba428f", x"9e2383b9dba44496");
            when 27602290 => data <= (x"f77264e9b0cc24b6", x"515ecbaa37a87add", x"f79a44afcc4c817d", x"ccc787013fc457e3", x"442c407e03146d61", x"ed54034c765efc7a", x"1ede218ef03c8bb6", x"e5c1347be4660fc0");
            when 16854902 => data <= (x"80bccacbe8529eba", x"4724fdd978f9106e", x"87408e9a153204b7", x"f375c08090398dc4", x"b3cb3e7bdfd641c0", x"18ce5bfd72bdb096", x"4b8a68e4fb43010d", x"610ff1fe684ca92a");
            when 26140997 => data <= (x"1f026221baf64f11", x"07badb2fc665104a", x"68da4a09d081eafd", x"4d6050d1c327b222", x"e09f63db09ed0c2e", x"8b0ed38c0004600d", x"c295b4e4dda39e5e", x"c404c7e9849a1ed0");
            when 22208521 => data <= (x"f32644dbceb19bb8", x"306f9c40c1e5a802", x"bb6eabf360ed25a0", x"b0dcb2c3c930c3d3", x"fb6cacb193bff64f", x"8c1d37e0d8304cc8", x"be13263f73f7337c", x"e3ead5a8bef7d554");
            when 7215655 => data <= (x"f62b5a199accd8f1", x"628f83be83ca545d", x"a8711218a624e064", x"c45a04920f4243ad", x"cb5562e1ecbfd524", x"d1440324211e5ebb", x"6946a6dfc67e35a7", x"853fc0d3801eb0c2");
            when 30628092 => data <= (x"ffd79ca223025200", x"d9059df3c16506b5", x"f24a3a41b5790640", x"c907fe5a31f0b65e", x"ca2c01483b0462c3", x"aaa5627d3c091515", x"3278dd01ba27e9a3", x"23f3fc11d6139461");
            when 33539411 => data <= (x"59569029f5cfc0f9", x"5a93d0014f6148b0", x"f438f38bdbf2b848", x"8e911ad683c2fa22", x"05fba5fbe516af92", x"a33b65d3cc0c49a1", x"910d9ec699f0b0da", x"1abdc7de1b74df0e");
            when 32527876 => data <= (x"cfd081028b030b79", x"98aff8c8c1b45899", x"856b6200284275bd", x"d4f8a5365581fd14", x"bbd8e0d86c2d597d", x"1b92f847655bb7df", x"a107194aaa907942", x"07e79ee7a9ea7114");
            when 27329874 => data <= (x"a488b066b0c55519", x"e71b570580247072", x"e29dd04f2a890793", x"72cdd10f9160313f", x"9502fdab2059de6a", x"2f0193cba5f5728a", x"5ef5f6dca80b6775", x"e89745a4aa961abc");
            when 18609595 => data <= (x"89d69c452976056a", x"df493a3d650dcac4", x"cf8f3ec97a76476c", x"87f55d77ecb2e6f9", x"f1feacfa3b99176a", x"831c0cbb4f9ad08f", x"73affb2c4e04c89c", x"1a99f03e55d8d2a8");
            when 22157980 => data <= (x"3d4b0f3ece7236e4", x"f7a4c9dfc72f8b4f", x"7014f80cb1337d58", x"094d0cee3212fde3", x"917e8c006e9ad2fe", x"49fb6075d695576c", x"d2072fb066172235", x"ffba3a218336d138");
            when 2200489 => data <= (x"d2fe139044827621", x"532209d8153cba9e", x"4d99718231c6efe4", x"3a23c8d659685175", x"97dfba5e94eced8d", x"d7fa9eeb50f5eff5", x"76e6184e14739ab3", x"5bb8a2836aba0b61");
            when 2959208 => data <= (x"6038ca12acf4c1cf", x"0b8dd201d3d85927", x"e29c955e406f3c7d", x"899648d30d5f920d", x"b95aea5a0d13e367", x"16d88e0a44ba97ee", x"cfd1c1ce71166fff", x"7b6e3d4676c478b0");
            when 10424802 => data <= (x"5b9013413115a309", x"400fb50b9145ca57", x"ed64593b4cf9401d", x"0f9031ecf1b1b7b0", x"aa6b33cb44c223b6", x"9b459f2dbc98dc73", x"c649c7f1890aa834", x"911cc806468c55c1");
            when 13850383 => data <= (x"c7de1a00452a82ed", x"d9b819567766a067", x"55bf7337662f07c0", x"94e8c5946f2e1ecd", x"30677e747d297d6c", x"ebc2f51c19690567", x"725603019b96a4f2", x"930704bebbf38d79");
            when 7782465 => data <= (x"ce0a9055a8259797", x"9d3ec5d0868a47b2", x"9b4162255a44a466", x"223edaeddda3a5db", x"1960be68de1946ef", x"43b9a993f8a96435", x"cdfab9ec578c1266", x"db3fdf2ffa696b02");
            when 13101847 => data <= (x"d46bebc74155da63", x"bf2f58fcaaf37061", x"e79ddd5a3f3f3c32", x"04d638160ad5c8bd", x"416d4479007b2d4e", x"618d2367a49344d0", x"1454c3c3b49c939a", x"6e162e722dbbf485");
            when 4984798 => data <= (x"2a3405719a923526", x"5fba3cf9a5f0eb2a", x"36c3313fdf6afea1", x"09a0c45984f8419c", x"1cdc5bbc373b2778", x"d89a57f988a3b479", x"57663f8151353278", x"4487c03dfb44a760");
            when 8406004 => data <= (x"5630478721ef5e78", x"af1ff9b8bf1014c3", x"434814f9a372944a", x"d8111f91b2227a2f", x"d00293f73f00cf6b", x"5148537a25a7316d", x"f3d8e3e88d64b560", x"16ba67878497bbf1");
            when 10888502 => data <= (x"1529ad76f8f3beca", x"91b2c97b5ee1ded7", x"3a85e8037c9a2e86", x"1bde1d50aab3f06f", x"552f649ea14192d9", x"2f028a54937d5bbf", x"f8cf3a8c7a28580b", x"1d8e30adc669b9a3");
            when 11444496 => data <= (x"9e13ce2820f92bcc", x"078d4788e890091c", x"f93e6ef2aaa14cf8", x"3ff85e28aaea026d", x"68907cd199b78850", x"f8d234fef7b88f1e", x"e0766d3fa7e1d7e7", x"67d8c59566cc04be");
            when 32898339 => data <= (x"85f55125a64cd5e1", x"608cb12ec09c157e", x"61fa1678550f3a8b", x"9bacb955bea5ca3d", x"d59b076689d5e512", x"0537aab7e88e3ab3", x"f226c15bc5f4cca6", x"f08fda1d823ce984");
            when 29191067 => data <= (x"09bce815eb2dcae2", x"a1bb36dd898b2f59", x"099c21d886f131d0", x"68bae08209025377", x"19ade4e5777d3c5d", x"0d54d93e20475eab", x"ef35bc3bc5f6a0ee", x"0d79daede1792573");
            when 10027977 => data <= (x"11283a2a0bd5cd0d", x"bdbe4e843a80f071", x"a3596d15bebf5090", x"65831544e2f898b2", x"aa729f0e1fcc3617", x"e31f9edff5652aaf", x"3dfba20222d321ea", x"4a5c7b0e0e6720fe");
            when 20097713 => data <= (x"c6f0f24a5cf9104d", x"b029177726630010", x"125a03806c3b3499", x"bdbc7204fa3fe64a", x"0120999d156c0dd3", x"07a0f770d3647785", x"b67e69e014b645d1", x"a57eb93bd6b0e9c0");
            when 31297781 => data <= (x"6f29cdac4fb7db34", x"9ef1b03128a7a5ba", x"96d8ebec7d02eba9", x"119a71a8ddb7e752", x"095d4931bbb816fa", x"28c72dcf2a47a666", x"77af8d1732807020", x"7cc787c6e34a3120");
            when 30322146 => data <= (x"576c37e75ccd835e", x"08a7089cdcb46790", x"6cc92e814e49a31f", x"116cf54e5df02762", x"78b760183e212637", x"ea2fad0f5a8638b0", x"a5c8f73dc5bbcd1c", x"37d3d916c0f5cc5d");
            when 19121659 => data <= (x"b9e006acae470065", x"f42520fbccc62c2a", x"44a45c56124cfcaa", x"2b7568433c20a2cc", x"2bda18aee6654e23", x"233e79c3da09b9f0", x"6cb0e9681c299175", x"2ed08b4e058441a7");
            when 4157777 => data <= (x"95663091397c1aab", x"195e4694af14c23e", x"dca94e8a5c1e8ef6", x"13f03a67cad3e971", x"2702520fbfe837c8", x"6f5b2d82843f2e32", x"177c23bb7a459cf7", x"792e63f9dae0f65d");
            when 27910866 => data <= (x"b0ff25b1d9181b64", x"0262cced235296c1", x"517415a8064a0fd9", x"93d7222475a92a39", x"231abb0de07cad9c", x"0ae91a56550c6c76", x"1f98d2fea390de33", x"6954c1c790b9bfd1");
            when 28262854 => data <= (x"d38a645dfceca8fa", x"0c9a7abc58312072", x"c51b160066ba813f", x"7cf0242474e3ed1b", x"1e34ad367cd48bcd", x"7a06b4976570bdd8", x"1e517e236fa76f61", x"56ce0794e287b262");
            when 10473912 => data <= (x"3116cc932f42a283", x"be10961ffdcdd2a7", x"4daeaa3950e5d592", x"ca8e0a3f191a91cd", x"6ffcf0509c1916f2", x"c5ab5209d668e15a", x"f624325d3275c53d", x"987ba1342102b316");
            when 32159631 => data <= (x"cdba9fc4bb7f23b6", x"7d9fbf33a0b66633", x"a2cefc0399f59a8c", x"bc3f843fd7cda6bc", x"e8864639b465bbd5", x"1a1fe8947ff0f7cb", x"e6cbfdfca16e4a04", x"7196bf11c7f2599e");
            when 833739 => data <= (x"5800f041fcd2635d", x"45a1710e5e9a7c43", x"a16af9a580eae76b", x"a5331f0c2483b8ef", x"0af679c99349feda", x"d59c120f5c1b9d97", x"24e4fd1f05cf4094", x"f56bc186f552332a");
            when 7241640 => data <= (x"1acda60527c76a0c", x"75170a69cfcbba03", x"29e7b246ba2fd916", x"a8e94d1609c6a545", x"9fd0140a334b5c53", x"97e446df4adb3212", x"3809469cbd639993", x"eb8fe67753b2b0e2");
            when 20381423 => data <= (x"1d6b98ed4aa8268a", x"ab113cb52888cd21", x"ff7ada301865def8", x"464f6b4887180ed4", x"b86fe571dde13bb8", x"8917f938ca454e5a", x"007ef7f092d26455", x"c566808856875a4a");
            when 2439738 => data <= (x"c5e065759eee1c14", x"a543b1203c294b8a", x"9955784e5e86f44b", x"b73a1ebcbd593bb6", x"70cd9d3daad17f87", x"5263dc71626e8e4f", x"9ee56a679bad212a", x"a02d75da8220be64");
            when 20280777 => data <= (x"2018edb85bb13307", x"832d44b62ae1b2aa", x"fbfd31a3acfdd227", x"1af787c4b25459e2", x"de4ffff1bbc62e98", x"2606b09d49902b39", x"453bd9096ed77f99", x"f1c8834f3f23e9f8");
            when 30154376 => data <= (x"3da23a6592c51374", x"72a033a96bca0cff", x"1014efdbb8ed8cb5", x"b0ee266bd810412c", x"11650bd1b1ca5b5c", x"761a3d607722aef3", x"81af7ccf3866ea4f", x"3ed409914bbcd8b1");
            when 27031957 => data <= (x"92aaf6d90f9b96ac", x"103974ea4c376648", x"1accf8e5c96ecf8c", x"1a06f90304f33255", x"9290d063cf8acb46", x"0106902f06dd1bbe", x"95acfeb6c5f3c0bc", x"b1ffd4a5501a20d2");
            when 9096909 => data <= (x"d06f991f1babf452", x"0e1b700e1faade6c", x"f9a753e5025f17ee", x"3b4640b6cd680c34", x"8eeb232f7b1aa971", x"0a3df52a5a33ebaa", x"8e1d4ff1aba8d09a", x"aa424d7f422b07ad");
            when 10843268 => data <= (x"272e8b567ae8db82", x"8b02c4c2b8840eaf", x"0dc264e01b15a1c6", x"7be2e35bf90a4244", x"d5435e463ec3fae0", x"f75f973f1d3377f9", x"250b45a596f7ed8c", x"e6edddd37b5b2e4a");
            when 17069402 => data <= (x"ef7b3e12d8febe84", x"d27b7539f0125223", x"acfd309ae6deaa5f", x"2f105a8be0b1f44f", x"3127cebfe0c771e2", x"5dcf9545b73a196b", x"d6516e9059f2c0f3", x"50fe7dc387ba609e");
            when 31637453 => data <= (x"4f59e1e5fe563998", x"3012c2d838976d6e", x"b57a6ef9299d95f3", x"281afe7ea47ef39e", x"0849e6a2da2e7acb", x"97bf4d52017bfdbb", x"1a77f497a0e8aa88", x"e985cbbfd8906a79");
            when 9112194 => data <= (x"b017e62dcddf75c2", x"2946e9c2ae4d7190", x"ac73c8622c2f2ee8", x"ca83d45b53b9242c", x"c9bd23533e7c7ad2", x"3e999c211f756d16", x"772983407ced30a9", x"ab8893fdafebde70");
            when 18548279 => data <= (x"3e0e9e83c11b6be0", x"42c8398d2d12a280", x"99ed6d4e65c4f759", x"befbc73d0ec65f3c", x"4af8eb56a9326500", x"6d44c8d199ceef58", x"c6d58c0bfc18ceb0", x"d9adc7d3e126cc77");
            when 11812725 => data <= (x"2c481cb2a12575d5", x"52edd7d7e13cbb31", x"ef6c70e3a64214bc", x"9efc66a1ea71819b", x"a335ec5a151b1234", x"cf895a4b8ac18c8f", x"9a876f74d802a67e", x"e3f3ec9258e0d5f8");
            when 32583624 => data <= (x"7365c4bea4542b99", x"735b451a0cd4e63a", x"2f8cdc1a661f4021", x"c9daa9d5cc0ddb4a", x"8d80560da06acb16", x"a5a438ee5f5c4dd2", x"0325cdfa795c4625", x"1f3af20bdfd77012");
            when 28837675 => data <= (x"7f7e431db5835a6f", x"7906106d1943117a", x"dfa23bf00e885017", x"3b34791af65f21d2", x"2714a9c896d62c6a", x"8fa1ed351c4edc5a", x"34234932e3a4b3fe", x"d2d9740a32925e46");
            when 20852687 => data <= (x"28fba6f22be4c29d", x"250cc22ab690072a", x"b30df304ecbe74fc", x"27ca996e6ded8e78", x"ce1064eb15ea2234", x"c0ef96cd3f44c56f", x"42679d6458e36af8", x"c34a05d188380b01");
            when 19857182 => data <= (x"53f466a14be5b0f5", x"bbb30f80addf961d", x"edd0f2727572a01b", x"a0df1dfdbad83819", x"7e3f66b35fb143d0", x"5ca1070335257d3f", x"ecc1ee48b959274b", x"5563bdb190c3aa19");
            when 28255406 => data <= (x"b7cea75553345da1", x"19e590013f50dcc3", x"ff31a974f0429773", x"d9a5bac324e1b18b", x"ba8876e46aa0c356", x"94df6a6309535789", x"a7becd767c618cb2", x"29974e2f1531ffdd");
            when 32570887 => data <= (x"3533392b87a55454", x"7ac672fc8481091f", x"a89492eb604040ac", x"253a9dece98889b4", x"0f6f51d6233d0a29", x"b042c227b2bceca4", x"386796e3c69a53c4", x"3049c1e3a0ba77d5");
            when 33168395 => data <= (x"a841a9ccdf6c5473", x"fab8fa537e4e42cd", x"cdc2b413a07a7f13", x"701d797b8e737930", x"1d55dae0427d9975", x"7e1e6c74aede4dd6", x"66c539445c9be8d4", x"5d9787cda08e0dab");
            when 33470662 => data <= (x"33d000c32c9a7d8e", x"392b5a14c7731c7f", x"7eaf77cb343c5c73", x"3f43678b82fd4e7e", x"4ff8d939f00369b8", x"978b73a674b0a6cc", x"aac11a1ee43e1ff4", x"d0154605111cd1a3");
            when 21136762 => data <= (x"420eeba766196ce0", x"e813cc94aea2756b", x"309ed0a9f9154ec1", x"dbeed7c05e4209bb", x"af157e0a5be60f02", x"145d897ea00e85db", x"86c4739a01313614", x"029d222ff6a250d4");
            when 23780618 => data <= (x"70527938d1c32aa6", x"0eb2695bceeb79db", x"bd09f9954c5d35e1", x"30ca6b25359f8a46", x"1e1156fd61e409fb", x"2ded67708da54f38", x"584e178128d9f232", x"bd2eeb4e121f3d58");
            when 17885500 => data <= (x"b93b70110429d2f2", x"1ccb919ee54dd66c", x"96bc3fadab5b1b16", x"3c5713c712308431", x"b03dc55aa5e94573", x"e3c6aea3a0c7327d", x"13ef3044a5377597", x"944fc9fc8d4ba53e");
            when 21583212 => data <= (x"148695afddf573be", x"9a8a7905e4335691", x"32bbeccddaf37275", x"0f2a58ad42cc71fb", x"40ad48e7bf8f0ab5", x"6a8d5a9e21d7492b", x"56bceeaeae927d2e", x"ef37b9673c6fe478");
            when 4030096 => data <= (x"6bf7aa0966320bfc", x"de36241b3d14f6a2", x"2968fd7d81e07b2b", x"54f2b866b89b22a7", x"98aaa41c0e586cba", x"b77d28b1feeb16eb", x"6d625d9de3560a12", x"f361d76fa3c406c1");
            when 15876374 => data <= (x"a24f9baa8a959822", x"b65fde3258e4c39e", x"63b318321aa27298", x"65d7fad6612cbbfb", x"2446114fcf79d15f", x"583bcd48e4982e70", x"0e0ab3683d05e69b", x"6c149cc7d3213afe");
            when 15910045 => data <= (x"f295055cc077bd50", x"5d9b4c946cac92b1", x"8fe6e84600865856", x"c08c114a8dec30c2", x"92cdf9b3e688eaff", x"3d834176f8e0d7f5", x"174cd4adf5c6dcba", x"a6702f49fd4d62e9");
            when 27538283 => data <= (x"978629814924a763", x"47b3509ce0a12d5d", x"eeba84fcdff3eb3b", x"ed0136151d1ec81f", x"28e4abce6a7bc846", x"d6c11bf88ba0a078", x"a61972f5d0935b61", x"8571710114a129ee");
            when 23045310 => data <= (x"b9c393bae7eb558c", x"32dc100e363d3977", x"255387e3aef3ef69", x"cd8ce155f066f935", x"f61f887fc7e7930b", x"5745a66a54b526b2", x"505721c34e3de987", x"f427b21c68341a71");
            when 13955895 => data <= (x"2d15f90adbd60506", x"517b549a334e4c7c", x"59796a205012f1ca", x"cad7989105fb4d6f", x"a894e8ad7a28e3d4", x"55775cfbe3e98ad3", x"cce5a33431b38d00", x"2eed202315135b1b");
            when 4991223 => data <= (x"2e7b051b3e9795f6", x"0dff960ecdcfb36f", x"236aec4b30645c50", x"f731c86ed474fced", x"4267939c1dcabec4", x"da0cf54fa830900d", x"4011c9b1c5332549", x"e4d3b0f7baefee87");
            when 10348747 => data <= (x"01c39db4a16b6893", x"c6f5cd79c7725032", x"9b4d11e97a16bd5f", x"d68fc8ca67ea0359", x"ea92b5d462cc5967", x"35ba188e62f945da", x"115a3d30768cae5f", x"31a5afd1b553484c");
            when 20321406 => data <= (x"3d2f07b9adcb52d8", x"72cfca2a532e2856", x"617d9359fba9a963", x"9b4e4deff8e06912", x"a93bf2577ea66ffd", x"033f59a82ea1ca01", x"c4d9539aced8bff9", x"b50522a82a6fa107");
            when 14334867 => data <= (x"a3cf0119eeb36bb5", x"bb8510d0d24ba7f1", x"2839463d01509b72", x"19ae2aa2a7f238dd", x"0a7b329a02d615dd", x"873b36c1cfde3087", x"f0068a65825d2747", x"2286c03cbe07c1bd");
            when 33843333 => data <= (x"6f77ba81e72a2576", x"5fadee8826fc18bd", x"7b70072b256d48c1", x"1e63a54a16cf91fa", x"101e02a31b3a5c7c", x"511977d4d637bc06", x"716cde1ae36f1549", x"2042d0a0a054b855");
            when 22371103 => data <= (x"336e42796ce79f7a", x"6cecaf4bb33b6bb9", x"e6723b758b5f3c12", x"945511eb42d0105b", x"1227e2403296bb0b", x"08b217c5c9c08c49", x"3fee602272d4306c", x"5f0506f57c0cdcc4");
            when 2066122 => data <= (x"d90ea0d64a94c4a3", x"7c0862ef15847cf7", x"59d7ee4ebe5ab5b9", x"9884d713ac58780d", x"2dc067ede7a7f620", x"214f1ffff501c6b9", x"2e5ead119f2ecc20", x"94fb41d39fd57dd7");
            when 28263166 => data <= (x"57e25ee49325842e", x"81ed43e80d24a2df", x"304020bd5cf31d6c", x"ff86774a4fe7c075", x"44d96c65753ba79a", x"5b23379425aa2d01", x"579794f4c43f8e96", x"495ebc03e2bd9e51");
            when 32074158 => data <= (x"f61cd8688e845dac", x"609d5d30c08b1705", x"95bb76eac923156a", x"c666ebf2a2c5a9c1", x"25962dba78e7d819", x"2913ae45bd6c8410", x"966a78d8722ab883", x"e5e260cd6a8ea54f");
            when 8461196 => data <= (x"349883e0526d70aa", x"c9b59a3fb4a87019", x"6c022b8b71d4f8a0", x"8c912b66c89acb83", x"90527166419c9db9", x"d08266afbf6d2643", x"9af9654670a609bb", x"f7113881859b3d99");
            when 12566880 => data <= (x"2684a50c434bc914", x"7280d64d57dd208b", x"654a2df2125785d9", x"ebcf3cdc268a3280", x"377a979b2826ee7b", x"2b024caca903070b", x"34e7da7a509d6b1e", x"6d9982b6a092feaf");
            when 19173362 => data <= (x"6389f94bf9cabe01", x"97b85d6e07299bfe", x"17ef823a200cbb17", x"89f2579061859e49", x"8514afb9657631dc", x"fff336beb5d514b8", x"ee0a3652f655b6f9", x"090ff72467bf1080");
            when 3323384 => data <= (x"f2d6de3984d4e01b", x"ed20085d7f5c6878", x"64942859e7e2f893", x"ec8208e0d60a7be8", x"44271ac380b53cec", x"19f5fc8176e2be52", x"b468e98182bcd271", x"112fe4df12b1bf02");
            when 22873705 => data <= (x"8fff767d76c770bf", x"0b5dd687171bcbae", x"a9aa6a74a9dcd157", x"133cbaf0a7ccd085", x"f641a4b275ed5b95", x"6b6aaff81be1ebcc", x"5e6db7f853ded1ce", x"4a48690ba92a9498");
            when 18441653 => data <= (x"7895467276b7b907", x"8e545d92fd06e4fb", x"6944c4dce6f952ab", x"bbca10cc79c2c61b", x"f9abb4beb1258bfe", x"708ee7e2a520ac8e", x"7500579b0c51a527", x"2030eae8270158a1");
            when 17915659 => data <= (x"bca62edeac993963", x"c854185bb35d43c0", x"5efcc8a116213bfe", x"d5e746e36056eca9", x"c40e14b592dfc248", x"1b963659022d678f", x"f0ae53fbab871912", x"a21aa03fb72de91b");
            when 16584959 => data <= (x"a3c770a74b789cc2", x"e107369602f196f6", x"35429824f840a5b9", x"bd41249ccfe97654", x"da3d64ee958603ac", x"30ebde7a3499f157", x"5df6987a2dd7e01d", x"b7eeec095ea7c894");
            when 31432486 => data <= (x"e75d2b678b5d39be", x"4ac80f9780616390", x"0c7544b5e8ae3bcc", x"477df48b189befdb", x"5d9a3d81eba19706", x"1307b0ef00afd3f1", x"6bd23ff72ac523a4", x"bd37e06a427fd7b6");
            when 26614750 => data <= (x"2725757e2a4e7b0f", x"d9490a8a2be463e9", x"f722ad3290702262", x"a958c06a41694216", x"d8a1edb9e58b3a40", x"39f353b7f4a4e969", x"0b91c79df6039f40", x"87c475445618af98");
            when 17874132 => data <= (x"6e3e2b8ff1998973", x"7a6b06a2eb2a51ff", x"775f3bf87466d7ed", x"bac9f73b4532fc18", x"a934b17c2da57ab9", x"e42e72c81b952c89", x"165dbd47bd54061d", x"8f5b700ed2827cd3");
            when 27472908 => data <= (x"7b380e2963e7bc57", x"d1d090f8477635b8", x"3bd352bc10bd67dd", x"44491ccdc2180e72", x"bb08aeceaaa7cb0b", x"a01b152511f1e8b5", x"0d7d2e33d788b308", x"aeefacb52e6ba6a2");
            when 16600340 => data <= (x"b2a7ac8db7397c62", x"72e38f80cc7e6c71", x"243a50e94358a662", x"4465096daa0057e7", x"e2660d3b3775a915", x"09023af82b759f67", x"d5e3ea30e4cf33e8", x"07c03fd4179b9724");
            when 7533966 => data <= (x"7e96619eb135a1e4", x"0661f2f458dadd27", x"13dcf9b450193ade", x"18dc064a5194cad8", x"062d08b708013c93", x"03577136c073b67f", x"86f28476303c188c", x"580e7c5b14e8d0a2");
            when 10789213 => data <= (x"a8d1f077ce76469b", x"22f56090afd8ef6a", x"3baaec92d796b107", x"70e2ab6c1bffd4d9", x"7ec9770a88a4bb6a", x"7d01611b46f9a595", x"64fd48988b74907c", x"0dcffa7042298713");
            when 1141073 => data <= (x"2cfb100d9eb81612", x"219825e9168b7779", x"e18ae65f12f0d471", x"2915c609de727d09", x"a65f2e263438c40e", x"18e5c62aeca18ee9", x"a28a1e273a442dc8", x"52d777454ac37768");
            when 28801101 => data <= (x"feba9770ef6680a8", x"46e47ed0944d7e9b", x"1e32e21e2bfb92cf", x"e92d2bd9012e3c82", x"5bea725cf1392c3b", x"c2dab1a935a6a760", x"da4be5144c657911", x"dbcc89771be4f47e");
            when 31009537 => data <= (x"aa532b1f40de481e", x"fed14f1d6b0b9e1e", x"73385563b73110ac", x"6a51e78d45209926", x"4a500ab59ecb8ce4", x"357a7baf0520cfc4", x"1f0a4218788644bb", x"34eec4b8e0c673ef");
            when 25798743 => data <= (x"60d6e3fea9e07299", x"9d7664dd774918cc", x"f38c0ce81404191e", x"80b11126f1197cde", x"af063cb64d0cd692", x"8a7c1c25651e07e4", x"f9ffbbf73442530e", x"8459816c48c166b6");
            when 29519872 => data <= (x"17fee036c120d72c", x"dd5d6390b748c05e", x"68bbaa05279eaff6", x"12f500e219a34440", x"e609f3e100f1fdac", x"abfbea9b7a609557", x"dc2fa9ea225d2dc7", x"854deded2a894983");
            when 2108706 => data <= (x"0db0d77ada00bac2", x"0d59ddadff040d82", x"fb69932bd4da8c28", x"e3969e79e94aedab", x"67d63bf4f7f88d18", x"360297f3a4c40bb4", x"5cdbfe208b31f224", x"6bc9b056cb155767");
            when 18489013 => data <= (x"65f727ca55079187", x"4d38a2343773a526", x"7c7c792d8711df97", x"2119202b1ac3ff5e", x"e26806b627f58af4", x"a79a290943b7185e", x"f4fd4df011462de5", x"c6346e42aaee2554");
            when 5630209 => data <= (x"7c3529a1e5ec8c33", x"35d8813cad864a08", x"219c6a65c2ef1b86", x"c51e8b609d3190d4", x"90b0cb057f9d7df5", x"f2b7bb2b7ab43757", x"74921ff9f3d7d10c", x"04bfd4e6f336a071");
            when 11746742 => data <= (x"5284cb4673c70baf", x"14e6e98b07034fa6", x"bf603d1a5958d589", x"7c684fed4b0c3d86", x"fed2e281dfb5a2c3", x"b1b6eaa2153b92ef", x"2e763dc4c8b607ae", x"e1a4d1a7f13080f7");
            when 7563345 => data <= (x"fe291cc3791072d2", x"b16e9679afa2ee8e", x"d259160511ba1968", x"581576ceb8c23cd6", x"f616c301caa6d703", x"4b90785bc1ec7f83", x"b54f8bf893eb92eb", x"a02d3ba4b5a6b06b");
            when 27584916 => data <= (x"a55c3dbd2f6e3715", x"441b7ff6b84d619c", x"02f2bcb948ed7be0", x"dbdbbfd51379f51f", x"9c2f5acc4cfe3e15", x"e6b70bfaa7c503d6", x"7ca35edc87a14fbd", x"857913f2671797d2");
            when 16492751 => data <= (x"07b7f08cc39e705b", x"bbf46ee301d7a999", x"37411755976c9f96", x"732368814882b31a", x"9b9d22a898927acf", x"7223a9b45d640848", x"ea8b85d664b95635", x"1465cd6b549059c9");
            when 28944288 => data <= (x"ddfd7f2bbf3f108f", x"e41914e74c8b8834", x"a23701c6d1fd3752", x"4b55a06509d675f3", x"cddd6f805da7d9e2", x"9a3e48519cbe22e0", x"1f7bd3bd99b1f185", x"5668ff5d8e61da57");
            when 6399023 => data <= (x"a12fbf972aa1ac88", x"a80ef71298a08ed1", x"d914c6d4f0b1eb71", x"d127c8720ec19e37", x"0ca7f2b3abdf2b9f", x"07aaba7788450fda", x"5cd7f00cc15ae1e4", x"64ed358f5023dde4");
            when 22581512 => data <= (x"2b2b574b2fd33032", x"921b72a2531037f3", x"c3d6a3514c876db3", x"53ae95ba816439c1", x"345ff0c60350b8de", x"a2389246fcfd3292", x"87f556badb724844", x"f93a341046e1a046");
            when 7062964 => data <= (x"5bee600779eed2a5", x"354acb3bc3cacbc9", x"dac6b2b890e2c960", x"9c0c83a52f2a2ff3", x"ba62826e19f86ccb", x"a09451c3549e0846", x"e1672ed434b40a09", x"6ff9cbf31fb31fb8");
            when 31465810 => data <= (x"6f6752f02d2a7376", x"b8a989b42bb6fdc3", x"bfd725879c4d7d12", x"f635aafcfeffa660", x"090bef03523b911e", x"078adf8785f77589", x"75067c64e1306c1c", x"712dae396d6f2919");
            when 13128246 => data <= (x"8b9e959f87ac7d69", x"0580911d2e5771bb", x"b5238e4c94fcc635", x"eaa3dde9071d8877", x"b12edc6f5408991e", x"929dc860e81d0f91", x"2c5a3a50ab2fd887", x"5c54807f7163987b");
            when 12345117 => data <= (x"1689c4299d26d0f5", x"e45d957153223185", x"80cd4ad4257cf6b8", x"d7525e580de411f2", x"faadf4a380ed3738", x"b3a1dc905d8de623", x"467b45d00d4ea72a", x"11cfe07780ebac4d");
            when 4817190 => data <= (x"55e6cdae691b82cc", x"33bfefa2de595ef7", x"2f21c19520656cff", x"4011189cbb40dc5b", x"7d28026070dfc86f", x"c04e44d5f452f1c5", x"2ddfb7a451595211", x"a39c8c89d11cb4c8");
            when 30542560 => data <= (x"0777935336d75c9d", x"e4e6fc12b49b7d27", x"c56779557bbdf955", x"e75095b0079e911a", x"6a454aaedbddec95", x"37cc763017d96a09", x"d9aa318f7b9e8020", x"5894b5fb31442951");
            when 5452336 => data <= (x"1b6a16e3274a4d56", x"125c14004ecf0344", x"b189d36806c5391a", x"45dda9da9337e75c", x"36afb1252c1971d0", x"de2d26d15a450ca5", x"d009ad448da037dd", x"a82620c436e90e70");
            when 31660112 => data <= (x"f4d7a805de1418e0", x"5c3f6b7f4671eb4c", x"6d5809a8d3dbb78b", x"8b32c6c71f0f9cc8", x"a566aeac2e93b741", x"bebbfcd9fab82938", x"c9c65f78cc2967b2", x"112bf35dd3a49657");
            when 7917953 => data <= (x"0ca9bc17134e62a7", x"ac4220ac3f59012c", x"31f2da146cedd032", x"351b939ba35141be", x"70790ea1373caf65", x"014d28950087c0be", x"ea80078c3ef8814a", x"e26693cca785b39c");
            when 15784565 => data <= (x"f8bc110e0fa00d21", x"d585ad1939c133bd", x"042120da1289190b", x"63c489a7bba72319", x"fbc92afd0aece202", x"ba103df139870e9d", x"31c0f63ec29571fc", x"6e152f7929c80990");
            when 4680584 => data <= (x"440f7384b4a3597f", x"336685a0e8abcfbc", x"024a6c9a3c87237b", x"8afe956f5f1f4292", x"ee477870512bea76", x"529f6e649feec8d9", x"b5f4f5e9bae6bc84", x"3745596377cd2e5a");
            when 5948039 => data <= (x"800c0a1cac7b7584", x"607d88f825de6887", x"769b425699d98fed", x"1a398529a37e5726", x"aebed22136b6231b", x"0143853c011c9cbb", x"cd4aa23c4a51fd59", x"569debfc77981adc");
            when 4721315 => data <= (x"a1613371748ce1f0", x"fe09395afadd91b9", x"6f428f8d60d131d5", x"f4d8a5731539c717", x"b8166b88961103ca", x"71866939ed32a5c6", x"e4ce1a79b096fdf8", x"0806b4be4b38faa3");
            when 615748 => data <= (x"18dc929aeca7ce2c", x"f917045eed3cff86", x"9b39c9f5efdc3bc8", x"42ca05fdfb4ffe1b", x"ea52385d303f02d2", x"c4e0f0179dcf7d79", x"53dafa342b694d40", x"1a9d67478aed3ee6");
            when 13293083 => data <= (x"38576c4c567636da", x"2df1c66b25810c92", x"0c0476148cc4b132", x"1029bbc338688ae4", x"279ea94c8b3f4b2a", x"8efba262ab0ca292", x"b687019cf5492e93", x"699633e63486170f");
            when 32328992 => data <= (x"77579830df831bbe", x"4dbfc9ba89450441", x"431b64502cec867a", x"0b99e496076e8f39", x"81fb7ea33de34832", x"a3c9c65f0c6dce83", x"80166f16420fe217", x"9b0562c7271b4b36");
            when 32887744 => data <= (x"4a9ffd9d8ab370e1", x"2e6944f6253212f8", x"26f81bc03d5d16ba", x"402f8d62e32e5125", x"ffe044fcd26a447a", x"3d3a4abb3de09761", x"eaaf8d9b83b980fe", x"655b28a7b2d284a6");
            when 8545299 => data <= (x"5dc462bf43d8ffd0", x"8cec89fcac20a64d", x"7e81f0c888175e7d", x"411e30cc8004950a", x"7ee6c855bfb33ec6", x"9b17d3307d33865b", x"da45e46b71255a01", x"06e088f032296f55");
            when 24300163 => data <= (x"1ac9657aa0968bbd", x"af7d4c1849b261f5", x"27ae859343a348ab", x"7c1450b9cf748cb0", x"38c3f57823d28203", x"bc16590109cbac29", x"647ec69a90b9b792", x"731f25ef612d7a7d");
            when 13282167 => data <= (x"e55a34da0faaf347", x"ce16f70fa95ed7c4", x"46559e7060767648", x"8e198b4b2bf8c512", x"e06a2db39beceef9", x"9707e6328e9ee107", x"95c535a3d6beeb09", x"029bf490c199beef");
            when 20799720 => data <= (x"6fb7df566551b6a8", x"f7eecbb47c94724e", x"d290f13d5f5e5c8a", x"f5382302a846bb47", x"39cb171d991ddaef", x"fe86c91307bd49cf", x"a44c28ed956dcb72", x"0fb7a29a80dd37bc");
            when 19196595 => data <= (x"16268a61bcee7436", x"1269f4a8e984aa6e", x"596b2cc154a5c163", x"54ad11723c09ff49", x"f88bcf5628e67e01", x"c62a61b7b334894a", x"149205cba92aa163", x"45223e2998ec237a");
            when 5078603 => data <= (x"de58ca0a66c86808", x"5dc3860bcec0e3e6", x"fd8fcfaa5a6d3ae5", x"27c8a5e5040ace54", x"4870f8375dd95090", x"65fd471b01882fb6", x"4b92be26c766204a", x"6702f2fde2e07baa");
            when 1164133 => data <= (x"a828c487a2dc9e3e", x"128b5eeb85c25d58", x"4fe33653e8d1fca2", x"1c7d7800a93cab07", x"a45c9d55a7cc5bd3", x"60ee3126ea37f4ab", x"84050141661dd559", x"7505d1e1ebf52348");
            when 28820521 => data <= (x"20a5205a5ebbfa48", x"c4b8838e0975823e", x"36746090f5d4d033", x"19c4abc8267a3722", x"79c811bceb374add", x"8266d55e9e3e591b", x"f851c88866a261bd", x"5916d85407c486d2");
            when 858783 => data <= (x"58f663b8a576bd97", x"cc85253be72a3524", x"2bad86cf332f66fa", x"51505fbc615482e7", x"a6180458724d9e87", x"34133b606775b914", x"b21f39f28022937b", x"e76484a4e66c7af2");
            when 32200204 => data <= (x"ef307cbeebd51024", x"ca73144e2f2ff5b0", x"239342ec50e20541", x"6b4dac53c2850fcb", x"a0c7e76388668292", x"b2837f7d3e7ac86e", x"a5c47c1661a39e3e", x"8e5ef656782c9d26");
            when 6321849 => data <= (x"0bc0df8ccaf6c750", x"d3bd5092f3431b18", x"5fda908647448b1b", x"3d90e413f493cdc2", x"78512a011b10d44c", x"5dbb0216242708eb", x"d705b1a335892bf2", x"35cec07d16029821");
            when 6975706 => data <= (x"67dea55ff95bdfc3", x"cd2405318682c4c9", x"5fa8ac2a56495395", x"4ae841f8d36789da", x"70cd60674fe71978", x"4da821f94c9e42e2", x"36ec8cffdf4e2a07", x"eaa94268da50ea5b");
            when 30264416 => data <= (x"954a46973d943c96", x"458193e330a9417d", x"befd8d1a4c86e02c", x"db61fdb0f8c6197f", x"02c7322a191165f8", x"6812b842686a43af", x"2836fe28d613daee", x"0e253a2924d1fc0c");
            when 5335469 => data <= (x"4649c3c993ab3dcd", x"28dc23b8244b684d", x"692297052d91302f", x"8f0585c864211300", x"bc8d1d725bf895f9", x"c41309688866458e", x"3b0604ed286b030a", x"f93b78bba592f677");
            when 22284126 => data <= (x"7100acd5ac9b98df", x"0a7eeecb2634504b", x"4c16abf6e81eaa49", x"e2e4c8ba92a10ff8", x"b65047b95b9b66bb", x"8c0f457af040ca0c", x"22c0df23810c3df3", x"0a13eb68d68c6f92");
            when 5919340 => data <= (x"32a6737ac6a730a1", x"fab1c9284c2f0da3", x"ccbebf9a0a0f84a9", x"f6501429cb80db23", x"c4de9f6686768196", x"be0555df7a9aeb5b", x"0be2869ff4b0f6ca", x"146efa3833cd4d61");
            when 7704633 => data <= (x"887f3fb5214ba993", x"abfebe9360d3903a", x"b85324e438bc102c", x"c2b8d5258a93a89d", x"9e023964f4351bb1", x"9e76d3dce05529b5", x"325295ed124893b8", x"3b05d387cb996778");
            when 27519803 => data <= (x"c3e47b4c1f413548", x"e205c4fcb08e699e", x"821476ba9b81e36b", x"aca3695784af77e0", x"6edb3c580ec94675", x"35e877a363319bfd", x"53d471ee5789609a", x"ba29fe0485837139");
            when 8851680 => data <= (x"0b865ab1b1ccdf50", x"c2f66916f973647e", x"b073fc9001f1efd0", x"e503be57a4407d1f", x"446c9617917e29c3", x"9d9f1e8c77acc6a0", x"eb6dbdd74fcefd59", x"5b2f2e6b0e71f46b");
            when 11117854 => data <= (x"cc67135ab5e5b149", x"0f513a28cd3247e4", x"dfafb1caa9b3f819", x"59d1a0214d251d0f", x"788fa18c840edd04", x"ed013563a952f30e", x"bb3194107189fa3d", x"9129245267fb63fe");
            when 3454488 => data <= (x"64a6cd6bc785be49", x"c22ad2f4412290fc", x"9bc765fa36887903", x"93a44a9fccd27e3a", x"1ee580f0b5220932", x"08be09b0e950d2f5", x"50fdccd7bcaf3ea8", x"3385158a6bbafa4b");
            when 2224969 => data <= (x"70bd30f814d6c8fd", x"88eef8ecf28e7fa8", x"b785d531b0046540", x"ad1514a6d9aafb59", x"3859e365b337af01", x"a8d470eaab501aba", x"ed1842a0d3980100", x"a53fb241f622b56a");
            when 24413521 => data <= (x"6fb274b960bf6e55", x"9cd33d428b7a3e18", x"ce763b930b26b940", x"0dd428002f0dc360", x"9988dc4dc68e382a", x"2ffbe754228def74", x"cfeab41211522a42", x"05137bdf6c57f28f");
            when 1837141 => data <= (x"e41a5cf6f5db9189", x"f6caecb0753ed76b", x"b6ec0163809f2be9", x"28da7503ffc762ca", x"69f090ac85b0350d", x"14d96860412bc790", x"4df429257a3a95c9", x"4541e6a7d98a27ac");
            when 14127159 => data <= (x"e1f8f321ee8612d9", x"68bd219d8e3e717e", x"8953887a5c87ffbd", x"770cbc669c7057d9", x"7c3409de2de2ddc1", x"3099e887ff037650", x"d626ccb3ff63d7af", x"55651572c8d2af50");
            when 14902036 => data <= (x"a71e17b2c6a511ab", x"34d475a79d731760", x"527d377a2084fe4e", x"377b62aefc5cc7c9", x"7747ad660633c61e", x"17a8a31280f7ac5f", x"af4445dd79770362", x"3fcaaf6d25c89dac");
            when 8558509 => data <= (x"cb49f4244acd3666", x"7ac9e8e58427d5a0", x"3dc94a6294bf6348", x"efa52904a7f77531", x"b35da6e82fae507e", x"e65abdd8859d10ea", x"b3a09b14419cad24", x"49db74ee6249f76f");
            when 22670833 => data <= (x"58e11318dba6b031", x"d45af22620719d8b", x"9fe7292b83a290f3", x"66f4c3d6fc5f0a6f", x"e1008d8a4545e0f5", x"126f5d2f3d3cea71", x"baa3bb5c0dbdff27", x"7868f206e5547673");
            when 11325444 => data <= (x"493d48175a95fc40", x"8cdf78035f4f93ce", x"15f39559abc0591c", x"73d6d41fcfe999ab", x"b00694ed4f2980f9", x"717e459ff9211cc9", x"0ed45ddf692afca6", x"1da41f13656f45ac");
            when 20047496 => data <= (x"27fa953050075aba", x"f22b140f9b0f0a3f", x"5394102f9c75c912", x"77af24475f7bd866", x"ea8b96444475dcfb", x"15a930f9567b4a0e", x"ee9b3bc22461828a", x"e88ed7865864d68e");
            when 1816545 => data <= (x"bec97c465b4909d2", x"5d1f7b5d19df6c87", x"e80fc2fa40792728", x"5266e8b57a833d0f", x"7e81c45ac88409ec", x"120a43d4ab655e28", x"fdfc07ec869df5d9", x"31bd2bf6d3925fe1");
            when 31647922 => data <= (x"20e93ead373213be", x"85861ffc3ac52890", x"8721486314fb2cbd", x"a49aace1cf627138", x"0ca88371fad3e463", x"51fdb7aecf7d81f6", x"d69b033b11d00b8e", x"6bdd1034dbf219b6");
            when 22251480 => data <= (x"37af55ada080baa6", x"d68c5b59af1f7149", x"71637f1ae2815980", x"d8183522e7db0dfc", x"f2f2adfa65650859", x"de3f74cf277c7c95", x"94de66a6ed7a0078", x"4d064512dbd1b7e3");
            when 6635937 => data <= (x"374e65c6fa122ea1", x"1a9347c6b967d1e2", x"67da59de4fce3280", x"e069b2cd51e1a031", x"8476ef4fa26761fa", x"44030fbe8ff1bd56", x"9ebe9da94fde0cf8", x"bfa6e13256866c5b");
            when 24817704 => data <= (x"6c644192ec82dc1d", x"7a6854f47c8a2db7", x"7de378fb603e98d6", x"74d20c66d16d9490", x"78adab99ea16328a", x"94940281bfb633b1", x"cc582a538d3d6a0f", x"3b75d25d5dbd89a0");
            when 16888012 => data <= (x"2903d9c1af8da3d2", x"4cbd1fe4ff47d934", x"a236f15db576596c", x"3cc8f759a046a94d", x"a60137bcbeaee10a", x"4f9d2f489d9d5a52", x"59c0c54ad0e7252e", x"72417141d4a3bec5");
            when 14967559 => data <= (x"76dcc6caf5ab156f", x"02ebdc07e5d82db4", x"8bdb9f62611f33d4", x"a201a91151c26852", x"3dd51ac40de0fb34", x"ed45f8a918838599", x"d6c15cf19f749452", x"f6bb6d6eed7b2116");
            when 22011943 => data <= (x"ae0ef04b2c8ecc05", x"7638d4a26d08a412", x"63c18a59ddd5e3c9", x"cd3f3e771a0e24e3", x"4f61f188631c3c77", x"d8b893ef87e2679a", x"a5579d5caf9c936d", x"4c38da08071d7484");
            when 6644164 => data <= (x"946a34ae21c1d34f", x"7d15cf56d3ed4cd8", x"813f13874d008114", x"78eea14e0ff544e8", x"6598d9bf1a1b0b0f", x"835c3cd7b51df043", x"71483199f7381c27", x"5061d1b40f831271");
            when 1845592 => data <= (x"bfa142ca96c8ea4a", x"659e73e31a5c33bf", x"7b456bdbef5a6116", x"129b4da335b85592", x"f41bf50ca861bd91", x"aac9ee07ab05afa2", x"57f5f1dbda80b5a8", x"d8cc33f89c329915");
            when 9328546 => data <= (x"9019afa6a9a5cd87", x"05430be708b3867a", x"0d33a352c377c4c7", x"17126ad6c4d93056", x"88dff4d9923a939c", x"03f6ddd491bef5de", x"386c2ef51f661a27", x"98c7942cb4585ec2");
            when 11595190 => data <= (x"1328e6cd2b0c1d75", x"05deb614f7a603c2", x"c32c7fc9cb444a31", x"0c223fa6e6683cde", x"510edfc1c73dd0cb", x"d3d0d99e0a70ffd2", x"3b2b8b5d422fa987", x"0f9ab4ac6a53cd21");
            when 8382261 => data <= (x"707c00cd1d5413b1", x"93052c9fb80684a8", x"c43a5e962f9a1934", x"46e62d6d9c855d8a", x"899a38c2822dcbd9", x"eb0ece830ce6597b", x"efa3ebd04c5a0b0d", x"62064238ca6ab4c9");
            when 4702460 => data <= (x"04ca5c2c79ba8289", x"ca79378d29952564", x"e9ee7cc95a0b9bf5", x"f0c5679aa0adb896", x"9d134f39ffa25487", x"379f2b501e15e831", x"a7b5c13c3fdf250a", x"cb5af78ce9947573");
            when 31475382 => data <= (x"1bfdee88aff32762", x"362164e0c94ef0ec", x"e4dc48de0c733852", x"5f6d8e61992e8fee", x"78685b64128c6bb1", x"f0482064c7e0f0f4", x"ccd4906a929dda7a", x"b6101fd658aeeb14");
            when 18613755 => data <= (x"86d0f290c05bf9f5", x"e641f69a2e63918b", x"ad8d2e8ab5af4d4b", x"fee4669fc9495331", x"1c3aaf355a8e5df0", x"3f96e43156a79d2f", x"9aaf9a25ea703d2c", x"7ade0ae166a14b7a");
            when 15854133 => data <= (x"fe45b31d6acf1c91", x"23bedf22086d1cdb", x"a6c166bd02b21fa6", x"a880316428bff999", x"89acbb525916a0b5", x"b0041e919c9a580f", x"304cbbaa4c769bd9", x"6ce3440d8844e514");
            when 5962004 => data <= (x"7c3d6ef90519dfe2", x"1cd56549480a8d14", x"f81ee539e64a615b", x"3309a87d944140c0", x"9d9916df132363d3", x"f2753deb64bf6eb5", x"185b1de8e7adf990", x"55c06570be30de07");
            when 4236909 => data <= (x"873eae5e19a6249c", x"e80e69b1eb15b5d2", x"a2985be1c93e6bce", x"d408ec76a27722bc", x"50fb4234c6048969", x"b054e91186f649c5", x"c01a5ea28d6d0fdb", x"20623a55ffa73801");
            when 21244829 => data <= (x"af2c3109204b5d2b", x"4cde4fc05bbacc80", x"170b3c6716ce6050", x"aa37144c9c6f026d", x"877483dc4739ebeb", x"9f7dcc9b0d343e96", x"ebf0e993e4839ff8", x"f08f78f3f4435135");
            when 9330940 => data <= (x"d29d0f79b4666060", x"d9522ed75799c8a2", x"e347e6af5f9bb9ec", x"46eeaf0d976c8888", x"be1290d2b3f779d2", x"52bf48dc9a1e3255", x"b977984ca6bbd0f2", x"c0ef484e99962ab9");
            when 19068335 => data <= (x"3953182acf5561b2", x"6b8c136a3a88d51a", x"1891a22a30b8319a", x"f4d208ebd2894bf6", x"db458b1a6be87f3c", x"6fc016d82bd6c048", x"10dd6e2e440b2bcc", x"f8f8a9c102b0a526");
            when 14500240 => data <= (x"71a874722e53c6f7", x"76884d9809b927d8", x"2dd1b7fa5c1941be", x"f5e75de9b5758043", x"d730117ddbabfe1d", x"6019a17079400de1", x"98f38017d1b56e27", x"43b94d529cdf7331");
            when 17172476 => data <= (x"e63f200356744867", x"c6b19dc101aa1d96", x"052ab2bd67b4fee2", x"68d7f60c76621fc9", x"487a61e467c9202f", x"b932fac4f41cfe6f", x"fe61c53af652278c", x"6a8a1f6d96074c4e");
            when 16663757 => data <= (x"2ae4d4822cb16fd7", x"6442d0a9f79f8a2e", x"1666696192215e15", x"310db55d97ae6bff", x"9e5ca83de72f94b6", x"c471677214b56320", x"63706e9b937d2a8c", x"684672487b98b485");
            when 27872029 => data <= (x"ac7bb53a5ca0aba9", x"4043c311a0ea9d1c", x"04dcd306650ae4c2", x"abf7a90194fd3e18", x"a9149a60462a3ec5", x"e0ebc9c8fb79dfe8", x"1a920a935809f233", x"55949de66c728fb4");
            when 24763560 => data <= (x"c57ccaebccb19787", x"23f49feb50f1a32a", x"e71fdd1574eac796", x"c58708f606d07597", x"9414f64b67c686c1", x"e42829acd6cc02f4", x"17f5551341fdf54b", x"c85185762d0cd714");
            when 32121028 => data <= (x"09a4a8430d1abf34", x"dfcdb6ca24a3079d", x"737ab06ee1d8e88c", x"4c003429ec45b34f", x"d6186370a3d2b5c3", x"d4c49f341905529b", x"8ad725a94d526819", x"9b77e065f8c4ba16");
            when 23086653 => data <= (x"5ef7caa83c14ce64", x"ff5c883c272e6706", x"0557e2949d6014f0", x"b7360055d0b07393", x"9de31a599f8b1772", x"45b45482c5ac0347", x"6438c84897fea940", x"33ce0d49694ec6e2");
            when 23527647 => data <= (x"32c3dd317067edca", x"3b3809b8fa5b60e0", x"367d234c215c33e3", x"e0aa2fedaa3fac1e", x"22a254d401b47625", x"49a4a0a49d7b4b17", x"6469cddf922e1468", x"98f8016ee5e0485d");
            when 29426195 => data <= (x"80f5f61fd366003e", x"2ccbd460135fe3e4", x"0891bafda682ba03", x"a8f328ee12294032", x"ef47b086f5df49f9", x"8296c3285a7753de", x"2abbb9fd9c114323", x"f3461b3065f6d578");
            when 19004771 => data <= (x"f0c20997f994f1f8", x"ffd0cfb261e3eff5", x"f43b15dbf381c971", x"8635f4afa4cf9872", x"f02e6c81ba36ace8", x"ef060b4c43068847", x"19022a7d0a36f516", x"7084b368f8daa6cf");
            when 13938474 => data <= (x"ef1fea1e8ed58b5e", x"90609315702efa5a", x"bcc212548c9f96e7", x"1095eca1d90bd187", x"90e1af07942d3b6d", x"36fdebc168d5dd4c", x"66e0de3ca153b9da", x"5bf53aa5e228a639");
            when 5689812 => data <= (x"3798b3cdb24c8926", x"445dc67158a6d62c", x"5f526cc055a7deb7", x"0ef670a1dcd8eae9", x"ae9993edce1b9862", x"31c926d3136aceb9", x"445d152994b34a34", x"d4f2b516d97809f3");
            when 6042610 => data <= (x"658e69c7ea050bff", x"4520ff5b5c2006c7", x"c7fabaf8e6fa32f4", x"604c3f5347461f53", x"294cf20eb111c260", x"ae283c8734be6543", x"d7473193435bcc30", x"c31f0186e8dbf038");
            when 16573421 => data <= (x"1b4cd146354ee559", x"df6020a8ae0bd5ff", x"627adeaecc18dd78", x"0fa2469f5d9f6b02", x"66bf6727737754ad", x"197f5c8029267079", x"5337133fa2a5595f", x"56bfe120200b0b8a");
            when 28408553 => data <= (x"02864cd0d5df421f", x"9a91663f681d06ad", x"50a69034dda7d0e2", x"083d702e3ba4d987", x"4a68a21c77fa8d0f", x"4f0d48232cc4898b", x"d4ecc56daf25e893", x"aa2bbcbc09bb5d91");
            when 5595781 => data <= (x"0a863067d052698a", x"70df0cb5c6acaa27", x"5c6aa2e7e019fe10", x"93e57bdaa817e068", x"6c3ee855ac5544ef", x"a31b248d7a2785a0", x"4d065f1992b949b2", x"fa44d3c6fa216b78");
            when 8075416 => data <= (x"7fcade1041800dfd", x"1b1533a3eb58a61c", x"9e6d5ba3789d2344", x"ecb96abb54db9037", x"0aac2a2a325d5005", x"4795f3ad6ba4e16e", x"530ccb1e1616b529", x"4b3a68f81bae145f");
            when 26706150 => data <= (x"d09fc65750dae8c3", x"95f2f11a1b994697", x"d6df8c10eb4f0775", x"4308f27f29542a63", x"467be19528ffcc08", x"d01dfb09e2bdfe18", x"bfaa67eaf07bc3ae", x"e581ad67fb2aa7d5");
            when 9635755 => data <= (x"a6f65bfac778bc1c", x"0259790711824d37", x"a0d333069fa1f66b", x"e973eedded51f6b5", x"4cad9c13c254b08d", x"e2b2c25bedb0ae99", x"21eb0127d790e96e", x"e8e5a2acf06c4e13");
            when 26333364 => data <= (x"b2840cc8d1a3c11e", x"9431333493345f4a", x"0e5b9e94208b1855", x"75b19ce90bd8f952", x"b1d9dcae2396581d", x"35f1d9f99b0b16a9", x"6bab323bdad2f8db", x"eb613b7e30690c36");
            when 16566768 => data <= (x"e446b52d3f1fe5fe", x"d600bb25fdbd9806", x"f6285e952a8864df", x"c33a9a14ef7c4e8c", x"3d091ab0e0d2c381", x"ea1d40dd03bc0868", x"f6ff81cd2e0c453b", x"814d4cecd9f31a7f");
            when 16039942 => data <= (x"78c34cc34dff4cec", x"e7b483bb6fa9fe4b", x"62f01be6b9f2bef7", x"12dc21ad660535a4", x"f5d32462d4b879f8", x"deb4c7eaa6523e3c", x"d6a2d025cdeb6fb9", x"a698a5c20cb39acc");
            when 13191384 => data <= (x"39c61ce1dd219b86", x"49575581645d254f", x"a4bc446b24580478", x"7e62d8a10e89ba66", x"1fd6d2639716fdae", x"6ca61ffeccc6503c", x"58315470038a0929", x"bc759aeb59563064");
            when 25380263 => data <= (x"2ecfeccdca14a77f", x"96c50ccaced2b788", x"19601a066353c8d5", x"cd343a458ed018d4", x"e233933ead00745f", x"3bb4751e43d7eedb", x"1db7d7613c1e5d6e", x"06e4144c4097d278");
            when 11635011 => data <= (x"193444ac1968b89a", x"005592713acf7a91", x"2329a2c0443e901d", x"5d34aaeed67cfe89", x"fb72236e97ad180b", x"48bcfb2b43237eac", x"4d7798f311936122", x"ecf0fe73322e7c81");
            when 27210827 => data <= (x"4ad424f61b9b9fe9", x"4d5693a9d0fb51b4", x"a3c0a51389c5f967", x"a9efcbc15058918d", x"c9f592bd705702bb", x"08317545b52b50dc", x"4b2f1c618b725aa8", x"cc5b226b0c89e3a2");
            when 1753954 => data <= (x"eaafcf55856feaf8", x"10010a4426c152e5", x"6f687b1a85527802", x"447347138a8b6b0b", x"3776609a8f606d29", x"bb3862c3a5d0a9c0", x"292b1f8adc974493", x"3462911d8cfc87f8");
            when 22195930 => data <= (x"a06e843f5edb7331", x"1504f12f2355d045", x"d18d48ba2c4ad785", x"0a5f262601246a8a", x"b41279b6f083562c", x"a14fa01910110dc7", x"bba08bbfbaa6ac6e", x"3427b931667569a3");
            when 7908290 => data <= (x"b43e53de6241e590", x"7e3a3c8c30fa6cc2", x"8e16faaac19ba8b4", x"47895bd170dc8eae", x"c445ece19c111d86", x"e6a39d3a9d0aed63", x"37b6e6fbb66ca56b", x"3b608e0a3e263e07");
            when 18633970 => data <= (x"76db817a07fb4479", x"04807a11b90f1cee", x"3af9e7c27cecb3aa", x"e57169717cdd2df2", x"eac88e6a88d60e1d", x"1b60bf9f74005a34", x"f6fee77c0c54ac35", x"b5bfff10a857e8d5");
            when 25354870 => data <= (x"aca0bb698b490629", x"eff92e1083525e3c", x"48219b5feeb8a980", x"0351f46d4dacec97", x"6cd4f2be1fdf9890", x"04bd66e2310b7390", x"2da1c5e8f86348f7", x"75e7358231a0e987");
            when 33032658 => data <= (x"cff17ec8c5c702c7", x"27032d996cb35988", x"4127659fd8081435", x"0f406df3b193b74f", x"7a5f44a015aebdd3", x"985ce1b5a2986dea", x"bf04d45d927d5f37", x"673c395765162f20");
            when 22250751 => data <= (x"4196cfbad1501c97", x"d229b85093a20a0d", x"e131eaf973e61046", x"d626c6c7b6e2e688", x"8b3e46931e2488bb", x"64cec8ad0dd8994d", x"da68e02cfaf0e567", x"eb2009767aafb2e1");
            when 11478895 => data <= (x"75d254ae291db485", x"d682c0281c9dd07a", x"bc9c333d3deaa5c9", x"42e5ca60351d6807", x"9935e1079d5001b1", x"e606587b15c78b4c", x"7964f7521448d44c", x"b7dc7911bfff3638");
            when 12376094 => data <= (x"6406ce3c71afae80", x"bb9ec7eacb6dac16", x"1dff68f71f29d94b", x"c20fb63c6576d78e", x"e18dbf9638e2a186", x"98f5ff137ec6ed6e", x"9a58bca369f0014e", x"7459fec0113b33f3");
            when 11177502 => data <= (x"92bbcd6b349e69b0", x"9b22dd55905be608", x"12a0c157432e3658", x"a6c49764285284e4", x"1f6d50536b08b705", x"61e7771631f180fe", x"7b7daac438d6a834", x"ad7a0c334a8e6acc");
            when 19931161 => data <= (x"d1d6ae5b2c2f6754", x"26d76ad1125280bc", x"f0d1bba5d5e8dc64", x"f0d26af00cc2acba", x"b1982ce61e23ccb2", x"05d466329879e646", x"0da7e6207fb81d25", x"d7ca2c0c59cee22f");
            when 9483614 => data <= (x"b50b720ec819d744", x"b0bdebe74a0f5aa8", x"465c6774ab1b3053", x"dd04040fa457db17", x"75b375aacac622cf", x"74c8509214c182ca", x"70ff61e8f42db141", x"ae0b955984156a02");
            when 20404898 => data <= (x"c3779dfa23fb276e", x"90f356f77fd65ebf", x"55d48a084c84d62b", x"d46aea7a0ed3f234", x"1a5c93062848146e", x"3bbeec5779c27213", x"eeca1e840aacc63f", x"4a9609fcc8a88d8d");
            when 14525613 => data <= (x"e04914c3924b24c1", x"8e619b5a85d7a2c9", x"e61dc1c959894e3d", x"9ffead9101ee3713", x"9c315a5093e876e8", x"7661a1601ddb7b94", x"ceb873a34f9aa06e", x"6f3dd10207b4b340");
            when 28173180 => data <= (x"d6b51af9ec79a906", x"b224b7c263b1cf95", x"8472016a17269e70", x"855f072279ad27c7", x"8393760b41d9ae89", x"67c5282fcb4f32a6", x"ac54a54942cedf2b", x"0d70c1a37ee50ccd");
            when 16574210 => data <= (x"18cb70877872d84e", x"6359dd35d6174d28", x"bcf31b9c922a4e01", x"b159d175e0dca6f0", x"e6e7546c76fbb9fe", x"6d52f0a04e4ae763", x"ed925d8e62336911", x"168773f188f8e237");
            when 21267952 => data <= (x"6bd4a8958b6734ef", x"7ebb0a5e49db8a71", x"f33b9cc70d2e6d9c", x"f636f3768b77c89b", x"e2f9222f81a9b35c", x"0870efcf4c55e250", x"9516da8b1dc54464", x"2576ad675281ebb2");
            when 366321 => data <= (x"1d17839992a658cb", x"8ce15fb4aac10934", x"fa3d63b4836da4da", x"66c4296014276275", x"ab02434e4553a759", x"819937318de60d11", x"0c6e7e72cca6b98f", x"8a6be5b5f62e4dd8");
            when 25635317 => data <= (x"a67a4024e029f0a6", x"78ae444751a7f65c", x"73ac87ac45f234fe", x"eb1342773839fa4a", x"0c54a26c6b63380d", x"07b96d4d04547620", x"92d8b9f2a1abdc63", x"4097d0ed208f9266");
            when 18077162 => data <= (x"9cf08376853ea048", x"008eea2682aabb93", x"842eec33bce49031", x"5d2c0ae682f03a55", x"c5991e0bad21845e", x"5e334b52828a32ee", x"18dd29e8c5af5afb", x"d5b30cc4badc163e");
            when 11672656 => data <= (x"7c8e05d975878865", x"96a28b826ecca06d", x"30f977a155719264", x"b84d2189951f2760", x"dac39eea3739257e", x"410e7012145c5252", x"c28d24ae9ec6afb7", x"29057f84c3b607c6");
            when 15366372 => data <= (x"c5839f288891d1b9", x"28684bfb79463c35", x"6ee0c0288dc54390", x"1ccbda93d2770bc6", x"759efc68244e6cb5", x"6a91a0701f7256ef", x"e6dd7d7cf46ede40", x"c35f2b7aaee8e847");
            when 32559573 => data <= (x"b4b70fc78c184b5e", x"de4795a4a4f7c93e", x"f7c5ba305e4257e0", x"a99c02e1ad9d5891", x"230bed495efbba00", x"2c2968966a0c5dc0", x"04361e6f5b5a1c15", x"3ef19f15977bb994");
            when 17474779 => data <= (x"f2e090f4da3fbda0", x"a9bf2c57ee481ef8", x"70c785108f5df21e", x"791be18a82c878b3", x"f655312cc105a878", x"aebd5147ea9af8e2", x"ee948fa069e14356", x"8214f4f09a3bdaab");
            when 29272792 => data <= (x"0a64f64219b901f8", x"da07ce3ec7c85cea", x"59f8e08b9903ef5d", x"e43e6174a317d748", x"6a47803928f176a1", x"aea0957bd0504012", x"05510a5d51463946", x"79eeaa149c09b49e");
            when 27790251 => data <= (x"3d2b5ced21fb1246", x"6f192f6d6bf28c07", x"4b85dec7a9d4f455", x"33adef2bb709c52e", x"6e3e9667b33205e5", x"99ac064ca7846197", x"b3a175185cc386aa", x"70b94308fbab9c85");
            when 29149702 => data <= (x"90865e3a6e1ea2f1", x"9ff6cc2c034afe04", x"83e88168d5649c23", x"2eea066b92f9a2ef", x"892211e505eca9f1", x"b50676999e770874", x"526cd55767dc63be", x"8a56f033bafd5b1e");
            when 7712586 => data <= (x"6ebc72e8ce818a14", x"5764db5b2e41260f", x"d57498d2b8c8c12f", x"757de44b4f9ac58e", x"c55428e0d6c8f655", x"fdf92b1e5ad3761e", x"138edc07df7b50b6", x"de8f4b0db4345df2");
            when 8225082 => data <= (x"886a658bc0adc868", x"8705e8b0e5ac4fe1", x"4a7836e7a2c01e8a", x"b690a2aae193cb36", x"0132ccc9c71abc9f", x"111146bfa2892881", x"8b4cf0b24bbf3731", x"cf09196faf61ab65");
            when 29507734 => data <= (x"17322fae385fbc92", x"9b30afc1a3b8107e", x"487a6f1fb2b7b2f8", x"c4e3aa1352457e8c", x"bf8f03381b79b781", x"29ea4839477e6ec7", x"868565018e2d967e", x"a4adbced147f4cc3");
            when 7857432 => data <= (x"cde19e239a4dfcbf", x"9e44d3e76145709a", x"e1602aea9fee6ac5", x"844beb08561cbe34", x"e427327123302278", x"c44be64bc26378ef", x"0942da3001ab0274", x"3a572e976615cc6a");
            when 11504944 => data <= (x"49538b593f11ddfe", x"64af28aa9b53587c", x"ae125cc949a7c533", x"2e78e0825318162d", x"5f6ba717fae97d96", x"069e4e2e05ca72db", x"99ef5b593c20e0b1", x"3e28f312b3eb1561");
            when 4585853 => data <= (x"a8bc92f242a4619b", x"9f1eaded3e1d9888", x"8856fd842021e741", x"df0bd0185ebd510f", x"54c3b4a7a7ee07b3", x"35a258ed463d5177", x"bfa55934359105c9", x"9f8496f0b88f16a5");
            when 9974033 => data <= (x"c3714a2b913832b0", x"952790972c5c9adc", x"34245ee758789448", x"104716d9ad399dd2", x"ec582d3c0e781b35", x"1817693c8b8deeac", x"a326f87051966202", x"bcaee5c993bc4e69");
            when 1749718 => data <= (x"7fd9d6c87dd07edb", x"51311d84aecb1176", x"fe19262d369f4806", x"bc290846b922a05e", x"eb3078208eaa3fe3", x"251f32662cabc096", x"f9121e971e4e8e58", x"44d5d012acc016f6");
            when 12672347 => data <= (x"33d73f1eb787c08b", x"7fb6814e7ea13d18", x"02ed7dc066730467", x"34502963b520c0e3", x"5d6c73c4ca2f62fb", x"4a18af8d0ec66f0e", x"a7e03a45f4fc7d9a", x"aae5213dda4ba1e3");
            when 3655821 => data <= (x"9be70f7ce6d04fb9", x"e089155a2fabcbae", x"94ab444a3ec80b4d", x"6f1ae243896e8c84", x"6d36a49bdd53dcc8", x"a45b62cc307380ec", x"63673f30d06d5030", x"754f0124e42d29b6");
            when 23610479 => data <= (x"e2a614a78a09ae09", x"a460a2e7ab2432de", x"c76e98ff28667e17", x"f455b2f9b2668c27", x"8b23cd37a78d8f3f", x"99c9b9d88cf37fed", x"9540f57e5e572faa", x"089d7ab3443eb5aa");
            when 10348098 => data <= (x"527b4fd40ea6606c", x"3deb26284ed75931", x"dde9dbfc4cc8521f", x"36a34e76287966db", x"0bce820399a62e53", x"3cb1eeb4dcfdca56", x"3decaf3c875120c7", x"305f4e920a9015a6");
            when 22394988 => data <= (x"5eea9a9a915ef77c", x"eb394ee94146fb81", x"d41013555da7c747", x"ab4d5928d0652761", x"6c289fab32924ddc", x"033f7495547c8712", x"78eb2f8e7ae38ba2", x"4ac2747683f46ac0");
            when 19288285 => data <= (x"7ebd8df3b48e2733", x"687113419c632e44", x"f76e6ff7c8e841fc", x"b7411a91226e466a", x"f5a1f3f8cdb99c18", x"0f6dcd0f6855fa84", x"a0849919081b0f1b", x"59ee8b631f7ac624");
            when 29629939 => data <= (x"fb3e7573fabd430a", x"a7dd7638fd91072a", x"3604e7ca85e4f7bf", x"42bd789c9061b40a", x"c10ff53338420f36", x"611a7c441ae6d7c9", x"1b710ada90ca2785", x"4f314e154297baab");
            when 5471098 => data <= (x"e389558d9d78851e", x"ee91236fe3d6e2d6", x"3cc6263a0390c26f", x"52f44cdee39959ab", x"793ed6d3e43603e5", x"47efd5291b94b6c2", x"4c98448f5a5fa4fc", x"b4889dc4acafff18");
            when 31999425 => data <= (x"cda909a2fbb2c797", x"f5e4a576990c08cd", x"1ae5e52ab0f84a34", x"2b520fd0e220a4a7", x"b397127db1e284b5", x"8a973a919a3cc86b", x"44c8b2b61ee58517", x"74e4146bded97c6a");
            when 33100252 => data <= (x"16f1cd216deaee70", x"21e463c47264e5c3", x"5ea66f82b2185774", x"68cda64e32a8e0b5", x"db9f7b940001c932", x"c82899bea4648edf", x"3c90294a67fa9c98", x"4b4b1933fc3ffbea");
            when 31706515 => data <= (x"b0f564a644e39364", x"aac04853ea5f743d", x"8affee3525224edd", x"92973287dce282f8", x"79a19579aae4bd3d", x"17bca8113addbc63", x"cb6091880e12de53", x"8662be590fd32ded");
            when 17427283 => data <= (x"34484f520509d742", x"990650ea8fd77278", x"4b50315769462702", x"8d2f5ccfc3691d31", x"d63e72e5cd562632", x"4450b4b520b1f3a4", x"31a92f60505fcb8e", x"f70f277541bc909e");
            when 31034953 => data <= (x"2fe585b0dacbe47a", x"fa528f919c762053", x"f4a353b056a19234", x"5bd51e6156b05cdb", x"1c907dbee872a750", x"f8b79b02b80055c3", x"aafc158356d00aef", x"48e3d9507053f3c5");
            when 21764739 => data <= (x"06f302c0834a5e24", x"1ddef4c54a1ac10e", x"6068ba4eb2a373b9", x"e6a741e6871b17c9", x"13b412e465464c22", x"54793f3908740b1f", x"d5b07d72ac304d33", x"b8dc067015fb3ab5");
            when 2910370 => data <= (x"d3a59a7e4acb4692", x"2efe3166759abb2b", x"80ad182986c5c3d5", x"75cfec6d2af02824", x"00b8c93c1cdbf948", x"a714d62d4848d519", x"1be2784b50d4a478", x"7bd7e8331f33f885");
            when 15188995 => data <= (x"77639122f80f4e10", x"2a942cdfa0762461", x"0a0f7cbc4523d779", x"c03056cc69c6f0eb", x"bcf2689cd72fc618", x"8ee1d30f4d29873c", x"a4b14344e19d052c", x"b1035265bbbcee4d");
            when 33205817 => data <= (x"194f28464caac9c5", x"73b13950c48a0060", x"a02b82a5042d4ad1", x"766829725866860c", x"cf2677d77dccdb92", x"22b913444693ccfa", x"f398159dd8b7d3ed", x"82d0cb231855a3e3");
            when 1539403 => data <= (x"9c32983f88d94027", x"d30898b2d2723992", x"76d128b61f7f48a3", x"133c071615db3b99", x"6b24c1eb2e0b428f", x"2ebe28503d6e5b08", x"b959a57b6ef6ec5f", x"88285bd5b2a4175e");
            when 18051724 => data <= (x"d68e3477be0efe64", x"f954bfcf844c26f2", x"853785b86202a4d0", x"21f65f665094d3aa", x"5cc6db0b13670177", x"76af3f8f3f659146", x"e429cbf83f759ffd", x"2bd054fc72c9c214");
            when 13101363 => data <= (x"dee15c6db32778f9", x"017ff2f90e7d04c3", x"ec0a1838dff07480", x"47a364f22aa0527f", x"015e6b51cb35a59b", x"63f0faf46c8cb054", x"5899cf90ec2cd3d7", x"1baa79af588f08fd");
            when 29239036 => data <= (x"b0030df247d02a38", x"491b22dc30eeec9b", x"f8ecfe537064772b", x"3aad4823e997a48a", x"3a8781779891814b", x"07e9ec97e447902c", x"63bac41a66764398", x"04a2ae1de8393fe1");
            when 18688078 => data <= (x"d57057529c4f9bb2", x"c5f2712199639ee0", x"f825654892919e23", x"2b4efc3d9d6776c7", x"a8620bd21f9a86a6", x"3548907e47f7e5f3", x"2b9b4aa642485536", x"28fce450168cfd98");
            when 16269962 => data <= (x"d8018f7013af719a", x"cbda76ccd6b5942f", x"066e5da72a25dd9f", x"4b94f054f89dc0f4", x"56ba2c5b1c0e10cb", x"c6bb3705596c29f1", x"3d87dc9cae7c389c", x"2cf5dab8a73ba1ed");
            when 18026143 => data <= (x"5092db19d23c4b39", x"8511e5b5677c5caf", x"2924c83684c1057f", x"db8042da8dd79ce7", x"c43593a666e2d14c", x"d60e6b0c75513267", x"7691ab493b2ef3b7", x"08c9b0b3f606b3bb");
            when 18381637 => data <= (x"94db6983533bc6da", x"b0ffa98c026be34d", x"adb2ac713c02beb1", x"e46f602b37686dcd", x"42c52ced02281a72", x"63d8e7376ed028f3", x"a755471530df9a3c", x"168410300b51e972");
            when 12015850 => data <= (x"619671f9775a905c", x"ce0d7ca47c867c60", x"5cc3bbb47b1196df", x"1f125bde1d18183f", x"26a0b5c733f9418a", x"decb96b762cc4ecb", x"cbb1107357edeeac", x"e5196e0c6dbb281a");
            when 11937554 => data <= (x"c23458a1ec263b70", x"cca118d27f914e9a", x"0342081fdb885453", x"681d6833ea314eb6", x"594b85b2cdee96ac", x"bb24a93c334d06ac", x"9dcb7d56e80f4431", x"b60dd93b0fdc66e2");
            when 8831273 => data <= (x"8982241748685d09", x"99981c0e82d4dc93", x"ff8abedece17cdf5", x"40027cd1626e3bde", x"65d9ff920575a22d", x"28a3d7c6e8a72c82", x"7540daf6e3d5883d", x"ebd0e869b785e8c1");
            when 28215151 => data <= (x"3fb3d67ac76652c1", x"6f87f40f8dcee975", x"3c55aebec952e10c", x"1b2f9bcc84ea6b52", x"7daee3d7114e70b1", x"1eb0fa763ca4d1fb", x"c1f14528008e4370", x"9177e807251792b3");
            when 14257440 => data <= (x"883f42ca197642d8", x"63f4fff6f9e52d6b", x"a690f4d4a4bed56b", x"d672d6bfa9906748", x"8da4429275f59033", x"05c7f95237c8a4d4", x"d8a25ca49ee50635", x"c05df8f3d31b28b9");
            when 25677560 => data <= (x"a84fd54f9f4bf06b", x"0b4c6247520d6c4d", x"245b635a0e91dc1c", x"b822a6b6ce2e6a85", x"43ee797230c167b9", x"5d90793fb583dd54", x"d35b07074f92bb01", x"5d212a750cba1bb6");
            when 33480559 => data <= (x"245dd701645d92b3", x"64624ade583ca8db", x"316b80d7de901fb9", x"aebe8c59ad147a60", x"235faec5aa9323ef", x"72a4c9e3498c6b76", x"d5595a329e4dbfaf", x"71e3501ae64b47eb");
            when 16832024 => data <= (x"c89e402aef3491b7", x"fbccb2db2dfea0d0", x"eecb1f5d290028bf", x"6f3d1ac47ca6a6d5", x"a2de952ce16ac351", x"d1bf2cfe65f1d44a", x"45e8c9114919ec75", x"76d5574dbf80965a");
            when 11910948 => data <= (x"d7f6a59a79b18bd4", x"6f3a0ebf009a0176", x"2f5bab3b3e5dd817", x"efe46f34e649cbdf", x"e8edef8a2cccfc77", x"646b2e2b5fd4a104", x"395df262ac0c9c2f", x"de899dd8bc0f925c");
            when 23327043 => data <= (x"09a8ed528bac0e42", x"18fe6ff1512a560a", x"7516cca612731224", x"73da883af265aa78", x"0bf6b3c3892a6078", x"bbf43f582dbcaae5", x"12372f37b828a63a", x"9360daa75126ffd4");
            when 12225425 => data <= (x"0909a241d566987e", x"e8a8480c1cf09399", x"ffb7af49d7957261", x"dce4e0e415b02ad2", x"051408681a3ba25a", x"e7eaeae31adcdd22", x"37056794461f7be1", x"9fec6886e211c5d6");
            when 25927293 => data <= (x"d812e26002f90451", x"be2a8d3c8e170a93", x"fa565578572f1ae4", x"c792dc17cb88d0af", x"1682ddd2e7d3bb74", x"3a5f02a6ea9848b9", x"2c9fef73a0854098", x"09fbee2db56d3e31");
            when 28454254 => data <= (x"70798b29a08ae0b9", x"b31f45ff019c5637", x"5ef3fe2aecbedfd8", x"84350d247527c5bb", x"5d822bf6d99ca698", x"e49bf2f4d75b9d8a", x"aa4c49a632246fd2", x"dd4d992260644006");
            when 3037974 => data <= (x"70023dc68d25fc23", x"a318205700e7defb", x"1523198f16ebe944", x"c19a07ee52d024cc", x"206b2e4a9d6bb3e7", x"4d682d1ba499facd", x"cdd6f9794cd0aad6", x"c70a8a5ad0a75314");
            when 7287975 => data <= (x"553aeb4315008332", x"75735d93cdb44bb0", x"8cd8bcc65727b2db", x"3051ab7e1a7ad65f", x"0a3484dafa9ae939", x"58fe6c03ab45c02c", x"ccddeca1e4a6010d", x"23af6e16f20839e6");
            when 9883393 => data <= (x"38082459fb7a540f", x"0d5a3e6437f3793b", x"5b36df9be767966e", x"04b305c364233b7b", x"18522db7475ce228", x"9120784cf25b5e42", x"574f7a690b3d504a", x"aa1203d30fb1be0b");
            when 4403076 => data <= (x"1f4a117c574b5844", x"db395e8ed9e9871a", x"d1b56ac6c6f8b5e2", x"4ddd08fe229ac290", x"b761b399ddffdf30", x"6415febbaf0f87e3", x"ef2aed927aa87353", x"0864014173e19d51");
            when 22273340 => data <= (x"05b8749f27323d20", x"bcc18dc32a9d0609", x"9785176df07baef3", x"8c9af4bff48785a7", x"21de30b835778a63", x"f9c7c7a1e2ce8087", x"80d06e001e856d6c", x"091b709b5e0514b3");
            when 7357943 => data <= (x"2a07f8f81789c95e", x"a44d2617f27bb93a", x"347b8f921377c929", x"aae235e6f92157dd", x"11c0e27ef58b0475", x"3942a5b54b1750b2", x"2a28c5ed42e20521", x"a61dde949b6a1046");
            when 27872272 => data <= (x"3372ccc62de29433", x"a9bbe6b9e1560b10", x"33cf2ef7b172db13", x"79937026c0c4b2ac", x"10e3273280ca1772", x"7a711de91544931b", x"d982d4a98c9648b8", x"fc8dda4e6667be57");
            when 7389049 => data <= (x"46a01b82e67dc359", x"de7f8fb517187473", x"809c4702ea107785", x"ca88671ffd5f2934", x"bac19d9fe2c33095", x"19fde2d60f8f2118", x"63c21f4376ca2fc5", x"2a2c92a074b9431f");
            when 21306590 => data <= (x"22180cd5b4f508b3", x"3b29d3093e5baba6", x"4ba34f35571b2485", x"f8122f2834750591", x"778304febc2e81f9", x"5301f54a57589775", x"c3df7ab91824ea7f", x"b938c4cbff850904");
            when 29601308 => data <= (x"7c1da759545cec46", x"9e3a1dbd5ae915be", x"33a64d4659209bcf", x"039b963b2024224a", x"07b55b14d9dd12b1", x"2f0f9ee11bdbcac2", x"aaff1c86a8d6ae62", x"646e44790b71df93");
            when 9527991 => data <= (x"c7a00a91cbeb89f2", x"b3fb74d5d283c0e1", x"f4262226d1c23681", x"78cfef5e4d1607b2", x"ecc8d23071da4699", x"424972b7d51890ef", x"c428ab823f00b7f0", x"05a35354a66ebc6d");
            when 15331672 => data <= (x"0548d9e42bf53486", x"51d8d3af87d05c99", x"97266dba553fe80f", x"23ab684d1ae5c84f", x"65d52117aadbdcb6", x"6f393c55488bf93d", x"0aa7c1eeb423685e", x"7c4f9b7f013c6356");
            when 21220034 => data <= (x"764851c6e90af4e3", x"a9d85bd5603355b7", x"49205e3849760f72", x"bb93ea5411f023d7", x"98d39cfa968d490a", x"6e555b0dfe171304", x"bced4e2a88096720", x"c970322ac83c81df");
            when 6735154 => data <= (x"4bbb7ef33fb0de93", x"e8522436e313ad66", x"5f5087be7a4efda0", x"8559cd4e9b3ea160", x"7755112bb7d25313", x"0a0b863b2a22454f", x"ad29ffb3063cd7f2", x"2b551180ff72b3f7");
            when 1612774 => data <= (x"ba4a109773ea330a", x"6d127ee4cc18f8fc", x"bf274573b8715794", x"302d3b3a2734b1ca", x"657491ab4bfc7025", x"9c2999f6092c41a8", x"43a18e0bb130a45c", x"79e3704bb3c796e0");
            when 2916356 => data <= (x"2fecce85244db2e4", x"a39c36a48ffda27e", x"d1b12d7b96285430", x"cc49c4d366b0b184", x"cd47e998692fe02a", x"593924c8d38059ec", x"a1ae46663ac8abf1", x"690bab02589b0ee5");
            when 16776793 => data <= (x"13ba37870661e8bb", x"580178311ad1299a", x"a063f8fa198afcee", x"e447965e0cc73168", x"474a249bba080b28", x"65e86a30366bda62", x"03b21822694525fa", x"a4140f96d4557f8f");
            when 17472898 => data <= (x"001c47decd39b13e", x"8593c0a98f38071e", x"6186cb58ee0b4611", x"5d7ecfd1b67f3f00", x"fe0a40ce10228d60", x"5e82cb5da2b3f482", x"7841d0c779d82ae0", x"fcf8b3737e481b45");
            when 13201633 => data <= (x"f45e92e460a93f8c", x"3fabe0a9a25b8a81", x"03d0e0a21760a4bb", x"21935e54582c2fda", x"11239025be8e3266", x"cb7ec2dc9f7e699d", x"0810d8b74cabc120", x"7de7a3c3f931035e");
            when 14407713 => data <= (x"2eaa3845c88afff4", x"4962bb57a2f9fee0", x"532a998d5fbf10c2", x"e4fe6b9d1a1c186d", x"67e876169057542a", x"3cdaad8b91f520b3", x"8bd077bb4b89f66b", x"c994f1417a006b68");
            when 20948974 => data <= (x"8702558320b068a8", x"a3aad18bba5ef468", x"098aa7ccee158efa", x"13f02d367901e577", x"3f1394afb6ce01ee", x"bc3025f95cf1e68e", x"a9f2b543bc0fc710", x"33d6267c7a6300d6");
            when 19310264 => data <= (x"970ab0c2325174c0", x"190d1342393bb4c0", x"f42fa35107460d43", x"ef810a6df784f423", x"ce752d4f03594f18", x"016fc41acc0afe58", x"9f7358cf8044c279", x"d467329db7854f15");
            when 7968052 => data <= (x"a6ad21dd185aa783", x"089ee90a9d7de1b6", x"d935f94b55c7fc25", x"ee042e0d7316ceba", x"f7adfafd8049831a", x"2cf074b5f41e2c02", x"c11b273630b5669e", x"5c65789238e8a9b0");
            when 31573845 => data <= (x"6d7b6971d4a0d5ab", x"ac56aa83e9633e8f", x"c0e6d67f4c92a5ae", x"d15e43486f5aa061", x"2d90880b9364318b", x"c83fc2dff6f2287a", x"49cfb636cbdf4430", x"26cac6740ef70608");
            when 27257525 => data <= (x"410af442bd752f77", x"d97da2090ff8f5d3", x"f5b9961842902fe3", x"5ac1a59bdb24e4ff", x"6513a72d26ff5643", x"9f3766930a35cf51", x"c77f87ed13d03cb6", x"41fef919258ef978");
            when 9268570 => data <= (x"d727537b04f8bb5e", x"7f5f4eadfdecb3b2", x"7a8614dfa160e611", x"c76ee4f94dba3bfa", x"e3886feaeb3fff49", x"e6b5cec7c750a89e", x"ee46ea34826d4dba", x"d799f20a246f6804");
            when 10050702 => data <= (x"71248d365cb88b7b", x"0ba70c76e8a450e2", x"3f8bd10dbb65b086", x"6b5fd21759c280f6", x"060a0168e24ddae9", x"367fd26390ca143c", x"f263e8688b37c7ae", x"f14d3f872a6119ef");
            when 20577086 => data <= (x"ad78d514532fd1e6", x"0de6e03186fbbd45", x"af62cdd8750097e8", x"248e52d0b3748a3b", x"3a3fb2a52888745d", x"68d3a37f714d7b0c", x"d947b31cc0894ebb", x"2d31c1cd6f84ad31");
            when 2030241 => data <= (x"abc7d0a41692b01f", x"fd21dc6edfa899b4", x"edd004c6c2efb3bb", x"92bd328f7050b547", x"740d1147312a8e55", x"4d2576e635644948", x"28ef426a48d06c98", x"ed44d74ab254115e");
            when 5839341 => data <= (x"9a8b364e7cff1893", x"13affc670bdacc04", x"249cb93ee5828d7c", x"07bb9b409663adfc", x"ecbc5624962f421b", x"d784fd77ea3f34ce", x"6eb39b408e2d410d", x"c1e7b991e6903a35");
            when 5660379 => data <= (x"4919513ce79a56f7", x"1488c955f18d1ace", x"001fab9450c77435", x"aa02cc07f552e312", x"2a19a30ee8116cac", x"d4b43eda0f6e36d6", x"ad343f3186822057", x"9032a9664a7f2b32");
            when 14027859 => data <= (x"351a4e5218deede5", x"b9f67ed0fbdb17ed", x"590bd22eb52c4aeb", x"c3796e43d3806871", x"ba718d0a8540e015", x"9dac699b73eec7a8", x"b496432f940704b6", x"a54889bd37ef28d0");
            when 27870214 => data <= (x"e6359e8fed969899", x"160ebee9f41a89e5", x"cb842e06186cf7a1", x"34e3773aef5a8cac", x"e92efbb90082857b", x"a825df047db10912", x"7c578ef676f54a4c", x"655edabf8e15139d");
            when 20703738 => data <= (x"a5be83f297d40431", x"da27ac11b588d3f7", x"bdd678b1d67daa84", x"cbcfa7b4e6581ee7", x"69bab7710962e839", x"9786750aeed64a80", x"9f353d8f0ff99891", x"71678c28785a003c");
            when 31101451 => data <= (x"4f8a22faa83c390d", x"92b88cacc6ee9f7f", x"02685dcbe87627e0", x"ad4794e6f65bb0d5", x"2b45658ff6871f9b", x"8f303ed0af32baf0", x"1585085b68c9b030", x"ae10c238663ed982");
            when 31015631 => data <= (x"ab56d66fc79b3808", x"ca4fec136a32726a", x"9dcb43c1ef531384", x"88ead10b7db56eb8", x"a31455107a11e056", x"909e8712f5442b02", x"b003a1e2f8e8529f", x"fca31897c12a4c83");
            when 21522081 => data <= (x"0dbf442106361ea3", x"54a3969ce49cb22d", x"ee92d2dad6256603", x"201fb83e500b4ef3", x"a9f39037959760fa", x"c0a51bd678a1d8e4", x"dbccdd204cc46566", x"1f4c982ba111b9b1");
            when 22343987 => data <= (x"7efd7be813ac1c09", x"c5e6fe8dc804b90b", x"004f411915f6c8e5", x"c7dcafc3cf448ea9", x"1ac69f03aa1e42a6", x"e0c92b7183c80e83", x"cee07899bb9db68c", x"c5677dcffecb3eca");
            when 28960309 => data <= (x"e5e0717cc10a17a5", x"620d6bcb6fac9ae0", x"cb054cca687eb445", x"e258803cf7c45a46", x"24dd4263a758bd7c", x"54f0974c47a7d7e1", x"9cee9b3512e672ad", x"b0e423953ac87ac7");
            when 28709994 => data <= (x"69f7a9186347b37d", x"32f476e5708a3608", x"74adbf4ac36f0557", x"5e45468381ba5f52", x"232da3ac20b96574", x"45901cd39b62d431", x"d79207ac55704f96", x"930ba0ec820c3d96");
            when 13259945 => data <= (x"4551d18e03e97cea", x"6896fa8856236393", x"00817f6475595d33", x"3b39d97ef3462f4e", x"5bed7f61f99e8630", x"f908b742fdcb1d82", x"c7134c1dc3158b0d", x"e8da8fe7efdbe3ef");
            when 18090411 => data <= (x"a502c43a6017c839", x"4bc755c99ff17771", x"9a7ea4557069637d", x"91449ac9d4b282b0", x"48ddfa78361c269d", x"07e1a5f91615c0f8", x"0263df240d64bf31", x"1bffa6ecc71cf548");
            when 16169268 => data <= (x"376019b95c649fd4", x"b9c7be28a83f8134", x"745a147ee06cd782", x"89a931969745e901", x"486892d1e2c4ea09", x"a1f17743565e09c8", x"72fa2c5b7a79975d", x"6e627a329c88bd67");
            when 30619547 => data <= (x"f9b69927bd8b770c", x"cd9dbce8b20688ba", x"be91556181a3392e", x"34b2194b3bcb9ade", x"6c4b6a9c764f8bbb", x"20f214c72ea9958a", x"df8a2cd640774207", x"6b35390a0589345d");
            when 13321464 => data <= (x"8ff4a820217b3f9a", x"cb20cd81fef07ac4", x"58d006461f6c512b", x"87456db1f08c4f2b", x"342e9782f7cb2cdd", x"c6ca8d3bbc4a98d7", x"9afac6b74e11b134", x"98ab43880510fcfc");
            when 14228328 => data <= (x"4808fa14de1f2205", x"224f61a9d11b991b", x"2b44bc1a8521bf96", x"a3652a50afefc11f", x"2648b4fbb1d02544", x"f3fa4b2b4ea06025", x"d1ed38998bdd23f9", x"32d8103baddcd61f");
            when 16549349 => data <= (x"7c9f2c722a4ab0b2", x"d1effb1fb7c8e995", x"3a7d47ddf53d7284", x"8d0cb2797286f849", x"558824e91d6a167b", x"92129f91bb79dcff", x"6a05c39ec17b4d39", x"8c601c99dc9536dd");
            when 21633823 => data <= (x"3b202ed28badbaa1", x"6c5d1815a271f226", x"33260fffffe6e103", x"a9085c0f4f68256e", x"6bb2ab1f2cfa3cdd", x"7ea6224e9afbe08a", x"cc205a662c2017b5", x"a1a4c686483e08ca");
            when 1934489 => data <= (x"40c550e8c050afc1", x"c325736c2ac9c17b", x"cda68753307999d2", x"e517a32c9aa218bc", x"237401b6a48054a4", x"4ca533ca37de9a1b", x"219cac83291a221c", x"dc289d1f14263a2b");
            when 23740773 => data <= (x"ee367d958790cabd", x"cad7f306d06d8a14", x"5b4c838dbd02c8ab", x"e770db5eee37d258", x"67d6150607a06160", x"7cce0931e0cde3fc", x"add88316a2499c56", x"ea6fa0f47138703c");
            when 21128233 => data <= (x"8a14b1e74e19b05f", x"7373c091657d8a59", x"bde28d9f2d5dd315", x"c5c839d4b9ddfe1b", x"0ec87beff9e7125b", x"25b8146df284f87a", x"f2cfc5a00fe90528", x"24a502adbf517f60");
            when 4781830 => data <= (x"117b0aaae66bc9f4", x"3e98b6dd98374471", x"d54de1d76868320c", x"eec1cb38c3aa6846", x"a632cda071b06847", x"fabbe8c56ea57d25", x"01da779d5660a9b1", x"d31552d12e9963e6");
            when 6529664 => data <= (x"8e40e50f0f877722", x"9f9846d08e2c2e14", x"694cfe8fa6d6a2f8", x"3404c52bb5099c69", x"ea4ae0cb4d75f62f", x"19f5900067f970b9", x"b1403ac71edf14d2", x"51dd48565fa8aa25");
            when 11055925 => data <= (x"5f06e008ae85d8fb", x"56e683fd5a2d8b27", x"b1bc6d08b5172fb3", x"d3d2ec5dba26604a", x"a07c74170a871bb6", x"3acb19e49f53a808", x"af49cdd8c0b535c5", x"dd6cbd1194394a47");
            when 8385789 => data <= (x"7499e7d15b819e05", x"65d585c4250843c2", x"15df56001a89d687", x"43a71faa2b70d13c", x"d49ffb45d0c2ff74", x"81d8ba1f4dd1a9af", x"d4bcd663ceb20bc4", x"ea8b9be2b693e1b1");
            when 15071601 => data <= (x"a34765357b71d5c2", x"e412f1af11d620af", x"b9a091d87a347e1c", x"301cc28c68b1522b", x"994e71abdf12da3f", x"b778d3f4d1f91cfa", x"e6c6fe0c9002b5b4", x"f17ee52d5324253f");
            when 12258268 => data <= (x"cb7e72f2443e09a8", x"c4e616fd780da023", x"67003708f1d6a731", x"13e5ba0fcea512fd", x"e4414271aa449b64", x"f7e586e563ea5bdf", x"efbaac97f92cfc27", x"85b3d21ecc7bad23");
            when 6934370 => data <= (x"8648529904fa6737", x"67a05966053979ef", x"c6650d1cb279cbda", x"f73f21ca4e699841", x"6d91af50e9f0195f", x"d9d87d2f0b2f7eb3", x"0de9f04ec58345d9", x"40382e7a2b179315");
            when 13042322 => data <= (x"eadbb2e2f58e9d6e", x"2a4d87a9a8b02fdb", x"b877dcf60415f2e5", x"164f46739a7f55f5", x"868a16a944d4541b", x"451c13b436d624f8", x"2ee6d2fe2b65718d", x"270c13d3f6c6eb51");
            when 15682818 => data <= (x"fd3c51812280798c", x"3c24e507a752fc71", x"5b32d4409d422503", x"1d50dc6f6491f32f", x"f6222a4439620d5d", x"0c562d7dab156d4e", x"cdd2bbf3656e9c2f", x"79bc80896238e257");
            when 15602025 => data <= (x"9d1b9976f285a240", x"675bd1785edb67a2", x"7b73c9285a02361c", x"aa9907e58d971480", x"df79d349562df5ef", x"ca45279ce0a84df3", x"0bc7fb3a0fcde158", x"ed6c4dc68a3bd229");
            when 13759641 => data <= (x"b1174dad03c293a1", x"a2989223dc585899", x"2e3961f5edd94190", x"e1c22d38f362c046", x"9a0523315ba0d45b", x"9f9fa3df2af4ff1b", x"df07934e01ab8109", x"c7d6941297af1a16");
            when 26559128 => data <= (x"b81996afa7baf63c", x"03cb2d5033a1f36b", x"26188dbbf417beb6", x"e51389433bfd6f54", x"d104939557f8a39d", x"da69e08b40f189ae", x"48074be9a8c5004d", x"ea678e9a1153ae5e");
            when 8493888 => data <= (x"01eba2418e489e43", x"85c7e62275685add", x"96d7fc3b14e2755c", x"8235a4c00dc3d1a6", x"5e1e16b81b1a0c42", x"b16ef3196b7986c0", x"47657ad237f62274", x"b7a70b72c0ddb663");
            when 11604832 => data <= (x"55ba0d9de41e51fb", x"a73cecc93b0bd2ec", x"c5c5a1d122839c9e", x"bfede1ea13f4ed04", x"157b6d23a12ca51b", x"435fbc68d3497749", x"c7f36a9887b8c4fa", x"fe8178d59065b726");
            when 26665462 => data <= (x"afa6d346fdf26f4f", x"2a9e075d16959498", x"a5d7c47bf3fe7d57", x"5d2f04ad9fa42248", x"e1d5ed353bb545b7", x"a400091a03b8fd37", x"35472517f7391d6c", x"1202137bb4b1bb25");
            when 26191870 => data <= (x"25dd7c6a4cb1d995", x"ebdd22e8fcde92e6", x"48328959dbcd3c32", x"d25818cdcda73fd1", x"89c9e764aba658e6", x"3244d360d7de23f0", x"fb0680ae80986331", x"86c87fb1a39f6b8f");
            when 27367910 => data <= (x"a92f6ec428a893e4", x"827e58f7a9299023", x"b77301e64e90fec5", x"7d3406af9b7daf83", x"bb288be7c994c531", x"11a937a4bd4c9c92", x"030870073e88de2f", x"42cad4a8ca2b68da");
            when 1012561 => data <= (x"ed466d5501fa8240", x"0bace652eab269ea", x"67bca4baee5614a9", x"ce451b0009408711", x"f2ab68e63f246bca", x"dce989fab6052946", x"585848ff39479e20", x"da6af67e469a4e4d");
            when 22957775 => data <= (x"005c9c86a92c9490", x"e470d85b4a03f7ca", x"2a6c05971bbf33e5", x"70a19f07520ad1bc", x"ec42aa9e718caf0f", x"74f07e6df660efb7", x"c7821e717d83adda", x"da8c1b68cd4c27d5");
            when 21436897 => data <= (x"268c7fe89f772a34", x"19f5ac1e44effa41", x"3fd705d907443ece", x"521ae5a7c3ef68cf", x"ebd991ea900465d1", x"8de3d47ee92a768d", x"080e7527fd83e4d0", x"858828bf5baf315d");
            when 19842258 => data <= (x"6e54ea4c5ecd4fa7", x"4c93a5807d089388", x"0573e7204a22d0c2", x"cf294837b6e674c1", x"f40a9b775f32dc78", x"d03d5a20e3672b46", x"28d54fb87c65d5af", x"53956b0e6747375a");
            when 7001975 => data <= (x"1bfe3a1b09ec2e30", x"a4e0f789cfdeba70", x"3d70d91d3cc84faa", x"974caf33108a42ed", x"640211dbee275044", x"911daaaba88f1df5", x"5baee7a9a8b02d63", x"e6290421ace028a6");
            when 6328571 => data <= (x"7baf354e6c47b25d", x"ba7780af885bf827", x"c5a99eb42d03516a", x"6f9019bb0e37a1bc", x"a6d8cb7b19f355d7", x"67f6fab69061487f", x"cb29f240e709baa9", x"11a6988d3cef4b92");
            when 1601677 => data <= (x"897e2050147a21f9", x"50570a5e475a3602", x"f77c79407f96c734", x"1cdc797c113add2c", x"ec5ce52b7dbeba5b", x"b1edb9fa595b58ae", x"4e119e2daf6e0016", x"555e02fabf07e14a");
            when 4665834 => data <= (x"a6f2eb0c158da0e9", x"f1a4115db6a422ac", x"1d4de1ebfab98831", x"8b559a991e1a9d2f", x"13fb3ce28d9aa759", x"f29886db620b67fb", x"da0dd644d8d7f6d8", x"658a7dfaa619e4ac");
            when 12842104 => data <= (x"c0e7fc11bf2f704c", x"c268c207caef771c", x"79d65b12193018be", x"b033d96ad5402a6d", x"c61a1e412fd4d7a1", x"f35e01807f79175f", x"e59b508e31bd8547", x"1b37b3628d085136");
            when 1350874 => data <= (x"272d4bbc20d68b76", x"9fbf6b31f9ab4c6b", x"d912279146d1502b", x"3af212478b33bcb1", x"f8e5306d64cb2f0b", x"840efba1e5700040", x"f49a4cf82437f2bb", x"472b01612daa1657");
            when 15549893 => data <= (x"26a8d485b23949d3", x"1b957a421a222c77", x"4e4257c57bd66212", x"dcae80fe821db995", x"41a345dd06213588", x"e57213a35d075ca5", x"eee708378f1e0bd1", x"4a78a50a6822717f");
            when 30360719 => data <= (x"96f058cf6cde854e", x"cd898914089e4f42", x"a6aaea3335fcc4bc", x"f796e21f9ee0c316", x"2f8ac760bb7952ab", x"6c4d1997c250e04c", x"7ac508252a6ddaf3", x"6be8b06860dd4ebd");
            when 32400337 => data <= (x"8a71dc911d6cdfc9", x"f7d87edb84008a25", x"6d8016c003cf91a6", x"a7351567d557b820", x"9ed4ed8473f9f83e", x"20d91f691b3dfb88", x"020906e1addf4211", x"bcddd3a5a6ef1f99");
            when 593399 => data <= (x"19de5bfd82ad54ff", x"9413c95d201d9ee6", x"ff7224f18ad6c21e", x"b12d5d58397794c7", x"38d1640a947ed4e3", x"efbc682e037b2621", x"5cdb2d1158fa6752", x"055a798485657b5f");
            when 16514868 => data <= (x"c56012aa49f552ae", x"ddad59556d7b1d0f", x"814c20c2503acfab", x"7d713480993f1409", x"e7a64496750c60d5", x"54560816f697d6d3", x"154433e209d924b6", x"bffc89b54d7edb34");
            when 17812022 => data <= (x"a6c1035e69d0e975", x"4ad113fb5484c9f0", x"f404089503c90e87", x"e123b2a547964e81", x"78e9a735eaacb9c7", x"7222f808f042b030", x"3bdc8db01da4785e", x"3a2dbf26126b7603");
            when 645131 => data <= (x"f77dc8e2c0755374", x"6d90b3199f1e1ef2", x"1b01beed6d65bf18", x"8b1277aac1692dca", x"9b8234d5d81c32b8", x"74821ef3669a0610", x"8bdbd3cca500597b", x"976a9208de3bedd3");
            when 22398445 => data <= (x"c34c85000512c73c", x"1ded441bd1de568c", x"9879d633dee84fa6", x"7f3b42c307a9e041", x"0c198230fc2c8b17", x"e2dfcd4dd5e18f8a", x"f93e485c21561f82", x"07044caad61e301a");
            when 32633062 => data <= (x"fcff20256feb983c", x"2377d06ebac2db4b", x"10aba41e4c2800dd", x"0d223bd7a4371849", x"55f8fa50e6b8790f", x"9968b3df1c96128e", x"8342051351d50834", x"e6998fa0d73dee32");
            when 16575496 => data <= (x"726f4dea4fdfdde4", x"71e0c7f676cc2a3f", x"151264e85f01edb1", x"6f63f299a3f84f11", x"ce1a1954c2521042", x"ff90dfd5d2ef4da6", x"0ee140dcbfb89c8a", x"37a95f30d4c0c136");
            when 31919309 => data <= (x"1dd57e7fa9aaa140", x"2f5430ac29bd24f9", x"3e284556986aedca", x"ae2ca6c1eab9adcd", x"c456faa5be185e54", x"b54a56aaee42b16e", x"2f2488f83d9b2541", x"f5788851a5220d6e");
            when 14197170 => data <= (x"4784db94e656f0ec", x"e42de5e9bb931cb4", x"e2f9c4a860109c30", x"dfc8ca1fceea5fc3", x"e09919e24aa32c9f", x"6224346262e9e24c", x"55a7b3985671499b", x"13fa51a351f57c37");
            when 4102152 => data <= (x"379e6e6bdd791975", x"d5cac7d9c5753870", x"b8f972ccdcbbdabe", x"51ee374a35cf3b91", x"26ee93423920b768", x"9ed61e123ac944ad", x"4bf7bb66c72e196c", x"65cf3238028fda01");
            when 5092548 => data <= (x"222ed33009e4e909", x"9491fbf6f5c9b18d", x"b01ebb61c9288c73", x"ae4114ddddd31fba", x"e01839bfeaf86e80", x"ffec7b97da557d13", x"30968147609120cc", x"707132e962cccf87");
            when 12272532 => data <= (x"bd434af5b968026d", x"d50274c6105b19fb", x"e3db16fb938a646d", x"298848850437eb8a", x"e0346a47c0c46f59", x"93e5f19ebaf15b0b", x"799536992b4584c8", x"71e156ba9e4488c8");
            when 20782394 => data <= (x"9b01a58895de2cc4", x"43f71330c5758684", x"d2ca599288bf71cd", x"66fa980b816225b5", x"6d1df7ab445e9689", x"af8a80db8982acdb", x"8015598a35a6c33e", x"256c62de4cc41173");
            when 31608019 => data <= (x"a12c0a2b596d0517", x"e255f3e5468f64a0", x"9d8f4ba092c408ce", x"2474f448c5aecfe9", x"345404d76a4d638b", x"fc7565901523d6cf", x"1e69dbe109799ddc", x"fbaabc7e63f97ac0");
            when 30049026 => data <= (x"8e791358d3f3387b", x"8133e02e825d9aee", x"eb79b0d3f0debf97", x"24bbcd1c6606e6f9", x"55cab9f5251b40d0", x"2d970b4bb89b8764", x"01386d2d8ed983ab", x"ac0f10019980037a");
            when 26463624 => data <= (x"851c598fad32a737", x"211f36e39011e9db", x"4d6a487e7ef80b46", x"0b948d73bc46ffde", x"78d0b7ede9f6a602", x"36d3cf29e427f512", x"5cf7f75ab07ed9ba", x"ef5ab68be9a05fe6");
            when 20940771 => data <= (x"c4bac9b519937649", x"ff38d71672efc842", x"b7dd6e1f3ebebeb6", x"38141250feea3000", x"48bd3b6f7076b504", x"f09e73389d2185e9", x"5616dc55d62a9894", x"fce6c72e532fb4fe");
            when 18996619 => data <= (x"3fc49ab30b8ee4c3", x"ee5dd11e6b20d191", x"19a8203a111d6218", x"d5f0b262e571dca6", x"9b6e656be4ab5d07", x"b1f6463a17d6aa19", x"06f98249a637d4ed", x"ee45b7fbdccb1dfc");
            when 28138389 => data <= (x"76c7f62186874b98", x"da9d0d3a6f1a09c6", x"33fd07e3b84982e8", x"c5e24a04f602870f", x"eae155f16b141254", x"392e6505f583ee14", x"fc2bdfe83c5247a6", x"26ed7a2b20f0fca9");
            when 16534977 => data <= (x"118a76c9efc5ac1f", x"d5577454eec18daf", x"2a7c2afadd10a300", x"f1bf3565afb4b90c", x"c61a544759ac2fec", x"5508cc6143974771", x"75513896cdd32990", x"7521dda5b4c30c77");
            when 23099511 => data <= (x"7fea45d0bb8dce18", x"244fe1e599fcda50", x"b9a6f56717f03b31", x"855a4933e82041ef", x"9e091ffa1611e671", x"59889e525006a516", x"f8657b5bae66992a", x"19edf0a78ce25031");
            when 23159034 => data <= (x"88f4b498c2c8e8ec", x"bab14422cdc3b434", x"5a6f87bd6f183ab7", x"802753f9c059e54a", x"d0ff36eddcbd3c87", x"f66b98c20562edd6", x"cd413b414544d4f4", x"6e710bcfc4ca5753");
            when 8644024 => data <= (x"96673f6e3b08de2d", x"407382f0016abddf", x"370ffe458d6606f3", x"5dd372e9ecfa4d06", x"131435fcde4f942b", x"2f3349c1542e56c6", x"ef9757e449ee9a1d", x"89327de863ac769b");
            when 20586036 => data <= (x"af0b00eba0fcf5e0", x"17e3c2fca730e8d4", x"09c83a4f14518be0", x"59fcf7651b8bd602", x"75f9e4d165f23fcc", x"eae76f3e6cdd81d5", x"e468e4a770828a2a", x"b3db2727325bfbb3");
            when 14204868 => data <= (x"cc5eca1279955cfd", x"3c3f8aa385980465", x"7a0d833cfb16581b", x"f648fc974e9cd7a4", x"10db4e9d22c3e289", x"f36e1bed6a59ea33", x"975d6435d89d9046", x"cf27ff97bbd6d910");
            when 9016273 => data <= (x"2ac8813fd2903fb3", x"9b02e166c662201f", x"5e37908180ce7292", x"05312e8678113d35", x"d2590aabefc6b187", x"9ad31f4cfda15332", x"29ebed25e4ddc388", x"334b5e3634715fbe");
            when 14784502 => data <= (x"7910af3508ce9761", x"4747f4953194bf98", x"e016c8c35ada8121", x"94d6eeed6d862cb9", x"be3bf089245b2bae", x"e8ff3e1d12689cbb", x"5f7a5761262a3a33", x"7ba971f8e807950d");
            when 8539289 => data <= (x"9c8f92169d2e989a", x"1ace5e2142cd340b", x"70c324048c0c1ca0", x"81134d4c18633f2b", x"4c342d0bc5d373b8", x"00f66858ef56ca96", x"2ed15b6ce5615749", x"ff47a984db54e372");
            when 16416247 => data <= (x"ba921e9f3593d954", x"cfd309ae6a03ebff", x"047ab4e806b41d55", x"51ab657137180d6b", x"42d39793a758c7cf", x"fcff7066f7408d05", x"6dd301e0f0623eef", x"5f41aec93feb8144");
            when 13519005 => data <= (x"88bfae81417dffb8", x"a5744fbcb8c8e8d7", x"02ba3b1b59bca5f8", x"d9f0bb1e476fe4fa", x"23f8af10f9834bf1", x"0a710dd92176e701", x"2a9830bee72afeaa", x"e0e536150350e6d8");
            when 10594099 => data <= (x"71da564e067732ee", x"cb409354f5deaa2e", x"7ee2ae907c779e4e", x"33bc7fbc1dc92229", x"fe02dbca21e86a8e", x"b204aa409dcfc37f", x"970531731eb62e04", x"28da887379b250c0");
            when 32299083 => data <= (x"fb4f936a793acad0", x"cfc89eba162acd61", x"f1939a65ee20278a", x"55b72c2781ef064c", x"a211ae3f9ce31ead", x"800ccab4c6cfcc9d", x"1ec41a568a716a06", x"d394619cb12ccfc6");
            when 8792027 => data <= (x"4a272d604d36aa2f", x"a67748f65943bcb4", x"e939b6c012c3833e", x"4aa2cff2f800f5fe", x"195f29a89fe51e5a", x"767955f97543c020", x"13d6f1832a3bcd62", x"5e3b956ce3204d43");
            when 13537162 => data <= (x"c8939115e99db856", x"b22ee48c26d32e09", x"8b3e8454c2ddd331", x"a7aede8e3a51bf47", x"168a47c5ad16b5a8", x"dc42c6a03e4fc4b6", x"088b56f088cb347c", x"4febe79d3369e8a4");
            when 26211767 => data <= (x"5db2500efa1140af", x"d6a14bfa5801fba3", x"e6edc0ba3de6231a", x"c7e09b7c5ca78044", x"2e1953c127a88f20", x"6f0654d0df5c072d", x"b0b22b7dfa57656e", x"bf8eafff6341eaff");
            when 29553039 => data <= (x"7968f14faf4c2a2c", x"df6f8e90905dba07", x"d95c5f92337d7a6c", x"1c6880d453c5f1b1", x"0671cd44aedfa102", x"1115a01fdea2005f", x"65d3117f0c0dacca", x"38901cd0202204e1");
            when 11229376 => data <= (x"06e04af66a8ef5c6", x"10d90de7ab3bfda6", x"b841a7a1e643cc9c", x"d5e235f943c5a5f4", x"062fe996c648a6a8", x"df9db96f4adbbb22", x"355490119ad37325", x"cdd79eb691d7c4d2");
            when 15406421 => data <= (x"dec0160d6f8e6d0e", x"e4ac6f2d3762f7c2", x"e3050ece8244305b", x"ae5d75d7dddb48ba", x"8678843c0e77ea7f", x"850034cc9d8186d2", x"975924b814730e36", x"90c269e2ecb5d483");
            when 15443727 => data <= (x"dbf76a580a7917df", x"fc4d8c5479289e08", x"1a52008a66ed72c8", x"0d8a55419eb63a62", x"548ae9431dd24b48", x"27a3796d60130f87", x"73af83fa6dcb1cf4", x"d69b695831b4a5cb");
            when 24088504 => data <= (x"8ae975d0db4db388", x"67f4b3b255d7810a", x"911f4b979e5214c1", x"e48de08042d667f8", x"d5eda1c1b317372e", x"fa6c08d8608382d7", x"a1dd1c8933dbe12f", x"a72f555756d138eb");
            when 5230069 => data <= (x"681b7d65e28cb16c", x"f7e83b5ea2e27666", x"3746de923ee1510c", x"99e2aa5304e70734", x"845d2245468a0e1e", x"c4f69c6508fa2b22", x"fee347da02e66731", x"4649b13385a98f4c");
            when 24827277 => data <= (x"fe26573bbd893542", x"3f424de02abf3e10", x"27bad40a396731b0", x"0a455c260875a495", x"d30514efb76e040c", x"2b15c7da63f70d66", x"7c56b7932aefaca9", x"f03d81ee4dfebaa3");
            when 716845 => data <= (x"4fd29159817c0c98", x"96551331a478cc3d", x"09547b81bf7f0649", x"cdd5593a56c3519e", x"acd1b714ce06a15f", x"21aee6dac1db9d39", x"b70c2eca7ecdb8cd", x"0b85a3994e1cf9f7");
            when 33042766 => data <= (x"63e8f38a919b75d6", x"0b1f797e81659b40", x"250ff1e065714046", x"4e493bc787fac356", x"1f3afe76d4c3ee43", x"1e4eb736fb12879e", x"abe6a9fde25ff6c2", x"6183f077a268245b");
            when 9192884 => data <= (x"ca54e67e656f2798", x"0abd60c31f63bf3b", x"dcdd44f14cf14010", x"49fa5821cc3cf2aa", x"60647b5a542440c8", x"f263271a89d224f4", x"31472bd262b32870", x"629e37934eb1d1c7");
            when 33329531 => data <= (x"68d71afff098b0dd", x"e4886dd10e0a4279", x"45630d525bbfb9fc", x"e481f9a486ece5b1", x"cc5e186ee2f9109f", x"d1a04bafddf6bcec", x"21beb5ee62d24093", x"f1f6ef1587bed0a8");
            when 1637612 => data <= (x"4b0163bc033e8b4e", x"feec441e75fc2bf7", x"8d80c1868f3d5715", x"baa45d0a4ea9b345", x"16a483c46bcc6987", x"2a502342b8a9ab45", x"43fd324e47e57b98", x"30b2cd5c43d6f05d");
            when 33588567 => data <= (x"07a4e58298f23c94", x"e300680dd958ea8e", x"20722fc6373f0bfc", x"c82c3e5ded51a873", x"75a33dd774244c0b", x"8bd6846d9cb35a7c", x"478c9269fbcd9ae4", x"fc65407083ce25a8");
            when 8034012 => data <= (x"ff045ecf2730d1e5", x"a943590d50c5cd04", x"da137e3a83dfffb3", x"6f4bbcdc88123236", x"ffab41f952196a6f", x"abfde0ba5cce83c9", x"984717a218debed1", x"b656ea6433943ff3");
            when 7203126 => data <= (x"8666eae55092baed", x"ab708991b90ed383", x"07c85a777b5cea62", x"f5dff7fb36092186", x"02dbd3353a4c2f17", x"75bc5543f5d4bbc7", x"7188a190a3058074", x"81d718315c1e6e68");
            when 29084220 => data <= (x"6fb5fd64601d6490", x"8d0c8fd5f0c03e20", x"f4e68f767074c011", x"c973de7f00d4fa2f", x"c309a3c3d6425b98", x"17a1f7d8d693eedc", x"590fbb65ca254ee5", x"acedb402d3a4cb38");
            when 15913970 => data <= (x"a9e9307a0772b66e", x"b85e4b38b80f7cbb", x"8be7ed42e332e690", x"6c44447ef45cbc6e", x"7a7f4e2d33c74d88", x"8eacb73a5d877c6d", x"cb50b4ea6f8cb9e7", x"b9a2b89e5b81afa2");
            when 16768624 => data <= (x"87f73b39c90fadbf", x"04bc0a0803407ced", x"80427f5cd0bf5ad8", x"c240c8a5678a4b9c", x"2bbee60bd18d76a2", x"2a67680e5f7b8a4f", x"9a264f17788c7e23", x"5f3b44c7b0d2c5bd");
            when 13142922 => data <= (x"13870ed6f619c003", x"971c85b05ba22e79", x"fd8db2bac2d4de9b", x"7c612a5d8f370f93", x"3b408e370d464578", x"c7f6edde6d03118a", x"14b1be1a269ac600", x"1e5b3c5b833bb53d");
            when 5444249 => data <= (x"c482ec989eb023c6", x"66e920a434ecf695", x"740511239e128ab2", x"fec0df06291f5412", x"2f8ec1c98943fc81", x"4a94bc2fb02f17d5", x"4fdd6ace69c85f2a", x"7ce39093f18a5b6a");
            when 14833282 => data <= (x"72a53c2ad1338cff", x"873881b3ff748229", x"2ab7d056b16d6c35", x"3b069a1c73c8c8a8", x"cc1b7b7c05b26cca", x"b5a75fca632e85df", x"026d66f87398b6ab", x"eb7dbad4ff830985");
            when 30967928 => data <= (x"4431581a02c0c47f", x"3044da240544fe0f", x"7e71abd6977db0fe", x"9c2372f599b7377e", x"f9247283dbea14ba", x"8dff7a53506e2e0c", x"1f2f561a173df171", x"709f904c53bd1e29");
            when 31618535 => data <= (x"c576337eab769cb9", x"c7e6dbddc8eff6f5", x"20d144582c78b8c0", x"2b28a0a316732554", x"6ee09f83b9bef965", x"f72468217fe030ce", x"d04a911814fa70fc", x"0ad2bb6beb09ed11");
            when 26026137 => data <= (x"e2960ddbd8d3cdba", x"573b86ce21430d7f", x"dd2492e99e22c766", x"4444bb88af3c48b9", x"db70437165317fb8", x"80c865249dba6335", x"54093698f6e506ac", x"1a56958cdac9a23d");
            when 8663546 => data <= (x"ff5ea6c00f80f3cb", x"bce1c30f898e2b20", x"c81e07aad8da3139", x"aa3c7ee3b12d7379", x"c4f86b9dbabcb8f7", x"1265775653daa1dd", x"aa78b5dadce78c2c", x"68b46326e8235747");
            when 9243910 => data <= (x"0835914e1641854e", x"32681828b1c0eaaf", x"90a9d3a90bb8cec9", x"7c8f14c43a2e0ebc", x"599ff20fff5ffc55", x"e67ed368e9aad748", x"9a1b10ec612520e0", x"11cb4db71b356f1f");
            when 28742507 => data <= (x"0d2d825571cb6060", x"3d3832b9eb3a77a1", x"4f98f8615ae17069", x"10ae238d7e56f00b", x"47f3efb8001bbcfb", x"d10bb28acea9c8a1", x"b89f32210544f773", x"d0bf05ce01e6f418");
            when 4702921 => data <= (x"f29454d3a118bbb8", x"280eaa091c997bf6", x"3de3ec16e130fc55", x"371988b3627be249", x"6311a0b3ce04a4cc", x"1a0a11fc65004c8f", x"032d1b0d5d50554b", x"d18e6621819a57cd");
            when 9838429 => data <= (x"1a1d16a2346b4be7", x"e16ad0cdefe121d7", x"6bc83db79916ba7e", x"0ceebfa719ecf4a8", x"82490612728f882b", x"ae7693caa3e390df", x"0ceee3a511cb6d70", x"9a8df4f435279324");
            when 27900762 => data <= (x"38d6f13c76db5d71", x"96b0b1be34bf4d55", x"8f35cb99c482f665", x"d8abf42286282a12", x"4b3f67e372a46ffc", x"06bf413f22176f18", x"2510c73b551987ae", x"2960b6f728018e86");
            when 30044099 => data <= (x"9a3a500b0320ac7c", x"a9fbe55ab631cdba", x"b2203e4f8a14bb71", x"7675bccb4c30200e", x"30aa87b61e81dd69", x"74ca6c9fb0c0652e", x"5ea858b94c8cdefe", x"2282186c71078af4");
            when 33278537 => data <= (x"e3134eaa31a37448", x"55f543bbfad84bc9", x"c59ac936a9d78789", x"4a7833774ff7e009", x"405aeb7ca8f17ed2", x"e0f8075ca1ac7885", x"62fd187b0dc847fc", x"0d83b57603df5627");
            when 2197720 => data <= (x"29ff5d4f0800aad0", x"5b3235d6c2a95af2", x"fd60dbea73d83ae5", x"d59d6853b16f1b28", x"85bd5a5ef8e07a7a", x"9589ec9417fec1d6", x"92aae58839342fe1", x"cfd62188b1361acb");
            when 19831848 => data <= (x"d62184e90c60a56b", x"3b0dc4fd7fe122cc", x"56a856960215622b", x"16a01d9f0436002f", x"ab92de844a26e831", x"6571bbca77fb81bb", x"1d45b8bc51d3548f", x"86c3ef890fcea757");
            when 20686410 => data <= (x"e541142ccab30c40", x"ccba17c243f5afec", x"79490b5be4dfe3e4", x"3ceb8d7af09bc75f", x"eb8351135a1e7f1c", x"a31535f74eab8ded", x"c83fbd66d3082c0b", x"9f85a0f889d79146");
            when 1115205 => data <= (x"5ca1f22afe8e6910", x"1fb92b19f4035fea", x"1e21abb80c0561cc", x"5a7384002406ea9a", x"30a812666ad30430", x"dbc97ca1b21668e1", x"62d952e74fd7b305", x"6e798d8e30a79c9f");
            when 13253379 => data <= (x"60be115d638cb1a1", x"61932b123ae754a5", x"f9085a723972e14f", x"fd5f5871f4b33555", x"079eae427657a62e", x"c3528e3ccd3b2bc7", x"eceb321612415f3c", x"0ee9b84bc2818fde");
            when 12468147 => data <= (x"5645db485ece085f", x"34401342446c40c3", x"23841c9d311fd8cc", x"d45056d89a4ff2f6", x"60cb1f9d451adb2a", x"7760b1435955984e", x"623411f2741e7ae8", x"77337c60cd3fc11a");
            when 19049152 => data <= (x"a9b97ae535a3744b", x"571dbd6eb02ff824", x"a49cac6d4512ef35", x"d944559e34864c97", x"805d97e3928cfb51", x"776a5cb1275534e3", x"2345cd253006e764", x"c0bb6c15bafea03f");
            when 30081794 => data <= (x"a2196cdb2b5081aa", x"7b3a2c5223e900bc", x"a0d61fd6d34075df", x"57899f3f181e5844", x"3e3daf9be0c1ed1b", x"cfd2b1a7a95885ba", x"8015d0369282350b", x"20e5573ac172ccf2");
            when 6809192 => data <= (x"21e92abb27d6c953", x"8e166808d6a595cc", x"243b21a2e516879a", x"87e12edba4812fd8", x"e855b9e6e0cb7c9e", x"0044f5f879e2e969", x"a4faf89ca7756d15", x"f10e0193564ed636");
            when 5294402 => data <= (x"b8a43c5f5630fc7d", x"0c33a1323f84c60a", x"7056de3d188781d0", x"da17b30dd835b440", x"bdf994ecd2924ff1", x"1848b0936402389f", x"9506861af7546770", x"77627e19263d55de");
            when 17247080 => data <= (x"2efde9d13089be14", x"7abd3b41001930f9", x"01e9717d73c1d9eb", x"5b05afc6cabd7d7e", x"b5b3f47231041cab", x"5306e5526ecb7377", x"53114eb2bca5e0af", x"c1deabf6e5787106");
            when 23528662 => data <= (x"f4bc2be0f08343be", x"c52c7984e5cbddda", x"326ea153ec7adecb", x"05ed4fb72d13df02", x"287367f07cd7fe25", x"1dd353610ac2f3df", x"b759192abc3be42a", x"f1ad793932d8330c");
            when 25795391 => data <= (x"52acfba8e74d2388", x"a8ded5407a15bb12", x"822892ea9b9389d7", x"85dbc41ed567caa8", x"53779ac033d10dd9", x"0abdc6674089ccd3", x"a3367c039202c969", x"25be3a5ca4c3a6b3");
            when 32752090 => data <= (x"894e9bab990a9a96", x"c9227b6a674b65b0", x"b2d4a4fc6e9783f9", x"220525cc5a1483d3", x"865f8c69db7100fb", x"19b467c9370c9309", x"80d6c0f03c6ebc26", x"8bc91d1ccf774834");
            when 33375061 => data <= (x"549e0a2895cf4602", x"ff50e53475733c2c", x"2ff8f60a6d66d87a", x"3e1263107da57a76", x"7be154412aa0aee4", x"95c3810c2480c435", x"c450471c07d67e1b", x"6dc78126557d9008");
            when 8197812 => data <= (x"6c2fae43b6496b93", x"fa3561f0d6b2212f", x"1dad526ef39c51c4", x"7d3db2c5338f6dae", x"7b6c4dcdf99303d3", x"61aa288cb87cf059", x"5ca47a7ed7055579", x"c98797fb9f597a57");
            when 27159887 => data <= (x"2aff68ce6e74306d", x"0bbd4148ea7b1291", x"0432caa7c7429766", x"22624702a7f90df8", x"3cc17fec992c3645", x"314b7288306cf062", x"f3ef0bf7bce54e5c", x"9e21f2a23ef15e7e");
            when 7250130 => data <= (x"55a3b1c74a6f00e4", x"f4179168fe68f6d0", x"22930560dfe456e4", x"d42cb0edb40cad5d", x"e995dafdd7bef235", x"e24355f7b6cc5f49", x"4716c2a658906b51", x"6049c3cd9eb7c7e3");
            when 23651030 => data <= (x"93136c4f492db05e", x"b65b1b74c63ec26b", x"0819adc54f0b2c9e", x"0fd5e7fdfdffbb55", x"516950985a3d21c6", x"fcdfa79ac27f5136", x"a74dfc0981b637c2", x"f9f9f05321489caf");
            when 14263815 => data <= (x"b5ed7719f5101c49", x"7406066ef5dbdc4a", x"4971ec2bba70c92e", x"addde73d0d5675b3", x"2ee7f30b8c987e52", x"c41c5d9e002a988c", x"bb06efc2113a49cd", x"ba3aa520f7989bd4");
            when 16711200 => data <= (x"00d6bbe9f33e7331", x"cf4f81960c67a740", x"d79145bccf8f0640", x"288cceac54e05e33", x"d5afa4e0c30f5f7b", x"41624646f573b95c", x"efdb893ecd86fbba", x"4b9bd6faebff5e17");
            when 29354038 => data <= (x"d5dbcf58e6b343de", x"11076b8cdaedaa4e", x"3242723a80f76dc3", x"8d5ae02724cccd2d", x"7dfe7b66b7f91a84", x"7e45dbd7fe021d7b", x"aba1f1a0aeea9d96", x"e85062c8b613ef7e");
            when 2861845 => data <= (x"371a104d308406be", x"e7d19a35fab18f03", x"f163341991335415", x"f14ad6070da92518", x"92a334207fb5c3c9", x"73d76a66ed692900", x"4c9cb57c38d7022e", x"ddab748a0df6d22f");
            when 7863709 => data <= (x"22f3c61db20e3ac8", x"73a2753110eefdda", x"8a749d2b32277ea5", x"b182849dbb5b975c", x"d99a5d6f8e9f6067", x"b676c034d21bcf60", x"53182e52bf8f609d", x"29a3b53aaad257e6");
            when 5174151 => data <= (x"3eaaaa8aeed58361", x"86e18bed84c18bcc", x"41c54de5f51685e5", x"fdb8f348bd6de383", x"3c1102e495077d94", x"6f2bf5ba3bb474db", x"2505d15efc53c6d4", x"9dafc6c88fdb18a9");
            when 20057234 => data <= (x"2dee008a93aeff8e", x"70680b6e45127a6f", x"9eedf906c0b76f46", x"b42fa3c25fc9ff29", x"91c4edcc4e8df302", x"dac094a9404fa0a5", x"4897b395863e27b4", x"df4403d9303305c0");
            when 17836943 => data <= (x"a5f36c40a188196c", x"2a92aa15650a025f", x"3348cc055d13aef7", x"24e76391bd623985", x"5735fbdd908f4525", x"fd888d698125edda", x"cb69dd594694a6c7", x"fe7d64abf3ff793b");
            when 28952661 => data <= (x"e9283b93d11d5ed4", x"71478872f1889ec3", x"1569d6ba75a74142", x"23b79515fe784cfa", x"c6ffa997bc3cd37c", x"83bd7a6bb7b34bb6", x"13ccc1f7c7dc2605", x"bffbdb9362d4a0b1");
            when 18423324 => data <= (x"00fd5a7c1ba9def1", x"6afab1b600755e76", x"422952929706ab74", x"f4396309cbafd979", x"910a2a005766bc43", x"0375a03adcf77c50", x"c94bd2eaea12b881", x"d2dd242ae0d76b57");
            when 4152125 => data <= (x"918559fc2727d335", x"a0ddbbc0fb512072", x"c75371114a41a104", x"853e0e91904afad5", x"d42f851c7d825e03", x"373c68d779e9f5d5", x"073466b9599904b7", x"93249e3ceb44f6d9");
            when 23520392 => data <= (x"f73ee89fc23cdbff", x"843840786cb7b750", x"c455c7cf9346ca41", x"e8b7371bfeafe68f", x"73f17e3e3a71aee2", x"8920eaf700bb18a6", x"1db73750cfff6e6d", x"b3c4954519ed7e79");
            when 25028877 => data <= (x"346cb84198ce1f26", x"d87c179e4a859d8a", x"363f6eb7cbdb2528", x"828321bfd3016348", x"f3cc9645007766a8", x"acd765a89fcab8a0", x"ba143859d47c867a", x"87be0f3093c7421c");
            when 8498339 => data <= (x"c9425bb87a96477e", x"4325414451d74eba", x"87bd00cb7ae3f382", x"0aba160efb24825c", x"ca1275f01297af55", x"06843bcd6b16a45c", x"2ced6c477b622a45", x"73dcd9f7579a4a4c");
            when 11163285 => data <= (x"5c1f3e6bae433a3c", x"6ba452d09e76f3c7", x"d089dbacafb4b53b", x"19755bca2db88976", x"57a17116553eb89d", x"f08464484f4e6912", x"7827d9e69ec4899a", x"e85177d46ca10ff4");
            when 30253359 => data <= (x"633f4d535c2fbddd", x"0b254203e3a967f5", x"7677d9528694a31c", x"8ffc77759c0f6ced", x"65546997b0ccca7d", x"06bddf9dc0868959", x"28d4dc03c981bf75", x"0a26e19caf282153");
            when 13989021 => data <= (x"ba67eeaf3ed4091a", x"650faccf7b5f7e13", x"75014dd282365f64", x"39a1df15c3c20c9e", x"93c79782991d1e40", x"cd1593630c008642", x"899a7e40978e0759", x"f5aa02f9078e0446");
            when 16791614 => data <= (x"c10c3fd6715c3b74", x"982c8af904c54a7c", x"e55f63e75dd25213", x"5b9c59ed27e9358e", x"d90dae567c937d76", x"02661c58f335b4e7", x"f895d9905eea2d66", x"27e7a4aea1273a76");
            when 11616523 => data <= (x"194766a4faa2f27b", x"f566bff42eb1b235", x"87c1d42a2b7c7da7", x"5661bc0ba519d74d", x"cb5f67041a45a22e", x"2b8d5f46fb3b7543", x"3eabd76a618bd636", x"0699292247f2a77c");
            when 27769496 => data <= (x"bb3da7187226156e", x"efe3ec7ac159c1be", x"4c05964dededa4c0", x"d6a16732eaf79732", x"b875ef2edc009dd0", x"2171b0558ddd3bf1", x"8354b03ce168b862", x"600a9703741e706f");
            when 15951100 => data <= (x"a36d4b1d329784cb", x"43502a528d59e68f", x"56e039900bf07bcb", x"55f4c1b90d2edc18", x"62fc2ea7736259e6", x"f2ef85d3525e9998", x"caba0d02abc877fa", x"b856f72db170ffcf");
            when 895487 => data <= (x"2cc709fc772c729d", x"4e2e92497400b3ea", x"713fa060ba60e59f", x"6746e9cfe01a68ac", x"8263067d2f70f278", x"386f9c0cdc893124", x"b4c6309d23ce417d", x"d00e4c85809b7c59");
            when 1222363 => data <= (x"851d012e66db4352", x"56b4e8ffd072e6b2", x"c8f7da204ada3576", x"17b05908c6a7b1a6", x"a9ba62f67eb46567", x"10221b2fb5480b99", x"e933289aea9f5c71", x"cc259e23e4f7a151");
            when 15204177 => data <= (x"273dc3c850586843", x"0c319fda102714c4", x"6b5f1a8169616411", x"15a5da9b96c9b9e6", x"66ade1fb0bb83c97", x"a4384ac22e04c4a9", x"00145007ab253b12", x"f09aba48e1be7c8a");
            when 26868191 => data <= (x"4054f274b04f554e", x"63054cd7910ab1dd", x"7350b398bfb87b73", x"92b6a0a2efb9c978", x"f00feed3e6de4f58", x"defae6fbf22b2de0", x"92968dbea70a0241", x"93d6147bec0dcdbf");
            when 31527305 => data <= (x"e31d719a6c439208", x"c306c7c47653acc6", x"4d3cc9302cfd6c67", x"50e0611eb7e2d861", x"71fbc9cd75d69cc0", x"57d0b55f2abefaa0", x"7167ea8bbbb2a22d", x"82de4ab8bc45b6c1");
            when 22357396 => data <= (x"3f51cd9980a75584", x"939b51e45a3be2c6", x"82d16d94a26856a0", x"00a6d8f67e25cbf8", x"94fb57065f539782", x"443b0c93b9d45b86", x"14912137cbaf12ce", x"b85a39dcf0025fa6");
            when 5594879 => data <= (x"92cccbc150ce3433", x"99c9e8b5585e7230", x"1c07582dba793f57", x"973795951d0ffc99", x"3f409cdc4d9b9a6e", x"d40a2f6013d8b3f2", x"658893830f2a2615", x"f6233281f47b06d4");
            when 24339578 => data <= (x"b3718998f4a507f6", x"8ccb2f081471eb55", x"bcd554acdcaa5d19", x"c1b00e2ecf49e33e", x"f15186179fbc471d", x"ca454316a5fd736d", x"7e30cb1127cad1f1", x"edc10b607343ae6a");
            when 24573562 => data <= (x"ce743205c1fcfb62", x"a97ae0a92b851e20", x"cd9922c229f47a06", x"49eb8e9ffcaf5a36", x"a7f6f16523275397", x"378654045412192b", x"8703f8ae2270ad73", x"8e1ad7a15decd357");
            when 9808295 => data <= (x"9e039d7addab4a60", x"f89876df35f31236", x"2f45eea5e5f19f13", x"7e24b2b5fcaed3e5", x"8257c7ce5dafcf4e", x"f76ed9cd3a1641a6", x"048e934a1f25bf78", x"4d75a633ea0568e3");
            when 22676128 => data <= (x"c22e419970f43d21", x"b54115476dc5f2bf", x"a0f28fc87fd7483f", x"5b4c952386569ffd", x"304d28b394a63004", x"1d3057e329b57d00", x"c5ce0071d3a48768", x"5366845dce13dae3");
            when 27600165 => data <= (x"619fdf0ad32087a4", x"e488a45a61bbf955", x"5ab5368a1d39777c", x"a87d788476473c92", x"37bf9bec3db7d601", x"75b3fbb7b867cba7", x"39235dd743dbaf07", x"9f269cd3482b51cd");
            when 25248172 => data <= (x"30b2d9d77e707ed1", x"fb95035d7cda5e57", x"bb9e5764b16ce871", x"09f41eed9da3cdca", x"0eab813089384cee", x"83c0514500819485", x"7b42a159d59de40b", x"37f03fb0e821bd0c");
            when 29336460 => data <= (x"852e16a0cc6ef16c", x"d2182b80b65f3478", x"53662d86aa8ecefb", x"3c15201faa8e02cc", x"1552f846900bdadf", x"916d077c2a58dee1", x"44e88f681c7c6e8a", x"5ccc293899ea9de5");
            when 6039296 => data <= (x"216e64aa71c2184f", x"8683784871c518be", x"f14b8844b2fd827d", x"d5a24ae795a6b829", x"26b8881f161ff8cc", x"96402f32d8f5d5cc", x"ad82396f7f8ae650", x"26f981e093c75b58");
            when 15659780 => data <= (x"2efa415d3e14c059", x"75f59553ca399a91", x"f1c42e695a9f1611", x"eef496d7a9b75da9", x"9f2cd373478af3b1", x"67470456f1e00489", x"fdbce9516b4989bb", x"65d4d01b2e893ab5");
            when 26775439 => data <= (x"389164dc150c92dd", x"c4caeb99e0dae2a4", x"d5c6231f806fb7f4", x"cce9c0d31a44dbae", x"62b6daaae44ce66c", x"a659ce6f9794a315", x"f30949b5a0ad9cdb", x"c3c0cad9d4e72587");
            when 29851912 => data <= (x"accc04119f18cc30", x"30c79125c78bd205", x"cd6bf37325062517", x"32412e7fcf0885bd", x"17a72ab3e2694ea3", x"868b62dfd5117554", x"2cd22367a7f47225", x"3369a40ede28a852");
            when 32622371 => data <= (x"2e188111b8f2475d", x"8b2e3e82e5a13c2b", x"fdd2edbc67552891", x"b7b1b0781c1c9c64", x"928b232d9a1cf437", x"ad21d283b3e2b7ab", x"ef0b8980017e9b45", x"d3d1419d977b3dbe");
            when 30795586 => data <= (x"405e740c5d74931c", x"c11f36add142bb5e", x"17cd42f6c5056eee", x"f23190305c1ab83e", x"6f4cf012601d53ba", x"0137412a99409f36", x"e23e3e7064116d16", x"7782ccf018d77be4");
            when 18291692 => data <= (x"e3f5c3b91c2b3609", x"66571068fccb039e", x"90af22b7752216cb", x"22ca21a5bba167c6", x"2face8145e846c2f", x"795b86819b25bdf3", x"47a672359d62a0db", x"3ac5abbb299be17d");
            when 366561 => data <= (x"1f6c060b6e9dc128", x"0dff184df3a2ea3b", x"6b8e9a39b82809e3", x"e3c415f0e86c6465", x"24aa122993a37e77", x"abb5bf043f4059f1", x"144e5d8e601571ec", x"27a3ec2478e8127c");
            when 1620846 => data <= (x"1f9fe482848afd3b", x"3d1059ce5597287f", x"8ef6d798ebfb941a", x"4dd194dfda5b3c32", x"b2dfa7d49f86b4fe", x"73f5607e4c54a60a", x"91d015cf8e209d59", x"20eb14f31d5ff21a");
            when 25382809 => data <= (x"8c0ac93cb27cd151", x"c4e0c514ccce10fc", x"2a9d1233ddabf8a4", x"9c83b19bd3b5e83a", x"30fcdfb69a565c52", x"62410bea32beb6b4", x"f241962148304d40", x"14ebbd1837dcc017");
            when 580354 => data <= (x"cc932f7e2fab72e0", x"1b5e94b6cb5e2ef8", x"f8701d28b588176b", x"8ecd697570f2f342", x"eadf2c7111e83016", x"e4cea39aebefa1ef", x"64cc6b9d7a2614e4", x"db8381cf2756c959");
            when 5412836 => data <= (x"135c563139fe4a48", x"22c95e7fa119c8ae", x"95fdc1cbfaa7c1b6", x"74c33f6997e6bb87", x"5937949315314cc0", x"5a53621c2b307ae7", x"622cc9ed57fe8c4a", x"82682eebbc5194d9");
            when 29326315 => data <= (x"f415e229a14d20b9", x"4a24a0e7e688ae03", x"951df1fec5c808c2", x"072bf3d7dd8e20f2", x"1ade1b1987960113", x"bc5f3b50208dc749", x"124d9d0c91036b04", x"572782630fbe8f68");
            when 3006775 => data <= (x"7905ca9e3ae9a797", x"5a3785428b41070b", x"504458a0fb42211c", x"cb4fd944d9a537d2", x"996a2c6fc22f1082", x"ceb1788be9577deb", x"7178423cd5d32381", x"d93430fcd2122a81");
            when 7201605 => data <= (x"4e10becf26d5fe65", x"304544a4c8c5dd15", x"e9080278ffc9cca0", x"1b113a9f8b7e848f", x"7ddb4a637eb99884", x"727ae35c67840457", x"bf6c13fdab1c8e87", x"8a8c9927881ac476");
            when 25590764 => data <= (x"f5c6627e2b5d869a", x"063b14061d2b3b58", x"d40745cd18ea0bc4", x"14b7a17fc58659fe", x"663691b6f5e99ac0", x"83d07fa7f92b5e0d", x"dba99906f8987da7", x"00f5280975d158ca");
            when 814547 => data <= (x"5f06600866bd42bb", x"ce61b30c2a90b5f7", x"4f53795d59a833e5", x"92cba7ac06e4a198", x"b79cdcf0e50deb4a", x"7bf197ef4f9fad04", x"c3e572600a30c9e2", x"b735f899c8644f13");
            when 24735388 => data <= (x"c221d23a981b9b5c", x"357f29055970816b", x"6e762b8cdb9541e7", x"b7e81b70720ba400", x"a2a3b592db2d335f", x"66dfd4e3329c0b4b", x"33a4248f7fcce873", x"9746c0e658f39af0");
            when 24361922 => data <= (x"f64085372b52f371", x"1afb3e8edbac28aa", x"48bb64d18173ddcf", x"9aa01a2ff2c1e7f4", x"372b908ac8b75495", x"edb98f12563f7164", x"afdbfb4882714fdd", x"9d02d1b89012b9ba");
            when 28477591 => data <= (x"e7370d4119db5fb1", x"f4ab8e504d1748b2", x"7a6d98d5e60b631b", x"f29fe3970b95cb20", x"0173a65ebf127ae7", x"867f9f20b34589af", x"d2932ab247b3f8ec", x"3a82a8c66314fe4b");
            when 29974664 => data <= (x"d06d4650208020ed", x"b8ef34e62f6f6b4f", x"6b997e5539635688", x"6842fe11a3a306b5", x"659dd650794ac302", x"68b9836c38e1822c", x"27628a19b094a7eb", x"fd786d1d2840f144");
            when 12322148 => data <= (x"f37fb8566fb3c1c6", x"f12f937fa45744ec", x"bd0dbff278da5f87", x"6e3e525d047a531e", x"07f7c3262a96a7f4", x"637b157feee90772", x"c000b5710cda42b2", x"4e4c7bd351174140");
            when 3760999 => data <= (x"efe48ebe9a187490", x"e45db5e53a481f92", x"d91c3a113ce441bd", x"20a54a315cd03403", x"dfd92594284ebfbd", x"f987e068a52791fa", x"7511e46106402d3a", x"4d7a0c35dc37f320");
            when 31261196 => data <= (x"e9fafc032dfe2d0e", x"244e3f8c505869aa", x"e7d4a7a626d8ea11", x"3e58be1abdea249f", x"73d4a68c34d8b8c9", x"7fcfd88df4cbabf8", x"55da119e3304f00a", x"076e7180d2ea48d1");
            when 1736072 => data <= (x"14387f160360e4a1", x"229825af4d03e715", x"63ecd1f279ab8d51", x"6a326f74d490d0d0", x"bfa9523cd22d9d12", x"3e1cb7ed3bfab3cf", x"6f49b28001eff208", x"55aaed967549311b");
            when 31209235 => data <= (x"af1f3c8e6473fe5c", x"8e5701afd1e46837", x"2ab245d243db7820", x"99f45084958c3c6f", x"65a5983e7ee65e6d", x"65c378147f6f46ac", x"3deeb715b901392f", x"7cbb7d4e23ca3c2a");
            when 8104187 => data <= (x"8051c3fe0f3a716a", x"51d6c99ed448a4f5", x"89261475cbc2cb43", x"a4ee7340bbc31225", x"1136bcf381beccec", x"c6bd9afa2c8720ba", x"e86fc39f49edf8c8", x"1dded70d2a7a65cb");
            when 365509 => data <= (x"e01ef12ab6516a12", x"938aec323d344698", x"7de73a69f73f492c", x"beda8d09a27feede", x"f66b910ae40b186b", x"72fe3cd344ea59c1", x"d20c252fc538a586", x"6939d6b0e21d0889");
            when 11877950 => data <= (x"bb0f44dead779315", x"2c8b602dad9b52c3", x"12ac665a35208c8b", x"688da7fd3b5f41a8", x"6b6be59315ae46cf", x"e03347cc0541363e", x"d394cf3eb05e491c", x"c964145654a6123e");
            when 9868927 => data <= (x"7083512a2526ef74", x"6f7ef6b23d670a5d", x"32545da0a8cc0393", x"514a6c70334c4eb5", x"c89b255b3b8ed485", x"5856fccdb334b083", x"09dc9db2c635af58", x"576c58e376151978");
            when 22991720 => data <= (x"c2c4fd2d4b9cfe04", x"6b0f5eb0af33cebc", x"dcd60408fc1de07d", x"02ce8df0b1bcd142", x"04a15d8054c49151", x"028c0b1d453c096f", x"4312fb0b00659d23", x"47b3ceafe3c747e1");
            when 10727022 => data <= (x"05bf5a55f8aba32e", x"25e3ed84a5584cb6", x"3a6c0138e912ee4c", x"998fcf91959eebd2", x"a7704ea4067bf772", x"1fc5692230353a7c", x"02d355bcb70fefc7", x"8a125cec688062e2");
            when 29918865 => data <= (x"913821bf20768ae5", x"d7c0e25f3659ebc2", x"0b00cfaa197b1bf4", x"62530416fd98890b", x"eb34ca9120f9e8f3", x"f1712dab3b3b8aaa", x"4bc4a8a95386ee85", x"e05c416e3a8caa08");
            when 1768735 => data <= (x"558fb52662465b55", x"097b6a4151b6f7c4", x"007bc5d39b407ff7", x"ddafefb5382da1cb", x"cb3e26be6b3a64a8", x"0537dbbab9bb2ab4", x"1b85f36c7d408c5c", x"f9ef85ba9eebaf22");
            when 32513160 => data <= (x"ea9eb4133eced684", x"e7a307ac2fd42aba", x"e256a177f80c88b6", x"83dae35880782267", x"06a9828da25f16e5", x"18c74f7faaa95c68", x"18f23fb555ee846c", x"b3558cb5cbf8877c");
            when 4115487 => data <= (x"2408ae246184dad7", x"815e8a5290c107c0", x"b4ba2b5e821864ee", x"1d04dbfab1404a96", x"77ee9987c2200bf2", x"95c57dc925be86ac", x"e8b19c6379baebb6", x"72ef479ffac54a8f");
            when 14497320 => data <= (x"7955d080687dc17a", x"9223d95fc5d29fba", x"45d55c4aa2b67acb", x"8393a65628148f21", x"312094618a4e205b", x"c7453dee722702be", x"61301e1fff5551ff", x"1856c275b676b2fc");
            when 19536410 => data <= (x"058e54c8093deba5", x"69731dc605f76804", x"1c60924059529d42", x"ac5e8be6934a1a9d", x"14225015a32f830e", x"a1cf597972decf53", x"4ca4e5d51bb12cd3", x"1bc9deddb1f8e8d4");
            when 7820290 => data <= (x"8bcf43309e0059ce", x"96012f470eaeee6b", x"642aad7f24160957", x"1e22b8a87de3b945", x"0cbb14dadfff202d", x"465b52a87f1a97b7", x"cd65703ebd98062c", x"8b39ccdba23dd1fc");
            when 9016150 => data <= (x"de69a5a67e10fccd", x"315a0d653d7cb5d6", x"4038e04cf54f454f", x"7d5ecfa009916ac1", x"887ef3b06a56192b", x"95be9e49089524be", x"c4db142dee7e0aa5", x"0f9b985d27dd24ae");
            when 30218703 => data <= (x"88e9a01960403466", x"36c74721a4d01e69", x"abed236c68f98056", x"6a1e3f443dfb05e4", x"8c3d78d1cf9fa285", x"403172f28f6b6225", x"97c0486dcda11aff", x"3a61016f1b0954d4");
            when 2960034 => data <= (x"f0ea323db4953c75", x"44e61f0514a05474", x"0c68607191fccc5c", x"284f9a910715504f", x"562e0b0c6df396e3", x"b56c1f9b71d629bb", x"06fc9e6485a91b96", x"56994f6cfe050405");
            when 28217342 => data <= (x"8b8d65085961b63f", x"31f6054b4bd564fa", x"7be231775750d978", x"11ee6cfa6c1a4a29", x"b91a6be44ca34ce0", x"120e5175d3fe2d75", x"643d7356fc540c47", x"c08bf7429916f8f1");
            when 28184442 => data <= (x"ef92d1624797cb5b", x"ff2d89ee59f1bc8b", x"a603cf3fa90eefc0", x"2de6839552bc0e9a", x"72150844ec02bd5a", x"a7dbd47d929a8ecf", x"c39f2d421969473a", x"fdf306d625e1d941");
            when 18234699 => data <= (x"36fa3ea386ebb792", x"19992b6d3b9bbc9a", x"aebba3256aead2f7", x"43bcfdec264462ee", x"6390c7bcc137a562", x"7ae1045933f829d1", x"c1e0fa47666b952f", x"59c05965c0778b7f");
            when 23231019 => data <= (x"5b5d4693bbb6d4e2", x"628db41deec56f5d", x"0541fbe2e61126d1", x"1a0ef5f3870949f3", x"49b278c95be1fb19", x"b5b302b6c5bad1f2", x"53945170e6c2a0fb", x"37e7e11c1e4aad9e");
            when 30428052 => data <= (x"ccac9779ea7d9c21", x"80b7f1ea50aca2cf", x"6a949e1f89a0b553", x"531bdb2290cddff7", x"0c9635fda6edf534", x"7dea857096b477e3", x"67e47b5b47fbcd08", x"5d403981cecdb872");
            when 8435984 => data <= (x"529df78be18bf3e8", x"9a5b85aae315cce7", x"151dfb0d539d2f24", x"ec36394407771501", x"94a9415f04544a15", x"829ad8e6bb00eb25", x"c26e44ed9f4105e9", x"996577510296c9c3");
            when 8396263 => data <= (x"5600b3737546774b", x"4256cdaceb078570", x"6f08de2efeb8e579", x"d6b6a354617808b6", x"b2bc25f4122964ef", x"fa1bb03f7db78a17", x"5d011d870559f553", x"ad07d0b72b7540b6");
            when 1482604 => data <= (x"d70212e9764f5ee3", x"cce5257fb0b0b434", x"36d485bdceb0fc3f", x"af307f1c8380fce8", x"11ec583b6cc78fcd", x"e462a41a96e902ad", x"1e878b3b43ca71ec", x"295ead41252d686a");
            when 22542970 => data <= (x"4ea30898a02012b5", x"f0152cd22840b011", x"350726f73cf2a5db", x"1b93968147a8b120", x"7f52018eea8c9823", x"89299a1d4c9e18a6", x"6a94032604ea8bed", x"b5b164c87214ad7d");
            when 28702410 => data <= (x"90248779da43cb89", x"0bde53a449483f2b", x"babb5ab91f5aab7b", x"e07856d17ff35952", x"5cfa6023baee1dc5", x"72ae577465b3b93b", x"aef132d7f1aafeaa", x"b3b0f9d571904908");
            when 18328506 => data <= (x"0aeb70e1fab88b54", x"4ce4ad575e9044a5", x"9b8e7c516ef55102", x"b7e230c3a1bfc186", x"9822dcf1dbe97226", x"e5c6e4dd7c7fdd4b", x"18d0a2118daad5a6", x"cfd53ff6c30daf75");
            when 4576549 => data <= (x"030949c9e6ba87d6", x"c3157e23c38f3378", x"6a274a553894cd62", x"02c485ce4d64192d", x"15a2874efa61de42", x"1a03a87babf8a17f", x"84384d8762ba8f60", x"f1d1bcfbd71a4966");
            when 16986597 => data <= (x"95a611616862bebc", x"a64393f8bcc02e7f", x"adb5f4f026e51146", x"ff503149b39dc2de", x"e70ace408c738f58", x"ea6c166ccbc88582", x"f9a399dc42813123", x"cf1df9e6d266c014");
            when 32822836 => data <= (x"3d7097408bce095c", x"3c9c9217959ff8ee", x"ffc48300b8381dc4", x"1dd2d92bf2b1286d", x"88633fbcdd179210", x"00b0b6a5534055d2", x"d637f4e29d28f0b9", x"2c674b3be9833e1d");
            when 7325045 => data <= (x"9717787aaa18a53f", x"fcaade104dd0d890", x"32353e2f7240e0ea", x"bfa01015b8fcffac", x"b8b4eedaf64cd306", x"6b8dad0c4d9eba28", x"65974ad448a81906", x"0227d8464c912395");
            when 32962126 => data <= (x"7bcb380c772a3a0c", x"0e5c3ba879a67c3f", x"9877183de3655862", x"ee17ee885d41f22f", x"649b6e9fa9b1f5f8", x"1ee467c0db58779c", x"d22a4b48416658ce", x"991f090347e678d8");
            when 21913700 => data <= (x"6e7ea1b7441b142d", x"7e2c80e156d0aa45", x"ea26a869ba57c6ba", x"c4252d29d7cc5b83", x"192e7f68c912f03f", x"a34b2b8e5c919de7", x"15dd5f050c2ac092", x"5171ac402c66cb74");
            when 5590428 => data <= (x"61af1346f34e28e6", x"b12d043c8e29b3a9", x"ab6959f3fee98904", x"88ce8aad8d9748f1", x"5be6f3c2c089b276", x"48be8c2938906781", x"1b8bb912075f8391", x"86ab293c49963996");
            when 28969027 => data <= (x"8bcaba0be9c42701", x"99874d9f09f25c48", x"385033ab335b6ee8", x"19c8cd4d3efc159b", x"37889bd98b5bda13", x"99757aa7639444ab", x"91573ecb832ba531", x"21ce6d6531eb218d");
            when 23737443 => data <= (x"19b643f8c1cec41c", x"99d6cdf83f23b930", x"0a2581bfe29d169f", x"818c4fcf0b1200c3", x"80b3304ec1633a94", x"bf639e584434d0aa", x"ecf092dbea4ab015", x"89956aed43d72ea8");
            when 30058965 => data <= (x"e24ddc6bddeff0a8", x"64441441a15f63bd", x"6089ae1f267d622c", x"cdeee6f46d975d95", x"c93d350f7ec6b23c", x"a9ffd615a072e09a", x"4962bd5d9b54f08b", x"78e160ec097f987f");
            when 16375362 => data <= (x"e587ee4b172d5798", x"6d2743b326a331be", x"35f1f0b1df170308", x"b97df57aae7f69c2", x"74d05d0384e143a7", x"31ec9eedbdf76f01", x"fbe12258a7c17d89", x"6744d1f8e7f0af6b");
            when 4770371 => data <= (x"f70db544a39c3449", x"240a6e6281dc3c39", x"ac748ebf9a4808b8", x"e254fbc85810036e", x"772a5c5904d5a218", x"d832e813c9acd50c", x"951b402b2626a0f5", x"e96350150e004623");
            when 24728583 => data <= (x"22a9305025f26aa0", x"8fcda98de2228390", x"9dd60635c982747a", x"8e4296e7dec9f9ea", x"0e4d5d901765a293", x"fd37d3b586a837c6", x"0c70104caec2dc86", x"c60a2ca10d68e566");
            when 1283603 => data <= (x"be09e6ec4749027a", x"b91deab762c7e13a", x"ff00a334363eda0c", x"7a07984dc82bf5d5", x"c6e45a10d9e8f61b", x"8abe8882c6c7c0f7", x"de3be80ba321d281", x"5fb244538387f91c");
            when 10573423 => data <= (x"0b15bbe576b12bc3", x"6772cc77c357a487", x"4a1159e8e057e558", x"a41ceddf69df05d8", x"531b094303090384", x"d20bc5210de1f709", x"8cb93e091b6bc590", x"499ed5f153c2fc7e");
            when 30377540 => data <= (x"e9631d2bd44c106a", x"e733eb8389926718", x"133561522166d3dc", x"4f79f59f91f39e98", x"da6e071adb41d68f", x"4c66a00357305d61", x"881aa2ea963e1dbd", x"1f74162d87ec4da7");
            when 16751949 => data <= (x"d65b512eb4fed61c", x"0215113ece2f8270", x"f605f17b0d945a05", x"89c3e346e5c9551f", x"faef4d3c2f645857", x"713fe8236febb8ed", x"612982d60303ad89", x"8fdf86e543bdfb10");
            when 12965783 => data <= (x"e5f7a3b9d151db19", x"f863f16ecef00093", x"4a7c1dee67da16fe", x"04ba321e7d811a1a", x"f2225440b2af4822", x"32ee217a3c73dc37", x"ec09cef8f314fcf1", x"ef11685a8c35eecb");
            when 26380361 => data <= (x"edcd8fb4b6b62645", x"053294fc9dc71ff3", x"ef459409460a73b9", x"35a87267d7c3d30b", x"d8939253c255567f", x"f589e1a5a7538f1d", x"ec53df2778216f5f", x"8852d6e34d923da3");
            when 16526528 => data <= (x"cb093fb0d014ddb8", x"e35e0b30acdb582d", x"016e014fa2a2195c", x"852a1e158561713b", x"e556036865b5b418", x"b8f77db8de38309b", x"cbbe877a90a856ae", x"3ca8c796d609413c");
            when 30116933 => data <= (x"7973facb5da8d41b", x"7c255d870c2aff58", x"70122c0b760a703c", x"20a0fa417a6ad466", x"2636b59cf6c1594a", x"6b22bfca9eeb9ede", x"7c82a260f556c04a", x"cc9af6bf02a583e5");
            when 14016970 => data <= (x"73c97317a540f2de", x"cf5bc6b64abaefa3", x"b554f9b65d53bdcb", x"a1662ef3b05da2ad", x"10052c79d73a2717", x"0e6bec3fdb79ce3a", x"67553e21e54daee4", x"e3408bbf037e19ee");
            when 23904564 => data <= (x"d7d0da2bf7901b53", x"73a3ff0211f5fcf1", x"bdbb0a02da8cbaa7", x"8b497ad54dfc0f09", x"6b9c18738149fad8", x"28c2be141ef13aac", x"c94852a4fb6d6949", x"4969779ba2be328c");
            when 19582533 => data <= (x"532549a19a3da979", x"4e50d86feb302886", x"6a5e8186609d9341", x"7638c5181d440861", x"8f0021cbb7b03ffd", x"89976f77c38737a4", x"b36e5e73048eacf0", x"2851467a4ee3c041");
            when 32602047 => data <= (x"12795bdf26988b10", x"d3586596ed5bbf91", x"f38c9e0b9d6e5def", x"6717bfb3500ca787", x"382a150214387e1e", x"40c98c0f9efa80c4", x"b6067beae21adaa1", x"f94c87de9886918d");
            when 14669351 => data <= (x"a2fce5645d537f19", x"787049e4a635bc9c", x"1e7325a8af96be62", x"4498d79b4f58e732", x"32564b353432389f", x"c91175f94ede2333", x"f0ad5b1ecbc2b24e", x"591ef83abb425a8b");
            when 24327407 => data <= (x"e18d823be268dc9c", x"653d0a04a846b4a0", x"d2e6fb5ffc9c99b7", x"bd5f0577a001ddb2", x"6a8ec6db6fc0c7ca", x"311759e3bc4446b9", x"e2bb62055a42b174", x"d526cc0c2074fc93");
            when 27131407 => data <= (x"21a9063e356f15bc", x"ab169f792fbd9d53", x"60d943b29f2047ba", x"e5ef5a2b762266ed", x"3deaf44137718638", x"3147f486e6a44ad9", x"9802f9067b416036", x"bf43862e551480dd");
            when 12157549 => data <= (x"711f0ba5a969c00f", x"156aa4bb7e840494", x"905f3a11c2256e3a", x"f3249073589958bb", x"7d22ee8ef0ef63bf", x"6d64aeb56848084c", x"936dae78222480e6", x"9cf918d06ba61a9d");
            when 13535388 => data <= (x"d28e05cf3f41899c", x"86e55d1def1e3b04", x"6082271f77e1e74d", x"b71ceac257afecc5", x"ff81872d4407e2d5", x"f1140985bf87521a", x"96cce4918bcd539c", x"1a6e207a2b5f4832");
            when 8496426 => data <= (x"7265aac92425078d", x"5bdd758919253564", x"48f3f3a3bd759347", x"9d78fccb5e6c9583", x"f7f64b1f6e6ca0a9", x"603db4696ef41d06", x"0e8910161928efcb", x"404697c45c09d8ee");
            when 26490426 => data <= (x"90ef54fc051520ef", x"1c52b49c1cea51c1", x"abc95646f61df5ff", x"bc95b07345723f47", x"fb382d503b312ec8", x"5a952e989ed85e58", x"73639dbf2192e44c", x"6898bb4db96ce3c1");
            when 4785381 => data <= (x"a0b4bb22ce237147", x"111ac2c28104dca2", x"5fa322109aa03638", x"88f26d4f6b0a88f9", x"56a5d74cc08050b3", x"7dec69f7a73f8c01", x"8f7850005ade725b", x"686edfa070b5ba51");
            when 21784541 => data <= (x"62073c5596f5ad82", x"301df17044a93601", x"af372c77418f2113", x"cbc7b8799a0afac5", x"8e7b1ac2ebcabc80", x"a55509f525fb9e3a", x"3e88c497590cb058", x"64e807fd77cc7b76");
            when 6153197 => data <= (x"77c1694572f90deb", x"e77d56177c25c8b0", x"612adcef7ec43c9f", x"5139beeab476a73f", x"0226c276c16d5c9b", x"79e635ed2ac4409e", x"0d225259492e6567", x"cc983331907a5ac3");
            when 5597080 => data <= (x"edfe491935340d82", x"0cfb1424e4c44e24", x"cd1e276c87b43ae6", x"9e03adffa731e8a9", x"2306a265b030d5aa", x"49874d1e85af98e9", x"41dbf7e246d75b10", x"09d4acb62cc490b4");
            when 33014947 => data <= (x"f0477036b84ee406", x"ab35abc76dc6ffe0", x"6119269e45dd7b09", x"d61521264386b65d", x"18d3197e78805ab1", x"b06c5868476b9fb1", x"6dc9c91c2bcdc1e4", x"fc67cadb657c3d4b");
            when 11716738 => data <= (x"0221bc12cf09fa0a", x"2d64ebf9f78d3726", x"3647fdc7e3555aa1", x"28f82cfea8512463", x"25ec1d498faa8907", x"d1717bbd97015c15", x"652ced110cfadcef", x"06fdeb9861f812a0");
            when 4755355 => data <= (x"c076ec1ed55931b0", x"e16de05d734592ec", x"9ac5a422b06d4e4d", x"4e8967e5c73a91f1", x"e2c7dc7df1e4f018", x"fb706ad01cb86f72", x"f092851f7b008c45", x"b381826ec60dafd4");
            when 27888581 => data <= (x"0777a9c161e269d6", x"83e4932551981457", x"cc8375f10325497a", x"87d65d8cb5845336", x"7c6fcdd288813ff1", x"f9095c6340dee53b", x"7573f446de19340a", x"06892c086126134d");
            when 20398412 => data <= (x"54b991400b988ecb", x"1a4d602136121fac", x"5f0e7f58d9284afa", x"4595c41971922b3f", x"051e029ff785e6cf", x"ba545b0972fbfc30", x"e804a64b7f13a4bc", x"a068b8ce5f20868d");
            when 16631487 => data <= (x"e9676c1f4bb1ad39", x"9c5409d173b5c36f", x"60850a0cf7b3efbc", x"b2a527fbee3c81a4", x"53d505158b19431f", x"13c56e3a680e7ea7", x"30f5ad7101876a51", x"9284dbe3c778b660");
            when 622529 => data <= (x"c835234696908f7d", x"44f0d00819497619", x"20a9aeaf6e956a23", x"3292c6256c3219a1", x"47aa4d56913cafba", x"364d37e12c4a1d44", x"6eea810085b0e4ff", x"8e109016f5b8d585");
            when 1375241 => data <= (x"4752d409a155ade1", x"f6855c0edebeb124", x"f032bfb54bd38bdf", x"060645c228de4aab", x"99f4d3983dfaaabe", x"6e04436fdaf9b9e8", x"58a7de05163c5a85", x"1a2438653911aa74");
            when 30253481 => data <= (x"b2bc57908dda6ce9", x"f9b5efa40f3991f6", x"b4a1f169bc34a27c", x"23f99c49454b86ea", x"6e6d26f3bd6f2db2", x"4ed31520129f8aa1", x"40065f97bf34facd", x"cd718c951efbceb6");
            when 6127169 => data <= (x"e9fdfa74a146cc29", x"fe99f39004b4d115", x"00f915f38d41e016", x"34337e435530338c", x"6ba548c0d08ec86c", x"9c133060ac8c652b", x"dc7c5d0bde2638f4", x"b49260701bebabf8");
            when 2809515 => data <= (x"97d6987651c02626", x"68701e71a0366332", x"dfe1293b2e86dad7", x"b9bdfb469a2aff58", x"8fb5f0a16e10b429", x"21e0d3b7b8e9e1ee", x"22247d964561b63b", x"c3feac594ff6e834");
            when 8998448 => data <= (x"96bf390e5b559a5e", x"950453c2df63f943", x"35846197dce5983f", x"18cb9d07308c8bb9", x"94ae02ca3818de31", x"e4728cd001cab1dc", x"632cabe9ec44c997", x"bec53f8e198ce5ba");
            when 31537984 => data <= (x"bc1aaf9ccf587092", x"55c1cd55e5c4d268", x"ee8cd7ebeebf8e61", x"8dc0a440b554daf1", x"dd38ade6c4ba3720", x"e26dcc2a0272ca39", x"52d3fafd3b6708d4", x"10b425b4c834d025");
            when 18167953 => data <= (x"c8a84c0c47e514af", x"633ba2e6202438e2", x"e380ea3f15935825", x"a1bc4d0f2ff20b52", x"81420b347d8c474b", x"7295b66c7396756b", x"f2b1149e532711c9", x"5dde093ad45d954e");
            when 7222559 => data <= (x"0cbeb7508128f7c7", x"091c87b466d3c8fe", x"0efde17ed64288a2", x"8e64b11541895f59", x"96c7efcac9562b95", x"f642f60819cf49b8", x"54e484fe53d88d30", x"5fd68449ee4b1b59");
            when 11116107 => data <= (x"e638804eff033403", x"d9e7776293fb8303", x"d23057417edfa7f4", x"b090577baea1d031", x"fb3ed135508399bf", x"2be9e660450fda09", x"e5a53f6a96f940f0", x"a39d1f2fdfef6dc9");
            when 7463236 => data <= (x"085f2cd2a41a1523", x"f04c430fdeec8006", x"7a1d4dcc70349f2e", x"66405f03f61d203b", x"b9b09a1b4ed62be3", x"da15fd01c69de97b", x"4c223fdd87370773", x"4b2045b1cbebcf84");
            when 17991744 => data <= (x"b4aef9c69e80cfa7", x"93eb91d4a4efff67", x"063de3206cf2d605", x"fcdb61e230aefb18", x"773ba1546d1b01fe", x"5342b97c45ce3a59", x"360ceadd418b7189", x"48aeb4c054223393");
            when 6796940 => data <= (x"4106c7a93275a9c0", x"a0725651ef9c749c", x"2bf4f4d39dca7e30", x"640c10c56a02fa5f", x"4e963f270f5fa69c", x"a1601bd98b6456bb", x"dfe02f0cae2a1f72", x"e1fb584272fc6e67");
            when 11058616 => data <= (x"5f6a55a88f942ee2", x"2b3a46796aa1298d", x"2468548fd973b026", x"33ab8df8613026b3", x"f343344535578b61", x"a99c6508c013805f", x"407d18ddb6e0a8c7", x"6f08b03978869f27");
            when 4679554 => data <= (x"d5a2b744e9d624d1", x"cb1f2a9cd074a206", x"714d20c4dafcc1f4", x"2f33b1cbdae84a78", x"5f1c8e1eaffc74ed", x"c2c19bf85486db85", x"3202dd041d7e3e15", x"b8f774c6ca5f8d19");
            when 31299640 => data <= (x"6ca9e9c6f534779d", x"2cf5758b35bd76cc", x"6f85d8c4cc63e335", x"86f8f0fbf01d6683", x"d9691413fe3d4227", x"6c018dd42ce923d6", x"874aa8890c87b8d1", x"f8ff027ef5ac99f6");
            when 22993962 => data <= (x"a15d02073a998ad9", x"39f98cafcf02c1a0", x"9a9322c879ae2e10", x"dd824c86750a722e", x"c1b8204ad04f6e4a", x"fd7a9d2b08113975", x"54f97e3ba2f31ae2", x"72c00cbe800d5d97");
            when 30417244 => data <= (x"39da3af7879485e3", x"5993e092323beb75", x"914f1198bba4978f", x"a33c2598bbf489b2", x"c38ace418451a39f", x"bfba805f16ed6b31", x"5a0f863b7882ba6d", x"ebac804f0edf2e5e");
            when 23018539 => data <= (x"516134e38e6f1331", x"aa3e90f7faebcc87", x"21bb458d6de62045", x"049b0315b5fdbf51", x"a5994e91595eb0bd", x"0ae72c40487c24c1", x"c0cd5e1e99d4a99f", x"8376c30e0a8adbb8");
            when 5017221 => data <= (x"bf8ca62e879823d6", x"9056bd32d5ccec26", x"ae80ae9d22f4da2f", x"0de43cbc82a38c46", x"4061fcd1b83f9f9a", x"8ff4efa0048fd510", x"7819bb58dae8f419", x"6b2a397597605cdb");
            when 25831935 => data <= (x"c816f23738dd50e6", x"6f1fe9a230254378", x"7a007bd3bbd6181b", x"b5633af2d33ef3c3", x"43c1ade9767a25b8", x"b43d7d4b80efbb13", x"71abc638145cd0c3", x"d2c9b1378a243fa8");
            when 24370763 => data <= (x"518f082460e5f9f2", x"42726021aa04310c", x"ad926596ae5c979d", x"73441b95ee3526fb", x"dbd096aa2adc8f22", x"a2ed15ca9689c0ee", x"ba193d150d8ab530", x"8dfbcd4c322fa74b");
            when 26746293 => data <= (x"9c9454c4d0cbd666", x"5596085cf4bd59e7", x"5ed00531eac63b03", x"260c9b4a7650b9fd", x"f3c374d81539ab3b", x"13b0b3d5bc83ad6c", x"c76876b498ec10ea", x"7e0967f8e84b05f3");
            when 32491340 => data <= (x"6955a9310b08fb43", x"ea9ae3fb2b90aa2e", x"917f5e5718f832da", x"c4f6c5dea3ec7b8e", x"37d997e384c9eb09", x"de4bb8b374bfdb42", x"bb9227c69834d1d2", x"0362e4e143868e5c");
            when 33222118 => data <= (x"f22436e62565a6a4", x"f29889743cc04b00", x"09f15d36ba83ced6", x"4594fdaf3b229462", x"2d0f8b9ac019eb7a", x"72b669f979969c75", x"5fa450c01168d030", x"391f62ae4081fa22");
            when 19022955 => data <= (x"2fb206e2b6b7c1b2", x"292a21c6e69765cb", x"5b61c6fe9a674ed8", x"86c2689048678d4f", x"2e39163434621747", x"555583ca907570d9", x"c882176c5842757c", x"eef35f93b775ec73");
            when 13576012 => data <= (x"49e1e8008a54ea42", x"c45a1000c4c3eefa", x"693563a58ea7e5ef", x"d2c4cff650891c72", x"46b1695143c253aa", x"3acbea2e87737e8a", x"4c39a95676cb4d53", x"54024ff7a778ff02");
            when 4299810 => data <= (x"92ae1ea119e2b0a4", x"e81dbdb1e7a3b9e6", x"5beecaa7ed3e008d", x"14bfcfc92d5c4023", x"18cade7b2f718612", x"8b7a4b9afb2ad7da", x"fcbe9931729164ba", x"c3b9be454b9dca73");
            when 10900786 => data <= (x"3c47d3658826607b", x"64cd3321d43e16b2", x"53af4965629cba85", x"78320b69a9cfcd6c", x"a36ce1e81544724b", x"b86f163b84018900", x"3e2a95673c8cc636", x"f89f7224baa283a9");
            when 1510652 => data <= (x"2336aa250e6b6957", x"28f4100a3f204a2e", x"6088443aa64a05a6", x"719ae30865fb2f1d", x"013f5e9f8cc33981", x"bafaf1736ff7f793", x"ffd98474044a2f48", x"5c0b0a7c63a306b7");
            when 5879251 => data <= (x"df9fcdb7ac4b3afb", x"28650deec1160832", x"959afe6605710449", x"6f3cc4ec29d82c33", x"8599dc36e68f2410", x"52f67ed579995dd5", x"aaeb8eab9218549c", x"f019bec876651c8a");
            when 30456581 => data <= (x"cdb8ff04a9510c75", x"2f18f281414e7153", x"2047d826f41bd5b8", x"744e422f2686114f", x"cd4450f5b78423c4", x"0f430939eab8c19b", x"9d125421e9506d10", x"3bd33ec609dc8d06");
            when 909452 => data <= (x"300c3969e20b5c9f", x"f2f13dda5e569721", x"6c653d0a73d31f80", x"612d5c90b497d9c8", x"2cd1f7fd2c251368", x"364105fa4a6ba8b7", x"1de14e7493689c8d", x"07e6f4535ef30b52");
            when 3903904 => data <= (x"151630a08de3caff", x"be0b8ac86fa3e157", x"cc89e1617a5e6c7d", x"0c3cf774787173e4", x"7d8955f79ce9a046", x"064f18e3214ff609", x"87c19c93fc211505", x"942213c27a9b2338");
            when 2902108 => data <= (x"315f73ffc8272bad", x"bd4e178520f6088d", x"196c350a2831add8", x"97bcde1a454c68fd", x"ba5754e4fa80766a", x"53a8ba7d03cef534", x"a778a8311b11948c", x"3dd485d0b5982bf7");
            when 32936242 => data <= (x"96c3b1a6bc45ef89", x"920e8eb000b54e5d", x"36c0e3085b15010e", x"9b870170b2c52a38", x"732a88519bc3da1e", x"1fcfc1ac26960365", x"c83ad1aac8a939b7", x"04d95b8ca2fb100f");
            when 21192781 => data <= (x"c1c18d8def84801f", x"37b2bd228230c6fe", x"ace0445b664c149f", x"7796286278e2c5fe", x"b4eab364e06897c5", x"d501972508d88b65", x"289f81925e5b4279", x"2080cd3c644af264");
            when 29421994 => data <= (x"6df645165e619285", x"fb58db9831d2a3e8", x"ea885eba1ae99387", x"0abc5a4fd0c01657", x"29efb26abca5704b", x"8f8cb55260caa351", x"c9597cdfdd8ed4aa", x"60091b99dbba3e73");
            when 29746606 => data <= (x"c2fc76f2fefeb41f", x"d0f7ce82ddb332e6", x"a3d354b3cd614f01", x"09edd3a8b388837a", x"33d1a4076c8b77c0", x"d87a7c4672b94411", x"adfc2764d3a7680c", x"da9a838596caaa47");
            when 14615824 => data <= (x"d82737c64fbffe40", x"d89274fef2df718f", x"040db39a1173aef3", x"4958cae3bba568f3", x"28f4debf9f4f38c0", x"3b31cdf7ae01199e", x"8524a316c8005cbc", x"51c67878992d02ff");
            when 22388853 => data <= (x"a3c017c8f26c9a83", x"42c578c58c936e64", x"5a46864f7faa7040", x"dfa14738d4ae9aa9", x"df22ed70b066ce04", x"93991cff179edab9", x"946bca04c01f3218", x"5f8e05d452bac557");
            when 30449827 => data <= (x"e2b10251842940c4", x"f373e3a01b7b27f0", x"b913493c00b67409", x"9d2618ac2cdbae12", x"f9a28079a70d43c1", x"35eeeec6e3ffd64b", x"078f5786fc2d4767", x"f1f1bc8cc7979be0");
            when 16617823 => data <= (x"a395f702cd4a26e0", x"b47ab792177ee27e", x"abb7e2f970ec3371", x"c900d6c473ea4572", x"daacfe19ea6093a4", x"876cbbf62e372474", x"75867e40f0a0f073", x"5b04c59b913d92b9");
            when 30987280 => data <= (x"8257fb3d338203ca", x"1412462dbb5019df", x"2a8468a0c0fbb51b", x"1742bf33974d17b3", x"f251f70fdbcf4065", x"a8b738046ac0d9aa", x"ba5bdf2121872961", x"c7f8981b4bfe7428");
            when 32858779 => data <= (x"2a27023503ee1d75", x"32851cd782ac2810", x"f641a1a9ae39a4b1", x"5efd07f85de298c1", x"dd6cdf7f05b87ad4", x"1e8f323741fca3da", x"3cef2c0f7240e4c6", x"432c5d07dc433f5c");
            when 10701657 => data <= (x"388ce1a9ccf2513b", x"bc174f079c01cc5d", x"2851295a6fa3cb1a", x"cd346145f955a82c", x"f70434295b47d0a9", x"ab40c83667b83846", x"f977bed524969874", x"18d4132a550cb2e9");
            when 11191401 => data <= (x"5da57dbe0408c311", x"5c6e547e403f1ce9", x"948595b394554849", x"3618c279b4bf35d1", x"623d4c5b8b3f722f", x"d3a0240028b51396", x"940e64de369681c2", x"f8d147a4c0fde17c");
            when 1146334 => data <= (x"df8f80850639027b", x"22473a3fa2fbe279", x"5316432feccbd174", x"f9740c92338ab46d", x"a2cc861dd1978547", x"fccc881240e527eb", x"4b5c85f14f29a0ed", x"370eadd7deea9ff8");
            when 23844621 => data <= (x"178107b140e18d7e", x"c2a912212ec06cdb", x"c8036b7721e34b16", x"00f626c15cb3ddc8", x"7b4dde40756f0425", x"ca211c6571b4a794", x"eba546b11197d60f", x"9595ce3b320733a2");
            when 23456904 => data <= (x"c7fef21b07208d7a", x"57626a972af720b8", x"a09eb71f3610cd59", x"d3fa909e8a8a3a46", x"fb41666320ef277f", x"bd37eeed5896d044", x"b4c93f1dce741e6a", x"12182252555fc89b");
            when 3663632 => data <= (x"f13be8d82e74cf4c", x"86ddf6bf830bcfff", x"d98fefb340291c2a", x"44b930ab020e7a2b", x"edb8a024724aa8ce", x"67bef8360f86897a", x"13199d1d9ebb6181", x"68f0bbda7fa5616f");
            when 31351123 => data <= (x"b8d5133d4d1b6b8d", x"7f5c406acac67aed", x"6282dddb28259626", x"318e30f9dda7a3e9", x"7daa6d046f5b6b0d", x"ba49ba8c0bae9061", x"424db1d513d6cade", x"07a6ca7833f8cf3a");
            when 3159301 => data <= (x"9b7207ba48edbda4", x"a4bad70139ff16f6", x"5c4c1e552d94ab76", x"2546f4d2ec2977c0", x"5f1f59051f12a0c6", x"2abe424dee703254", x"6f522dcdc0e09193", x"47edfc9e19b66115");
            when 23124361 => data <= (x"ef8311d78e2117c2", x"88a3c65399cd0b23", x"822597736772f867", x"80c8dc7b3463f0c9", x"ce4e0d7d19d73700", x"7a6088fdf82e89b6", x"5d665a89dff836d2", x"eb8613a8cc43d6d5");
            when 4959360 => data <= (x"2cea6b4055248685", x"798ec05ac35ea1dc", x"58ceb8a354e954e0", x"624949ef3084973b", x"dfd7057dc49afe67", x"8458d986d6031d93", x"748a2449d53e486d", x"b76d6cee087ead31");
            when 11673894 => data <= (x"5eb7983d6387a310", x"e3077cc674a97758", x"02e0cd12ed2eb22d", x"0f27b0ea218f7fc6", x"6348e5a5b96fd08a", x"90041bea9f633a65", x"8ebb1699b0ab5379", x"1628aa0a9e963cbc");
            when 28013886 => data <= (x"c4f83b2ac065670e", x"e8f70432d299f07b", x"943e4c1a58a13567", x"bd58d25a66ac7c46", x"6c41b9773d2fe74e", x"9d353eefac71b62e", x"fd264db272cae46a", x"00957b7c71c55c3a");
            when 33233782 => data <= (x"9d2a1a3886f57fb1", x"dfa3cd0adda0e1b9", x"9d397dcdd35c2e5b", x"ce370b71b2f79423", x"bab1462234901256", x"1903a63eace5b602", x"4004903cdae8a4d6", x"1175a1bb8f4fe987");
            when 1238884 => data <= (x"f4015047762b4a20", x"c1171226068e327f", x"69506a47aade41ac", x"958c4a18fd8405ce", x"7131aa2c972d4260", x"ab8a872134bd98d7", x"77af31e80b1dc3db", x"84d552eeca8186ae");
            when 28454437 => data <= (x"bfd590ffa6889bb7", x"bd4c31bbcb7a5588", x"557d4af9abe7de1f", x"1e5b43d7dc015006", x"f5250434a0db0424", x"027f749bc5ed1f72", x"2afb07c71bc87e37", x"846fb90696913fe3");
            when 25822325 => data <= (x"ae61313ee7e8cc5f", x"a58a4a73535af560", x"043383d9aef4d1fe", x"372e27e9da399309", x"767121a8222c7b4d", x"3cf039dead8fd85c", x"b54ea78fc17d69ce", x"0cf1c30267f69ed3");
            when 13515280 => data <= (x"3dcf088681e217ae", x"b8ea37a8758ea08a", x"f72cc40ea69786d4", x"604d1c18df674d83", x"d679590045256b71", x"798962ed42465f8f", x"40cc8f6367b18430", x"fdbd6806b4105c28");
            when 5341276 => data <= (x"da5d70d220829e81", x"63213ef63b13b0f6", x"6a447271da323169", x"b5d3728e06161cce", x"a1cb1a5715e58732", x"450d8cf6f382995d", x"e5ada4929251c42f", x"d0aec100398b2d6a");
            when 12489198 => data <= (x"cc5a418f31c8dc59", x"d531b6735352f15c", x"902166b8b0dd5ee3", x"ef2c85bba202213d", x"eb16162b192b604b", x"9d1028793f4a50fd", x"c3197fee5cd08f16", x"b7a36a8df49fd23c");
            when 14037203 => data <= (x"0fd9efb7ee6b3bac", x"45eb99d81380a264", x"4984275c53df68b8", x"5cc43bd37a63b7c1", x"b6c7017320286e0c", x"7a0540d3b1bafe48", x"25ac3af8c8707347", x"51df61c7f6bc594e");
            when 2856808 => data <= (x"2ef8108e95cff67c", x"8d1dff7a5dcc63cb", x"1499a203fb953abb", x"6e6ecb26f8b2a272", x"6fea93f0309bc1af", x"61931d8ad5563ac4", x"dbccd9da1d4c3d64", x"640c4a6279a5489b");
            when 4048696 => data <= (x"5296dc9e24d97679", x"3af5bb0d675b40d1", x"289e62fc462cc9c7", x"8c25d9553cb54ba9", x"31213c5096a45e77", x"94aec5c51f425aee", x"db8c0a9899bec67b", x"df7fe3f6f85fb8d8");
            when 818943 => data <= (x"c173e9e3e5ea4c8d", x"37a00651594b5f40", x"2a9f6fd973e974bb", x"339c939e38423fb4", x"4c7e9df6721ef45b", x"d4c21baac5799118", x"77c996051e545876", x"93e5d1e946cac15b");
            when 13050244 => data <= (x"6efc2846ea7a0967", x"b3c7bb16540f552f", x"d1d7c15b6e0b180b", x"633168000c750e93", x"d9dfdeb335559eb6", x"61d344b30ad18512", x"4654699689bcccc5", x"167ca578399e7fbe");
            when 9826221 => data <= (x"17f6bd22c2b2d877", x"1c74572a1cd55fec", x"674a49e6752609d8", x"684409c8da06ab7f", x"a719d213ef31dfeb", x"0324ae09860dcdec", x"7ecd101cd811f025", x"0ddd69b99f98de6c");
            when 4689551 => data <= (x"d1599461f559b128", x"d0993e661cf9dc8d", x"2ed3c136f7f3f2fd", x"b8ea8acb46e92679", x"ef9af795d6d120a1", x"1b750c236450b48c", x"eab15373f9319db8", x"1b89b8dc3cbb3663");
            when 33760742 => data <= (x"b65a29838475332f", x"8efdcd6afbef8cbc", x"93372323aee728df", x"d27447fad4d37e61", x"959e17a8f637b564", x"1afaa9c654019158", x"ef830946b077c38c", x"01d0b8c70e51128d");
            when 9634856 => data <= (x"4232773dd5acf1df", x"2e5c598b75f1a9bb", x"2f72a3567bd0150d", x"75651e784d334b6a", x"70058091fa666c2a", x"c5db37a65a674679", x"481b871de81a1bfb", x"527e20db95ef5f4c");
            when 21318340 => data <= (x"a725b42b933e3cab", x"d91c2e222aa25274", x"22c5e0e2ff361739", x"af6a53b2f99dd029", x"6202a1d644533003", x"f16f35b3c1a27f01", x"7fbeb327a60b3b26", x"31f88e6e0497c8d2");
            when 15142854 => data <= (x"e1aa4f2e4a6f7b6e", x"0b706ef6cd91ebd3", x"cba7228b2926e00b", x"2c4e7cbadbfbe2ca", x"fa878c821dd8312c", x"7af46ef5100c37cc", x"e26dffcd8c9f26a1", x"cb4010f70af5ca8f");
            when 18585660 => data <= (x"7f072ffee321bc46", x"b0512cbfc102b303", x"5e853be953350c3d", x"8d378ae9717ef48e", x"8560fae211d9bcaa", x"58ec86e997f6039a", x"757dbc8b491211a0", x"cd740da340821ded");
            when 21237738 => data <= (x"79e37fcb948df3de", x"6ff09d53c9eb160e", x"140ea6ffdfa7edc9", x"09940425dc9372e9", x"131f03b32b36710a", x"9b258ee592903719", x"6d370f365b3bd17e", x"a6d4a08fb749ad90");
            when 30823958 => data <= (x"ce032877d1156eee", x"74814e4bb3256845", x"fed54d7255d244f9", x"7c637631b11a68c7", x"5a1083b1be14e30e", x"9b16aeb5ae1fe8c2", x"36dc75b4d4941e9e", x"6b79ea0dba8e446e");
            when 7076717 => data <= (x"f973dddd6ee80489", x"8f6b9a28c53c966b", x"7513f39de25e0bb8", x"229e252dcfd23dce", x"bc6d26676a4be815", x"6f4232f7cf0d8d47", x"a6b0b943c5d727f3", x"ec627c741c5b34cf");
            when 28574569 => data <= (x"261ff1afe58fa55b", x"ca4c91294dda5443", x"c833fb6772affa0c", x"7b6019dfb9985585", x"a615b1c2019e5858", x"8f69070f485ee532", x"71da39b24505d4b9", x"257479a2e686c9ec");
            when 27256415 => data <= (x"86c5a82a11ab508d", x"c11a5ec07cb10756", x"1efc384909f87658", x"f68ef88b5c8db689", x"f75782be69f43843", x"02dc55a26331055d", x"70fb4788dce0b549", x"8854f3952c4741d9");
            when 29653526 => data <= (x"cae0c3e20e3db7e1", x"2b0261993aeee79a", x"9c771c1eb9cb3ed2", x"1ed4350d1f31d716", x"4e395014387274bc", x"17c9102def7368c1", x"bd7b2da57330bb62", x"958b8d6289fbddd0");
            when 11988865 => data <= (x"0566ab87585c029b", x"973c752ca770fd02", x"f99220ebf630813f", x"b58542b9666609d0", x"5e1620fac6df04a4", x"c69655d000e405eb", x"308eb14c6e6e8226", x"496a6c1401dd3446");
            when 6920205 => data <= (x"cdb3cf45f8b3f6ee", x"bcca4f7b85f279e6", x"a9c7471cc2b192d5", x"16e6fa61fab25cf6", x"bdb34340620e5ae6", x"2983ea5ed199be6e", x"12395def8056b224", x"f21cce1aab02ab5b");
            when 3708358 => data <= (x"5b70056b3d5f1edb", x"64c2cff7bd8f84a2", x"2a7efbee009e2385", x"fbc793d245b07f3a", x"1f576f6a5c129eee", x"f12e09c0f0efe1fa", x"08f257d800d96c1e", x"c518cd3576bdda64");
            when 7332046 => data <= (x"7b2475cb033bdc67", x"758023403f4cc3e4", x"0f8c9b4de3538564", x"ed784d04afe40a6c", x"ad70fe5cfec7fbe5", x"ebd21e95d656e26a", x"25675b9e2bda6248", x"b479cfa802dd7bba");
            when 17716743 => data <= (x"901eccca3f92c18d", x"46555d231586d456", x"cebd97edcfacfd1f", x"feceec35b514d341", x"4cae24c16fbf8fa8", x"3a536f98d4fe6f72", x"536bdd6945202a05", x"fcdcf0bf67e9f0b0");
            when 31758435 => data <= (x"54907e3cc6fb658d", x"7ef11a62878eb82f", x"7e64bf4038774def", x"8a6a434398c040c8", x"4528e5b27a6e2230", x"a27462933ebbee1a", x"099eda68b369ed94", x"092c7ad98d2367e7");
            when 15984537 => data <= (x"faa29b7cd523ab37", x"338298a9681c31f8", x"51d22bd2a88607cb", x"96b06662107524d5", x"0513afe5a315ffb2", x"cfd8937d935ba143", x"df92ba66970f11c2", x"d816c0abe93e7400");
            when 11891480 => data <= (x"aaa8fcca18f5e317", x"239dae39961adee3", x"7478e05561abe96f", x"ad40822a3cba86b4", x"2de37e06768106eb", x"a7d53e41a8bd598c", x"592343a7268c9609", x"c80bfdb17c350972");
            when 4650989 => data <= (x"c3d10bd3d668a88b", x"b8116096fc8539d9", x"f0ab664cc06b2d00", x"ecdacc30c0cf4b15", x"3d3732326f8133cc", x"6d299ee9f062e078", x"3c7983344db6bb0c", x"0837cad3b356184d");
            when 17419897 => data <= (x"41e69bb2250e04d1", x"d447510b0c99f720", x"f8195ef02c5b3b1f", x"86f4e6706dd3bdb2", x"c5ee6e681cfec302", x"370468863f06b1d6", x"7a7939f5d72243ea", x"f3690a556c5884d5");
            when 18132891 => data <= (x"748efa73d8651c05", x"29a6588bb3c5e276", x"b495b106171bbc8d", x"38dae0ca8d09032d", x"7bc194cfa2a721a2", x"fbfce906c122d878", x"0e93adce23097421", x"2723c3f63634fdf9");
            when 25322883 => data <= (x"3c21cb52185eebfa", x"8faa18b58ed3d2ed", x"0b411509c10be00c", x"1d1de17a5f8314a5", x"fc6561e778fd851d", x"0b0749040f36dfcd", x"b1802197d2d15979", x"5221446702672b61");
            when 15265995 => data <= (x"235ab5777a9a536d", x"4c62bf94d88a7497", x"fa92a7002062377d", x"75dc534e36c8f7c1", x"850c450d0a106094", x"966bc051b8e905d9", x"6ee25ce4c4f434c2", x"a91bdc3dcde979c3");
            when 20859663 => data <= (x"c1e83ce34991abe8", x"ae95c1cd69c2f82a", x"11d2af718b16ec4a", x"413af52c2a516cc4", x"2ac1118f67b52500", x"36cfcd90fe4f6f03", x"8227f466eef9f231", x"d5ba33564364de05");
            when 28101307 => data <= (x"472a94aec75cc1e6", x"f4ad7864c7526c5d", x"3828a331e5a9415f", x"e6eee883dc0bdbb1", x"54901d13b79baa66", x"9bc4b486716146b8", x"f3c53da0b59445a6", x"1c38356e50a79f41");
            when 30173719 => data <= (x"734771ef6b702b64", x"de7c9a8c360273aa", x"db1a08595c475096", x"81674371de44df29", x"0abb4cd4dfc6407f", x"dd429f4e7a620f6f", x"95c951b463829c76", x"556245fac9d69f63");
            when 31657094 => data <= (x"4a6a35138c36fb8d", x"22eaee80c48de83d", x"eb0756f66b4e6083", x"df8d5d9c5ca045dd", x"a6ba853c4770d645", x"fc6adf45ee9f5f1c", x"a86791cbd7af8856", x"2a27cd4fedff97e5");
            when 22831034 => data <= (x"7b8a78f922e6735c", x"0a7cea59dc5b96ba", x"aa600183f41fa813", x"c60f9f72de2277ff", x"17f02f64110ec8f2", x"812128f22e41052a", x"ad1fdc6dcabbb54e", x"41773d81a77b15da");
            when 13075666 => data <= (x"2a3353fb55307078", x"15c28021a4e11831", x"12b1c14df71afa02", x"bf21538e7acc13d7", x"43d4f6fe208be1ec", x"45a8726a3638fad2", x"634aeb3af19d280a", x"4656f9df68dc2e27");
            when 13913820 => data <= (x"297095dabe612549", x"ec77905b9a22de80", x"d7ea8c5126343ad8", x"f9e7fab954bb31f0", x"6fbd4018561178bd", x"fce01cf4ff8c143b", x"073a74109f03edeb", x"453ec6135aedfb78");
            when 857783 => data <= (x"a5579369a97a5373", x"46dbba7eac960ba1", x"b24c58b359813031", x"5f388ce5b4a975f8", x"fece208496859456", x"7f47ba4b49ca94c6", x"19f2cdaf00889e9c", x"1d2f228b1a7871d2");
            when 20285005 => data <= (x"aedb4ffa06c6629e", x"a82012da7e28ca21", x"b3f2c7e1c8db9697", x"28be57903d25bc8b", x"9ab5fa0f062a25e6", x"fdb376f4015d8828", x"57e565162eb8e8a8", x"482ee8578527b291");
            when 28548942 => data <= (x"29c1e9222fe7c4a9", x"378f3f15ca9affe2", x"94f4f9a4af147567", x"ae11943ffb2f098e", x"6a445f66248a6c0d", x"9bb273a701d44b78", x"0ceae6f4390e7161", x"0424c46e7b68489b");
            when 24730327 => data <= (x"45ebd1acfc79f677", x"feb77f6c5ca62ea1", x"14acc4f73f3a46b3", x"00c06db1ea608044", x"6dce16c2d77474a8", x"dbda14da3d29a52a", x"846916b8da08f334", x"e65bba460b640bd8");
            when 24355974 => data <= (x"ab668d800453094c", x"be44f3bd71e06c56", x"b521b1309915091a", x"d75f3b8ec92e71f4", x"2342608d13c05fd5", x"dddbb4337591150b", x"3fe8bf29537d561e", x"f6b55f51437c00fc");
            when 33732076 => data <= (x"631c726df3374002", x"0765db647a7256e0", x"0224e85bff886f86", x"54d93387fb86f663", x"4498770fe1225213", x"6acdfe4abfa44231", x"62149845ed5806be", x"d5a24f67ffd5c753");
            when 17970896 => data <= (x"1f15036c436b1196", x"678cfc8f2d3fff05", x"b97f39d788d39ea0", x"5a965690fe9bba45", x"be65e626722db368", x"a3b1c06e175216a4", x"e8d101730b9c0848", x"0b509dec499099df");
            when 18451395 => data <= (x"9329bec81a197c6f", x"3347c013788cd991", x"a01b41085f622ca0", x"c475046eb70eccb1", x"dce67186441a200b", x"d86d170fb7655bf5", x"735e77773822e70f", x"6b2e26c60907b45f");
            when 22632674 => data <= (x"4fc8079609358172", x"5efd5690f894ef83", x"39ba65c60a1b4543", x"7f2d33e7127c1005", x"33c0513ecb1b5b7c", x"abba40bc13cc41fb", x"a13e0744ef9b58e5", x"cfb51a58cfdbe0cd");
            when 15699381 => data <= (x"64afacae75870c37", x"c86533f71d6217a1", x"e6b4d24f0fac5a59", x"7dbb230889509de7", x"5b5a09f2a3348fb8", x"9b3151f4b6cfa767", x"893d02b987f5fa03", x"d824a07c7d0581e0");
            when 28689869 => data <= (x"ceffe0ca49a4b77e", x"8ca3797296b8d063", x"2842bdbbc7eb7f7f", x"d0a68a5b5365d82d", x"79c66cd1c87cc6d3", x"4eba3400dd0b9497", x"53d1fb5fa3e661e0", x"932c28ebdd2aba69");
            when 21575262 => data <= (x"685e179ca9435132", x"1f3cd5f247e37aff", x"1170cfc25b2db83c", x"d878501127389146", x"aaf92285f96bf962", x"8c961223888d48e7", x"6ce30f7f47c8e4ae", x"a5504b510ba183d4");
            when 16595399 => data <= (x"b7ed66f73dd610cd", x"7a467acbd20a26a1", x"66317f67c3e60dfc", x"8e31c9b3a89774e5", x"4402f5c374a0bcf6", x"130c0ab0fcf9c011", x"17d7da8b147ea852", x"f38e29b22ea67ca6");
            when 30716306 => data <= (x"f4ecda439b8b4cb7", x"c96844b4d1ae9255", x"4e67546527af857b", x"4c47338fa7e69135", x"544d69da7ff3ba4a", x"7e32034657e953b4", x"2945b20fcaee3231", x"91cd9d81b22699ee");
            when 17225281 => data <= (x"833c63681c79db81", x"f0b8c4d03a128237", x"8de05420c92c2b90", x"252071a2ae71f6e2", x"b0d87a970ea165a8", x"3d1eb5458a36ea29", x"73c1a2ea9d40509b", x"2457c945b19a7aa2");
            when 16913057 => data <= (x"58789c836ecf1868", x"220e5aaf5cd5b4ae", x"464753764a413928", x"a60b9eaf2a93f93f", x"5c30770d3472cb3e", x"a70d88bd3bb31f67", x"edff0961aaace794", x"c1548b45d10a1ece");
            when 19245974 => data <= (x"4644ccced0eb8a51", x"f3b6e25f3a4cf996", x"9b8523710e7a316b", x"ab44fd812fe2c920", x"ec735df5a35efe54", x"e286a076ba57fa4c", x"b96a41ba1497ad76", x"35a51d274166f0f0");
            when 11194987 => data <= (x"dd2fc77bcd13f12c", x"ab2f59d84d7af1df", x"47b0682a95ed45f1", x"8670d37625ba1851", x"0c39306dd704605a", x"c24e67a45aaf39db", x"176434638e14d365", x"828d9081fc7893a3");
            when 22423924 => data <= (x"f6ba3b7554f8f1ea", x"08a93a72ef3fc2e8", x"7d880145fa159ae7", x"8db298d2ce1ff44c", x"1becf86aa22da45b", x"ffd1cea0222fc12b", x"e5a4cf02e1d10b8c", x"d885e5030179f35e");
            when 12374147 => data <= (x"9edbc97217313e79", x"b8b22d3d46284356", x"cfbdd80d8045c8bb", x"0d6442bbbfac24cb", x"054b1eddd3558e1c", x"3f2508f4d8605a60", x"19cd7365f02dcb09", x"3a1ae2debe27b26a");
            when 32317774 => data <= (x"e7cd4b127d8bd5db", x"e560c0f0ee70cef3", x"4e0ca77553577886", x"363c73cb4bac1a6f", x"308a15d385f83170", x"3f9d0e1bf6f33871", x"1fecaaadfac7ad72", x"b8cb5fb2ca14e4e2");
            when 26553008 => data <= (x"c3b809e033ff989a", x"893c86d3a0be6d14", x"f9886a36b7525c56", x"fd9c5b076a467a23", x"665ae49b167f9840", x"ac140376f96fe94b", x"d3e38cbb8de50f9b", x"321fc7c0c202cb1b");
            when 24250485 => data <= (x"7213a491ebfe8aaf", x"2678c5b573ad743f", x"1b629efd767fe21d", x"c51848171cf5d7ac", x"acd65a2da604c6e7", x"75fb43654664d5e7", x"a023a37c357f2505", x"99d9b80289b656b3");
            when 6255792 => data <= (x"1a69323a74e8448a", x"e82baa0463a3b406", x"065dfc4d71c34f7b", x"c5ee8693990184f2", x"f3d4c8d183a60fbc", x"5d0886876c3e3005", x"bd4cb3f109a927e6", x"5cd5484993201fa5");
            when 18548817 => data <= (x"9a59b988c7c1765a", x"5b93dafbb614d094", x"030d20b7d3f7db0f", x"3292f75638fcd7fc", x"73ab49d62aa87630", x"7914f898c5992e11", x"255fc476cbcd5050", x"56d367fe53f2d2f2");
            when 4297132 => data <= (x"e2287f075209a73d", x"39d018bfda7456d1", x"b8e568fd2a6da605", x"804ae54c8d5edde9", x"ff2ae3fe0ea379a3", x"cdb2441aaa2e3f83", x"6394de63ca36f814", x"76c64aaeaaaae128");
            when 14289095 => data <= (x"b049d339eb0704b9", x"e581363d3229db93", x"42f4ebdafab0e48d", x"5ce913830a434eb1", x"84f32a1c6ce55d82", x"f06bf38e8b77db15", x"7ddf7eb9e00b065c", x"d88fd4aeacf8f73a");
            when 16721447 => data <= (x"723494ab640fc3a8", x"9f7e00e452daf8eb", x"fc7a22bb3fab2f52", x"79b5ef69f1793535", x"154938f4102f411f", x"27ecf19d78bd42a9", x"ba1abac7689bab36", x"793b1453f190d0a1");
            when 26313154 => data <= (x"45f844c02e573b17", x"6f913ca99f3629dd", x"1563306fa8932169", x"7af5f712343821e0", x"799a03c9fe87b857", x"7e9d70558403f707", x"11cc86a31a51cb03", x"fd092445d1c10448");
            when 13790855 => data <= (x"1c84b9daebe294af", x"8facad58e9fd77f0", x"aecab5dd7adc17a4", x"017dab91876c923d", x"d976c5f31204610d", x"5197ff1ae5bf62b5", x"0d2cf067aced19a9", x"c85d41196fc06ed9");
            when 18607505 => data <= (x"93474ee32aae3c97", x"762642cbe58d54ca", x"f755f412a2fa88ae", x"9a311923d2fc2830", x"d10f5767a5202dde", x"d22b3005336c6785", x"68a3459943cf6543", x"08dfe6ab058ef881");
            when 32817747 => data <= (x"dc7e289e09af9f87", x"818501eef85c7391", x"61f924aabfd97a75", x"eb044cdbc44efe24", x"91969c8a5b78d6c6", x"c85a551c3375fa92", x"42e52581bc35801f", x"cf50ab17f5e1c7a5");
            when 4358873 => data <= (x"9fb1ffeea6e45a6a", x"ea28a11836409100", x"cd39be0cb34262fa", x"bcee8ab89d6666ed", x"86ba8f3983ed3b64", x"b39b184367ee4f8e", x"8aad9ecdacdc6098", x"8ac73880ac68cb88");
            when 6794277 => data <= (x"0b2594714e137042", x"2b9c59562e2d818b", x"36ada812bf52ab3b", x"63a252c312d05514", x"7932f5955f0d009f", x"30a6351e920c49c5", x"297de9651ed854a1", x"6d8494044bff7f4c");
            when 20504897 => data <= (x"3c415afefaa88b6e", x"cd2c8429dd605745", x"79ec4b67953c75d2", x"a522395abfc247b9", x"977f1073727f652f", x"ed67dc7c57645367", x"244bd1e092e1e335", x"75e27f39ec738e00");
            when 17534787 => data <= (x"d90b7fa6ffc4496c", x"4af723c50d8e2206", x"bdcba2121c4b47c0", x"8f17f81f5c1c9fbe", x"5e482d30a6125024", x"66bafce0c3285f74", x"cc7fa12fac87c2eb", x"3445a2ed9e0e1b2f");
            when 5227516 => data <= (x"bfb6ffd481dc7325", x"4d1c16b8c1c9bc85", x"fd436eb7b381ae39", x"e3a543c2d98aafbf", x"93b3385024e37f1e", x"756a93a0c6ddcc4c", x"3ef99c017e6e902a", x"e05481faffa53dc9");
            when 25348284 => data <= (x"4a2a47cfb53f88e6", x"61f0f123e788241a", x"d1a4794d90bc6c3b", x"0ab26ebbfac06758", x"aca634d63dbe25cc", x"47800d5d27fb144f", x"8eeaf0c22b15cccb", x"8da8f6f2d21692d0");
            when 10632069 => data <= (x"4d234a9e0b206de5", x"19fe68241eb6451f", x"061eb2dab10bf2f8", x"b6d10c45cc35f9cf", x"66ab8d80dc9ee8a9", x"33a8360f281ccefc", x"be325eb2fceaf947", x"f42bb727a9070cb1");
            when 27094297 => data <= (x"bf0d73aef348e818", x"f459d9944105fe8a", x"e7ae0d9725525ddd", x"4612ac768f79264c", x"86e0037317bb354d", x"663f0677d3d6b6ce", x"96415cb11e04cf0a", x"6771234b1f80813c");
            when 11587211 => data <= (x"ddb036868ed18000", x"ed60c6717577301c", x"0c2b3f00fb4cc6d9", x"f1cab092052bdae3", x"a6848d2bf6824862", x"3c30bc00007643c6", x"e3c4eead782aa23d", x"6f4a2a7d2a818857");
            when 3531209 => data <= (x"073cbd9b63086b66", x"592ae3c4b2781e1c", x"a3863aa742edaf76", x"0976be75fe17c432", x"399f59ee26a425dc", x"f5586096c4ac1aba", x"052750c97cb7db64", x"2a6dae8235ed4dec");
            when 33435873 => data <= (x"7af9969f8d3911a2", x"7e24d7a57fc5ad5a", x"3190d269635e0ce2", x"b04c02c36f409d7e", x"147787c5f75e9de0", x"212025f0f141982c", x"7543ae1f5f26bb94", x"ad6f38c979f6f8e8");
            when 24740496 => data <= (x"c05756e1dad0b481", x"923374616dd0c09e", x"4f8cf18945a9e911", x"5d1d6469d0597ab1", x"e5baddc13e44c05c", x"38041bbd4c6fc254", x"67fa1657e97658ec", x"0e8ff850c8f588d0");
            when 14933246 => data <= (x"7d5b00c35703d246", x"584d4cfe8eedd53b", x"703757dc2b9d3181", x"61630caa464f9460", x"e44b8aaa5130ce32", x"8f6c882e8259f86c", x"3a665b11c4724c79", x"09e1258ae10d8899");
            when 9094875 => data <= (x"140cfd7b5543c141", x"a6fe8ba34b8ca489", x"9d96235614db4604", x"61aa35c09003bc65", x"36dcbc5e98a0d3f3", x"6d44ea8d9c512b06", x"79a52c2e4ac244d2", x"a45cc989e28e1218");
            when 26286621 => data <= (x"86e27e884f09ad91", x"4cf7a5f0a8cbe3ba", x"b19bedc6af283140", x"7d63e6699ec28262", x"3f6f1364025a6b95", x"529d02ddcbcc9a9b", x"e057cf585cf9b404", x"280b650d207faeb6");
            when 4813124 => data <= (x"f384068d56a7a767", x"2f3ea61ce1ede3cc", x"b2680a76a55a928c", x"13e97a76882c5d7c", x"aa362758df8de5a3", x"800897bfbd60288a", x"2373d6c2185c589e", x"6d997ca3c3a0822e");
            when 14057593 => data <= (x"57103e8d528d5fdf", x"d53c3e7f5e8bf5b4", x"b7ead713b6f15938", x"951ff3a1f2294e56", x"1457407d97e6f005", x"19a5605bbfadd89f", x"9a576ebbb2700368", x"1f97f929f7b6b652");
            when 8606021 => data <= (x"94dda7d644e4435d", x"78f35691c974cce1", x"25b424ffb408e4ac", x"cf018425cef789f1", x"c6aed133a183f2a8", x"750ee89c8d8ed8f5", x"e17ef53322774c40", x"6cdb6582389bb9d0");
            when 2128691 => data <= (x"80a15173bdd5d2e6", x"a3072dcbdc44412f", x"8fa2bc8ecb2f6657", x"a314188b3d5a8589", x"4c2391f7ac41699c", x"ff15d3c1e1f25b7c", x"e808299a7403d036", x"8287aa411b7c04d4");
            when 8971307 => data <= (x"58587749edf96438", x"0435917f0c8b21f0", x"de318fdc8f367168", x"1a0f2a80273c3ab6", x"3d2c72c5bfdfbb09", x"16a82890af89b780", x"82aa6755165a58bd", x"e2d240b1fdff43b0");
            when 25467408 => data <= (x"c1cdd6525d8d67f0", x"c20f77876391ed2b", x"cad040983d4c01b5", x"00bb4c5939a8415f", x"28c940b9056637e6", x"44ad3f3de39da12e", x"6981c548f52af886", x"5db8bf1fd21f84e9");
            when 2842127 => data <= (x"802203efb1782987", x"c4d3b25401842958", x"b82fe3acd8e4cf3f", x"92262c3e712cac2e", x"58bb333307b7f7cd", x"230e659c4217a9ab", x"384459b877c48a05", x"3c0021bde7c4cbc2");
            when 439366 => data <= (x"510024059a0315d1", x"7c12322a4f885a72", x"73a98c5e0577b3a9", x"1349f837e99597fb", x"37b01daf876c37c9", x"1f2ca1c38e1d0956", x"2f1c1b77a51a818a", x"9db3d47ce07dc12e");
            when 7943999 => data <= (x"60f4244b96193977", x"62a6c80e5729f22b", x"e0b51fb023a5f0d7", x"c95c2f0bd87a7f0d", x"67118a067a38c081", x"990fc66f93f0b6de", x"b6d93118c1a951f9", x"10c46d4a29a46364");
            when 2982795 => data <= (x"132d7169f7ec883f", x"d5e0c5ed1252b381", x"5a2a1bfe2b6a64ef", x"ca5da249a118c96c", x"0437a93f78e6c0da", x"107e5127e3acdaff", x"aa6f86a41d993805", x"17488ebb6c19b97a");
            when 28918777 => data <= (x"9eaeb2ce9d92ea62", x"4719bb6e70a8bd04", x"40cfee3f2a4453c3", x"2475a237ddca39f2", x"274d8a174d522315", x"e2f9a80715230cc2", x"eeaf28c2405161bb", x"c965e1c64ebf3333");
            when 18056667 => data <= (x"b029890e2ad1c670", x"5c062a9802f65bc0", x"47f4684a25b6c8dd", x"5722f0f0930ba82b", x"f4447b3e00801b3f", x"8938347a214d0869", x"35cf5021629dc27d", x"c93659aa3cf6eb98");
            when 19176626 => data <= (x"b9d722f295c92f19", x"0e6faa41dd5f8424", x"2075d657294fc4bb", x"5b0b094aa9ef2115", x"b96aace1128f76a7", x"1b5dcec90d564ef7", x"08912b35d0ddb4dd", x"7d4490afb0349e7f");
            when 13548292 => data <= (x"edf15cd7108daee6", x"cd10ded0f3257b8d", x"eb58c6dfd8d49a22", x"f96e3396a3f6a63e", x"bd65386bd16998b2", x"d48618f9f77b0bad", x"fab2b4e26fe91336", x"a8df695b6bf8b8d6");
            when 16089516 => data <= (x"4d8a767ab7d1e7a8", x"1e401ae48e9e4f63", x"4878e013369fcdac", x"97d88f8ce2003203", x"27ca0352b57ef2f6", x"831361decb16b438", x"e54ea78d4a3d55cc", x"a76a0cf785d15037");
            when 5096987 => data <= (x"5b5957c3fd0972f1", x"f13febf7947e5a43", x"531a38257bfda602", x"ede098b8a0587ea1", x"bf4c3df24363bf2d", x"39f54cf9c2ea69a5", x"cf922b06d28477ce", x"c4fcb0ee216da9e8");
            when 15471435 => data <= (x"06d0cdd747449b32", x"c172a77c725682ae", x"bf70b78871f46510", x"374d6af14c30c8c5", x"ccb4a92c5e3dcede", x"cc64bf7cf0451b1a", x"820b09006d0409bc", x"394b978eb3204f4d");
            when 26202262 => data <= (x"57f435314026f715", x"6d1bcf6167da27af", x"fcec6a53e141a10e", x"68a4b79a364d1654", x"8a55b5176109eb03", x"c39b268fbca73f36", x"dd449109e2f696e8", x"6ffcf0db43f89735");
            when 33673901 => data <= (x"ab3a1b2f68441e19", x"2d8035accb187348", x"3d8c3a60c4e64329", x"b41dd75e1c325aa7", x"e381e96c499897e7", x"d2128cd5dff7c879", x"48fa671e3015dd5e", x"8e4cce039a372196");
            when 28529131 => data <= (x"7ccc7d494fdd5149", x"e33003392769e340", x"74ca475585ed0b13", x"ea347e871527563b", x"d7b6c03c68748261", x"ed51081b23ed37a4", x"a28e1828dfc0d3fc", x"2b6cea7a9ef38ca5");
            when 2239210 => data <= (x"57fe44c336483a25", x"b7de4ca7c0a24196", x"08c0a540b39611d5", x"546ebf17b1969e99", x"2c97af735eb5e00c", x"94a03a676252242f", x"ea189cd9bbb8b577", x"cd9451f3a7349d1f");
            when 32866486 => data <= (x"7edd009ab9862dd4", x"02efd91195e637c6", x"3669a42e79dc78f4", x"99b064c2950cf1ee", x"898a3f3ab2e97cfb", x"9f166f0f06cf1731", x"010eb3164b3148bc", x"9a29abde597f5796");
            when 30844963 => data <= (x"6a3e3f338c9f14c4", x"c918072df456ba80", x"c262ee7386637803", x"10f989157c75976f", x"ca73083f0d7e6572", x"b32e0b3fe2beb758", x"c00de5a9e040ef28", x"f53ccc1d8b28c7b2");
            when 3186863 => data <= (x"cb83d335e1def65c", x"fbb0bfa355348a2c", x"78f5500e6adb177b", x"ba32125a0c808db4", x"9447c1d937062abb", x"7ab0c4c8bb6e6a51", x"402d3a52af2a957c", x"7c2c2453c2ca9f5d");
            when 23741203 => data <= (x"6eb1b63fc06073c7", x"6bbb57162c25c484", x"63312268391ebdf1", x"639b1d7c9b1b20c7", x"175c6de13d15c432", x"e5aff4a849246ebf", x"df50a79940188fb6", x"1c8e11ba0685eb5c");
            when 28966754 => data <= (x"a6ae6f7d62d211a9", x"fe9c3c5a58f078ca", x"ef90c8db9715d69d", x"61814055d3bfb46e", x"228ee328d8bb2a41", x"b691bced6ea4c426", x"9a1df5f0aa7daf7a", x"d1277772b44270ac");
            when 22346873 => data <= (x"99a4c4f747132897", x"b976d98ff8ed0cec", x"47929fda20e128ad", x"b00b8f271bbd40a0", x"b0c0e4e51648d379", x"e08075f3386e5df1", x"6c48614c11d5e2f0", x"110928cd9073992b");
            when 32498768 => data <= (x"4959e14a75600b69", x"ca1f48b9644d96b2", x"74be73233ec19d33", x"2f660e0e882bb1f7", x"60a39e17b70ddb90", x"1872f0da95d2f370", x"eff7ef4c1381004e", x"07b1a66df8fbc62c");
            when 4339052 => data <= (x"4ce63c3299cb7186", x"b6ce474187eabb91", x"0a6298d799d96e09", x"b1382132d8997ab3", x"878c2d1fe9dc1eca", x"9efe765b04f7e94f", x"e888bebc34273b7c", x"41b00f60884e19eb");
            when 27305431 => data <= (x"e5e19df51f6cb2fd", x"c4e6073189afa4fc", x"2d100622c18e7965", x"0363588f84e5eaa1", x"1d7694ad97510b1c", x"665520a0b5be578c", x"a395f0d60c91017d", x"40ac65f895e84912");
            when 31602269 => data <= (x"cd3f037ac93a28d4", x"9c22a396c68d2bf6", x"ea83a011b1c6104f", x"77a8e3299bfc0d78", x"65def1ff97012324", x"71d2d8a0a946ce1f", x"2fe45f13f788e2c3", x"255e36bdf49466ad");
            when 20873450 => data <= (x"83a035110f145b45", x"8de5b707eb04f626", x"6322ab5d261b41d7", x"92d137cfe4f34fc3", x"22a9958abe92bc5e", x"6165088f249364eb", x"b23cbe593102e136", x"17ec3ca65b7e4172");
            when 17784244 => data <= (x"c982157ac43e794f", x"5d2daa11d5cd06f2", x"dfdc3dbf0db59815", x"da5ef3d381b22cad", x"788726cad3be483e", x"e95309521c8d1828", x"715060d4e04937c6", x"e6445698f7bf619e");
            when 9657386 => data <= (x"e2f4764ec736414e", x"8ce7ece595a148b2", x"2daf4d5b6839cfc3", x"6aaf5ca009bdee5d", x"b3101a973bc75278", x"ce661d57ee7c320a", x"5934dff9c73e4f27", x"a82163cd171d83ed");
            when 7892042 => data <= (x"23584156fb5a4f74", x"f8e10fa1669d4dc4", x"282082854feba750", x"17b59bca5971812d", x"34b740955cd7f61c", x"3b80b255108940c9", x"e0ab367dbfdff85f", x"2ace361f3e1fa817");
            when 14702955 => data <= (x"f3fafdb822cb1c99", x"26ec8b58037457c5", x"594d209fd2523efb", x"9ee384c24a388e8f", x"5aa2db767ba188b3", x"d71b64c56fbba5a0", x"aad8ccb022f4161e", x"163ff9a99d9cbacd");
            when 13736728 => data <= (x"705dffa262fc8b3b", x"cc13dab4cf01fe73", x"5100a61ffb55fd60", x"2d5e4fc6d14e625b", x"e19a716b94b0c1d5", x"460a6cb33042e832", x"aa591bcd8d678ca0", x"b7d344c7b28ce696");
            when 18015564 => data <= (x"54d69633db74e015", x"82cc68abcec46747", x"1bec12b393327245", x"6a6b80b607a1cb79", x"86da1a86a93c920d", x"79076f3aa708f1ad", x"0a884267bb926779", x"87b13cd7c6b399f3");
            when 18491783 => data <= (x"da741e9137cf785a", x"7c52d464482eb1b5", x"b32cd2af4edf7358", x"8f5d215337464bfc", x"37f6ff7048da4ef6", x"e088f4c1f85e4728", x"f3c472099d42c9be", x"a1e1f03171c6dd24");
            when 5781756 => data <= (x"6ff298898def178d", x"cde1ed2fbe72e8e5", x"1841cc8c04477edd", x"1bd9331bdc3f115f", x"ade945110af7e554", x"fbca6cf95477a9ba", x"27b99ab75c9d912b", x"bf6a4df8ef9b7931");
            when 7042452 => data <= (x"7e241930fd3fcc13", x"5d584aef978e4cd7", x"985fd71c724d5a8b", x"3a4c3f90d71bca67", x"d6c25cba6aa40a7b", x"20a0492153fad493", x"751de37d75db8dc7", x"89253ae65ef774e5");
            when 5705354 => data <= (x"76ca028ee6111854", x"45134597929aa526", x"6d464301c41f912e", x"16fdd238c420f5d9", x"24910c2d113f0eaa", x"d1b9e66ef94f55ee", x"a3995891143f4e41", x"7d973f0d64e4067c");
            when 9593869 => data <= (x"d55cf97fbab3f119", x"1f12ee33fb9f20d5", x"bed1a979b53aed67", x"4fd335d83ddd5c2a", x"0ca3a1df58f34fac", x"8474d3df8ef9d96c", x"4d0686b35ecfbd19", x"976776467e051444");
            when 21612511 => data <= (x"c5c214e648d42488", x"0d7bfdc520ddbd86", x"b46c9f1260a9b7e1", x"07349d06b3953342", x"8af48465623919c5", x"eaf4081a2d35eb23", x"7485e3112db1e409", x"00fa1cdbd3ac1ddc");
            when 27508923 => data <= (x"6702b197ce744602", x"28d30ffd96aa75ea", x"3f239ea5229d23a9", x"b3b1edf6986e4227", x"621dd6649c952c2f", x"d98eb8c19d278adc", x"6189c4a9621982e3", x"22a07d3de715ae3f");
            when 31390496 => data <= (x"f389893e735ade55", x"49a8e6f12131f6d2", x"757531bb94020fff", x"7c050a0d0e188fcd", x"e975513cc1953325", x"4cd49da6794dc84b", x"b2ad510c960e1d0c", x"5cb287384a0461dd");
            when 5013670 => data <= (x"4028d3b044f35c8f", x"4dc5378ac1b74138", x"315e5b7d412b8b7c", x"59bcc8f98f0920fc", x"f994d940cfa33fbd", x"8f7adc56afdd9767", x"8310b60fb71b3cb1", x"aa4228a77ce24aa5");
            when 807656 => data <= (x"f0a529f1d9bc4c46", x"2bc6157a2a5d55ec", x"eef144936e8ab465", x"c047554eead2becf", x"edd85739a2daa700", x"8ace234e052a7ccd", x"28ad3aa32d8203ac", x"2a951d3dc3aa7660");
            when 28738441 => data <= (x"07169f372e65ef24", x"621d5b9d2838c292", x"996dce4a2ed1afe7", x"d452b854d313913c", x"616fc5a5eae249c5", x"a9123e250bc9ab9c", x"3de3d5a4c7398e47", x"ee53280bc683a928");
            when 2427535 => data <= (x"71bb967b75970314", x"98f337881b6c9d20", x"77aa462e6c2c206b", x"50ff63fdd1cfc31a", x"5df327119f4e850f", x"61a59cb815442c87", x"697ac5cbb5a70268", x"ca9a52c91d90f403");
            when 22697860 => data <= (x"d04bb16ae867ed3d", x"9c9e100991226ac1", x"cd5d2a141826b71d", x"89b8a0d232b2ecaf", x"0566f507c14891e2", x"9f2eab0b32f72090", x"2a9647d6ade5e188", x"a306ac40c54f0386");
            when 21854295 => data <= (x"a4454a4932eaef7e", x"3290aeda55d6961a", x"85e252f72c90e934", x"62df007d472611e6", x"648248cd64ba4017", x"b2df0004561e9e07", x"10e907914d54b61d", x"e0792bce817a00df");
            when 22472858 => data <= (x"44f26ad2ca2209fc", x"5e43b05c70968004", x"1d913f84a5e2a851", x"2922f6f63dd0b146", x"ccc9b3911d78c9fa", x"ac258ebc458a0ec9", x"acecfffee20352ac", x"bdcbcea7d23ea1e0");
            when 15675592 => data <= (x"83c6819efe6f811b", x"e958904b4b7dc69c", x"3e694ff93e8eb8e2", x"26666cdc9af4363f", x"a57507715019853d", x"a0b1c4a984487295", x"da836c4139adff31", x"4ede7c60ce020060");
            when 1367844 => data <= (x"1d150f029a61362a", x"2c77342184b4689f", x"3d61a36c9be89585", x"2e5c011be7d90b5f", x"bcc3a011e9c638eb", x"6929429905f80e7c", x"ec83a65e014f4688", x"9ddfc5d6c25809e2");
            when 28988214 => data <= (x"0565a9729e8b7dc2", x"b59fa6dd11953b01", x"7b403504daacccbc", x"8c039be8d91c410e", x"0d0a03b27c6f32f5", x"d97a277083fcd23e", x"63f40fe8462f2d93", x"58fa56d574f581f2");
            when 26632064 => data <= (x"62d8fa93230916b6", x"fbdf848978f44f0e", x"d537d0d625d66009", x"304296598e62c60d", x"2274accd0b14341a", x"b8c9e774134b84d7", x"264793b916cb1590", x"a88a6a55865f31e0");
            when 29268353 => data <= (x"18d03669648f6044", x"171b4054a99bb1b4", x"2b5c4a82e52fa34b", x"ade5a11bb0af0ff0", x"10302b656da16844", x"54fdc5bfe195492d", x"13ab46e897322e75", x"e0f510892f6a7844");
            when 17132889 => data <= (x"9c8cdbc2de230923", x"1bff26290d1f7376", x"ad4bb6304b948b9f", x"3365cbfcbc768a6c", x"11baeebf70a0befc", x"17c66f9ebfaa5e5a", x"b9ff5aaad68a0ae1", x"76202caa21cfbca0");
            when 6754370 => data <= (x"ed1d45f397696c5e", x"039dc798be225cef", x"b5134c53b2ab9168", x"30a676fd9005aa6e", x"619522a51b684f76", x"d5a0d151a4acbafe", x"29e8d7a9e3337f0e", x"be3f693a893e9d0e");
            when 29881364 => data <= (x"700493301391da91", x"be0c82c72a17fa12", x"a3e8f614c8c7ae24", x"1a880d957e881020", x"b5370d39a43335f2", x"e6bad3c4ca49be1b", x"3294d78c7552fc64", x"2b043d23ccb2e996");
            when 20189690 => data <= (x"b07087d313cd690b", x"a527346236e6ead7", x"0ca4563ac10f4601", x"5d624ceffdfaba9e", x"688e6ee0a2201316", x"436d769153b18a4a", x"27c796cf4d833c26", x"e466a025283d7450");
            when 18334422 => data <= (x"d1d3820bf340f345", x"b2c5ffd563edd5b6", x"e3c99447cf229ba6", x"7e3d22090dd821a7", x"6445c8a4b22354ec", x"73a3309590fbbb6b", x"a25271fd2b5f9f88", x"59ceaa5f649bd4bd");
            when 28148393 => data <= (x"b3fc331b0bd2d3f5", x"92d49b5e08916b9c", x"8f9a25b183ac1e6b", x"f6938f2d66f8e805", x"220804c7d8608291", x"affa67eb9bdabb78", x"68d3d80d4502c9ba", x"5e798b770586bb21");
            when 15994938 => data <= (x"5933f2c84510157d", x"a960cc3855cbcd1e", x"c22af57a3f6f8c17", x"044385f10d367388", x"97e830e705e4e663", x"38a1143e3fe014a1", x"eda88a8363fd38a5", x"d11bb94cf3decb5c");
            when 12921584 => data <= (x"b075b247beaa11de", x"ade2167329fef45b", x"6d2166fdd9c2547c", x"ca92f9d752ec83f7", x"cc87fb5b17371a02", x"514aeec00b4231db", x"04833a6c1d86f96d", x"722bc8ee9e5d489a");
            when 13700902 => data <= (x"e867171a5e6e0133", x"d683f95722f90279", x"acfcbbd156d6a0e6", x"a44575c6c05eeefd", x"085155f020957c91", x"c8e235eed843b4b6", x"603c74ef06ca320f", x"cc6c889d43e30549");
            when 4818104 => data <= (x"5c408bcc90e34609", x"48f2855e0ac29877", x"e974094892ce81f0", x"fe6eb2d8fa2bc5a0", x"6d4998a8f26a12ff", x"712cdd501b86a9a4", x"f6b98c9739cd3473", x"5107e32b526a8b58");
            when 31731574 => data <= (x"cfb4e08905c8c40a", x"7cb3914f7e6dd725", x"6339d7e62285443b", x"b9faff8934669ecb", x"d521359178f8b5a3", x"410f6ca495f89af9", x"51b6d053c6ea15d7", x"77e67602e47e721a");
            when 9697936 => data <= (x"4baa14982073ac56", x"886df9f4e8119487", x"7e575a5fde64e41f", x"a473e7992be2dd88", x"e5fd7b48a5a41a15", x"0db6522d3b061eb9", x"6166f7b1609a7e10", x"aa1181026bdf2891");
            when 27534836 => data <= (x"37ce6a5df34f7eb0", x"a72fecbf2b69ea6d", x"c2a1d8f574e4f459", x"8b1baf8b185b4a08", x"6e112199dd418e94", x"b2bb7512e928a2bd", x"f8d81784a28a9efc", x"55cdbd4eda7ba9b4");
            when 8988427 => data <= (x"1ff3cf38b0bec7d4", x"b398388972d4f692", x"463e4f6a645407ab", x"a1fcb1f035fc2556", x"cc978d761c33ef76", x"65b23d55d3305ada", x"d8436356c4eea6de", x"c03d907407a19f2d");
            when 8751918 => data <= (x"b4c2e1c0a909cc87", x"654d7acbf85f243e", x"5eb2ba32daedbda9", x"64898599bfed9618", x"967ef7d7751ae1f0", x"ead2e104e261600b", x"0892eeceb244587e", x"78560e6ffbf3118b");
            when 6916818 => data <= (x"f328555bdc525bd7", x"1347551041a195e1", x"0bc4eb7292954bc4", x"5afdda4fcb198176", x"12d7030b1e7f710c", x"57d51efbdca4bdcc", x"09d5969dc5a0f7dc", x"0cd4323ce2aa4137");
            when 8137595 => data <= (x"b8363b64ba4b1857", x"37490ea9c8990592", x"d9b2634177b61398", x"9afd58d62322d602", x"53ddeb6aa9b61ac3", x"843533186b7ceb7a", x"3ade3f73ffb61250", x"d2fa7e499a9428be");
            when 3316877 => data <= (x"dd7491d364481bdb", x"341e21f43a85f733", x"4936147d6e8886d3", x"56d098e9eac3e905", x"c9594bba41e513ec", x"2dbfb0f72ec7b18c", x"e0313ac11d88bf18", x"1c7b0ee719bc024e");
            when 14387766 => data <= (x"2d2d4c78c9a3410a", x"14396a1f0bedf8af", x"6f2b2cec378c321d", x"76826d6a227f923b", x"18777e3209c4593d", x"e7646004b30a3e18", x"96800ad1c952bc26", x"c3753d0f9270d707");
            when 1849707 => data <= (x"0e4d6976b4d610e6", x"1b4cea79388203e2", x"45ff0ac24d166c63", x"011ca1f29afbe076", x"7092453c1c3ad226", x"8a898b234ad0b805", x"22a38fb207d7cfb8", x"69ea11237b3c6024");
            when 2853517 => data <= (x"00e6a3ed064187c3", x"6cb299ec73197dba", x"69d1d6df522b585f", x"f5f8d61884e129b5", x"693c2ff6fbf5de31", x"8a5fffbd76e697a5", x"d2de9050e813c149", x"0271f341f091e02b");
            when 14893325 => data <= (x"6bdccc0edaa2fa13", x"4c516a10b6382f79", x"27731b94fa6c387a", x"703aa4f7c30d0942", x"1b78f3363610abbf", x"d04a09e328e121aa", x"f1ca13f5f61161a6", x"18cf1279e539c5ce");
            when 21487187 => data <= (x"3f32d0b312bfe7d0", x"98e24b3019456011", x"6f57319e979a5a4c", x"c9ae56d8e8abd1f0", x"a03a8b2812f5e038", x"34ffd193e7e4b4c9", x"19615548b6acaa68", x"d25a7f106115c57c");
            when 29694309 => data <= (x"c546baf7775582de", x"49fed9f25dd0f456", x"3e6305fb6d16e19c", x"8eb72dad47bcf1cb", x"538af89af92bf796", x"222a2eb6b74f57b3", x"1eda85c52b283263", x"2060e10ad1db609e");
            when 31048618 => data <= (x"2ad9726d6c71419d", x"8f30418cc698096c", x"f85633615fca4a1a", x"7b7a68df1a6a23a7", x"5387616373337ddb", x"e9ac4cf24ceacfc5", x"38c1e2ff282e042e", x"b654ed65d7cba07b");
            when 8837226 => data <= (x"d845a8fa2e6dc1b3", x"27078c2faaf9ee98", x"038f2a6b4e3e89fe", x"f85ddf8b4d572f62", x"447d5af9e4017d2e", x"7b9222a11eeebfe6", x"47c83f2d6e43f60f", x"ccd7805cb3102a47");
            when 24450937 => data <= (x"18471a644103a74d", x"576c261532ccafa9", x"37df2d37cdd12dde", x"e866d638d03d4888", x"91644a1db745e7f4", x"23d36c3b61f0db92", x"43c54ee4efa1f98e", x"1f9ea0821e4a67f9");
            when 373147 => data <= (x"9cacf26ffb34803f", x"d9287b2815af5902", x"d2546c22453b7d47", x"59059467db5a4882", x"1d45f5339b01a743", x"9d6ca59580667c6a", x"41d9bad48140031b", x"99b086c061f46187");
            when 30659241 => data <= (x"aa70270b3356b402", x"a3a5eca9dc674afb", x"226ad4fde5bcbb33", x"f2fdcfc004efb510", x"61977b021a311cce", x"8ab6065c7a9fb858", x"979ed5befb94c1ad", x"1396bb0c0130ee85");
            when 2118791 => data <= (x"76086457d7d04d13", x"93c7700cb4e85550", x"01345e6c191fb830", x"1218af85d9892449", x"c55ca61f332f50d4", x"593c9b5ee84f1fdd", x"2f1ae8005bb2f8e9", x"2ad160e01710bdc6");
            when 28655712 => data <= (x"25604561c5481682", x"54d82f15e66ee002", x"4ccb540b279da489", x"9206845cf2ab62f9", x"51ea43a49bebe1cb", x"f6aeea4b3f7a59f5", x"ca889f34f31e9b97", x"3e2522c99bcc66e8");
            when 21934540 => data <= (x"8d6c47014b9e40d6", x"9c05c3668d637e46", x"8cbc4430188f4150", x"375396eb8a573ce5", x"4c29355ab0a1be0f", x"6ac530a633c961eb", x"398f9d2803fb090f", x"294ed657b073da7a");
            when 1168886 => data <= (x"1b271734ea2a6fff", x"12f827a2dc6772c6", x"43f7c08d812515f7", x"c87207d3b02d79dd", x"b1dba394406bd951", x"e7dce20d9f786d04", x"1a5d8e2e70608348", x"4acd5f7cc642c9b8");
            when 6019241 => data <= (x"a90aba816754beef", x"7cc2dc35172a1be2", x"fb8b266131465216", x"08d30a2bacadc49b", x"54bce5bcfa06cd73", x"39356b492fdd0c91", x"84267c47f1f5b9ab", x"010c913ec237d9f4");
            when 33739376 => data <= (x"9c2ddeb0e2610cb1", x"481b8e0bd2c7b953", x"79f10ad84b7613d0", x"8ffa81c89c7d3b39", x"5e5cdfa2b0a94361", x"96f55bb6a3feb37f", x"e3979f34c96461bf", x"f403a7d53122b138");
            when 19136163 => data <= (x"56cc454b1b5abc35", x"859cee5e2a7f58af", x"d75f6627614d828c", x"60a25ec1960e936e", x"e454cfb5d943d866", x"883111da480a0d95", x"8f3c205e087734a5", x"51fc3615a5133527");
            when 10471497 => data <= (x"a58fd48660dc6918", x"e611241f440a99b5", x"1b8f7db8adeeab61", x"bc533c05deef97be", x"91c0ab4c62c72768", x"b7b45f786c056439", x"cf7f441ae96b0412", x"a2ffdc5d25f65c76");
            when 853972 => data <= (x"0d0314a1694f64e4", x"6fc68ac5711f836a", x"92c5a858b4d9b995", x"c2b81a3c2827d59f", x"475bfa6a7aa26848", x"7e8eeb35c5f97d69", x"ce44548bc857988a", x"c72201e47ace5dbe");
            when 18756850 => data <= (x"99b14f71b51dbcbe", x"ec3613233ad07a54", x"2cfe3587eed35655", x"d70b4d1483c11183", x"1ef5870af88eb86f", x"1e563c630170a5de", x"2718a57ea2225b40", x"62a788a6dd69a96a");
            when 9692661 => data <= (x"dab234f78ef593a5", x"1420f9f3c9054c59", x"595c053440caf4b1", x"44c1716721ecbfb3", x"3f94b3b1351a981b", x"8970d964d79b85fa", x"806d36b8911e10d3", x"0874e3399391a2c7");
            when 10555300 => data <= (x"cf6d5922ebd40d68", x"20c2651f88cdbbd7", x"a8f8542f3b6574b7", x"32382f3411839fe2", x"2473724cd8fa5a5f", x"32d8d92b925f9213", x"34897e70edb9cdc7", x"064f8fc9a8298593");
            when 10681661 => data <= (x"3d2fa9fec0ef36dc", x"ce868de5eda37f75", x"501135e498ce2f84", x"50d67828d6ef7525", x"80aed6e5a49d8561", x"de0f4543727dd4e1", x"ca53b190a573e2d6", x"5d8f4819ef9e5a35");
            when 3944881 => data <= (x"5dfc75e7f96a6354", x"da204d319b05f855", x"4581f0a32d31cfd4", x"08de9a3ee5e58bf4", x"e1f048a49215d6e3", x"f69c8e24576b54ab", x"ad8aae6587130f93", x"eb8f70622e578bf3");
            when 4781777 => data <= (x"66bb71f606a4f1f2", x"6f9e61be460276c3", x"e95dc75776e016d9", x"8e34a033ba439bf8", x"1bc42a5c709abe51", x"a5cd303b0109c4e3", x"50bb3347e4387e2e", x"5d4e90fadd043231");
            when 11733857 => data <= (x"efe0eea8ddbb4f83", x"2bb949a9319fc576", x"58bc36d62ced05c1", x"cc946e1bb46038ab", x"0b458da7949076e7", x"45db34683aedff15", x"e714da0c8bc75470", x"63fd199716d08dde");
            when 11577339 => data <= (x"c0e39b2df44789f5", x"0568b71dc7ea4db1", x"503880b44dc11eab", x"a789ddb612b6e6a0", x"cc383ed924e0f42a", x"695d09e8047a54eb", x"e0bede5c8667a9e7", x"99b0da127f8d4844");
            when 6793859 => data <= (x"b5e4cdd311e3502f", x"798d3a5ff843efb3", x"7218d1a8a046a384", x"3a35ea8e93845e3b", x"b872ae1abbbc8257", x"a34fc063d3b1853f", x"0f48e7441638573b", x"f3ca1d6362f88460");
            when 27826422 => data <= (x"01aebb2bfdbcb795", x"a5716994c30c9a43", x"d5f1f1b6d5da8fce", x"19fc94dbabdc8cb9", x"728db0f22f65ac35", x"9b18a6e3d6a69d79", x"0f931c66e43c77e0", x"0b340c6910fa628b");
            when 5413510 => data <= (x"c1cd95bc6ab44c3f", x"7ec70ecbe9987d24", x"a35a67f3f9db2dbc", x"d6738370d98cafe4", x"c568af4e5310040e", x"ff23c3e01abe49ff", x"bc4537a8427b0cca", x"f648dc333e38d943");
            when 19308268 => data <= (x"6f39c4995cd17a6e", x"54c0d484e871f93b", x"91824097fa10c9e2", x"a1299da490a1e921", x"aa465194d3104a3c", x"1a9604ebddaaada7", x"9d5de011950a8b4c", x"e56dc835db1b8b7b");
            when 23090610 => data <= (x"be0d99f5ee7ac343", x"3f98165538595786", x"cf924760f9aed678", x"5b55e3e84ad5c633", x"8088364e69e36945", x"58cb069a0e406276", x"4ec4fbb408a7215c", x"f98fb7075cb9674d");
            when 3692080 => data <= (x"c0304fc9bdeccdb0", x"c3af86c3d9de21f6", x"8097255aa37e5fd4", x"873c2fcf6b4846af", x"a30b296ac3ebef6e", x"34956e1a05154501", x"8b44893f714a22ec", x"7c941b679a2b0474");
            when 3893551 => data <= (x"e2076e8747877136", x"523e89d7ea9c04ac", x"96246711b488f64d", x"af8b8cad2eba93e9", x"302de3e4079a15bb", x"ab2b0237ee3e8f6a", x"59b7f8dc457d58d3", x"62dedd838a6edc92");
            when 13761983 => data <= (x"7fb34aa39ee326ee", x"628d9f4dd8cf8ce3", x"332ee101929678e2", x"c561183cfc561e95", x"8028810dd135d991", x"47034f4ff156ff27", x"f208fa23aeb96162", x"616e3df9a3dfad42");
            when 19206237 => data <= (x"42ebfa01f027019e", x"9d159639760b9045", x"bcd31661cafcf732", x"21c8678860e18927", x"d9e39980504212a8", x"0b5da52043291bf1", x"742da965d2cfe431", x"f9cf7bf5af8b3ffe");
            when 479657 => data <= (x"2b4502b6152c7e26", x"325b4f295be98d58", x"571582341084fdb9", x"cf55a252beece272", x"22053c5716f23980", x"9ac4410dd8660f70", x"fbee6c43e351f534", x"11685c842a4c959e");
            when 24056970 => data <= (x"4e9290e403b34078", x"88927c38315f2ece", x"5340a8311bec74c0", x"7470974b117fc344", x"60cd92fb8596d806", x"2546cc4087d8c99c", x"90562dea7e14e5bc", x"7b188f84f9b41785");
            when 2612068 => data <= (x"eba13516e6560e8c", x"f164751db3de6972", x"780b2bb396ac57cf", x"5aa65cf44a8c7d87", x"8b9a874645c34554", x"b16e83801ee12dfd", x"5bd15d4185f983fa", x"392e4a229b433c90");
            when 2019342 => data <= (x"3b9cd3d0e214915b", x"1e0f751fc4a9fbc5", x"bf7eae57d0a183b8", x"4b46d5c9cba21d55", x"df8d45c1267a56e1", x"cdcac43f7e8590c9", x"780d1a77cd702d1a", x"4db5171068e86500");
            when 6752191 => data <= (x"911923a5114eea64", x"c35654a1c358bb4d", x"634e7f26c1048551", x"4bda2cfcb3c0c87d", x"fae484e11f4a4acf", x"d2c8246fbdc54a1c", x"cad39a0041ad64f3", x"0cec3b5b9d350da4");
            when 10438494 => data <= (x"0851d183669dc0ae", x"1f8af547892a4ab5", x"3714e0bcba306f60", x"78e862513573b4b4", x"b6a707accd0e53d2", x"b50a9ea173efb4b1", x"aa9fcfd70dc37b38", x"dc92266d54b90f59");
            when 11796655 => data <= (x"042f4b804c0d1c12", x"704464cacc3605a1", x"4f97b46d580e494e", x"3e186ad443f3d335", x"77e08957656bcf6c", x"315063558386ec97", x"c021d5b6bd810c77", x"92e43814ed4a2581");
            when 5256098 => data <= (x"a1b80ee08f9f9acb", x"428090fd696a0190", x"9d498182732504c0", x"2206bdbc32a57687", x"dbcc9fe716bd27f2", x"9b32df0393425e9f", x"9a19b42415485b45", x"66c00499fcaaa6b1");
            when 13113849 => data <= (x"aafe81aec2e8f91a", x"e425724f6c8352f4", x"cc9ef76008556b45", x"fe9610b86bba7cf4", x"5f4d07dba27bb474", x"91648b59eb79de29", x"9741415dd1460599", x"c6563f8f6c04a1e4");
            when 29568459 => data <= (x"0b7aeb88455e4d62", x"47e9a5039d7e363c", x"4184934f37ffb0f5", x"bb8cc8afd085b550", x"e6ea64ab2813fa38", x"95c291fd3061b2ea", x"9bd9d1d971ec4282", x"c6f3f217450836da");
            when 29028135 => data <= (x"dfac18ff934d8b4a", x"80cc4949e6c5e73d", x"f7b06c736979a0fe", x"82074fc5b746c73f", x"e339e2bdd3e28580", x"77a37d69c7a16105", x"710c2cb512b1def6", x"1b28b578e2752087");
            when 11041808 => data <= (x"0dd4d108d58ff668", x"45d1752e8bd1939d", x"09cdcd25b62857c7", x"0c903738dde394b6", x"31496cdd145edc93", x"f120145ce4873dbe", x"a3e6c872f812162e", x"03b89face14a091f");
            when 18430445 => data <= (x"b0c36bbbaa01c418", x"0f7b52eb379dd7ce", x"577be90171ea87ea", x"6ccd6c9b6db54722", x"ce66af59465a4f5d", x"1bc1ea8f133800be", x"f4ddb78633f64a2e", x"1994c8331f607d6e");
            when 12885154 => data <= (x"3c18156c4808b3a3", x"abc069359bb354d6", x"54555fbb3380eecb", x"d0076edddb70b4eb", x"33935b77b4f8d420", x"04474a195da2c0b9", x"3c84f98847f6349c", x"2db97355e078c971");
            when 7616356 => data <= (x"da3b1fa8703bf421", x"39a5ffc75f5c8adf", x"31e9bb1c1f3c5e66", x"7903a181dbee9ba0", x"d279ba899fd86e02", x"7f2f87295b943b04", x"ad6871613fbe4b27", x"741cbb1293e1bd12");
            when 32333582 => data <= (x"a7f3ee0a1bd62795", x"5a1a797bf4ef88de", x"b94c41814393c3db", x"6ab7815991445fbc", x"40b162cb0373dffd", x"e29e835b72c66e76", x"9281ffbf59a7cd9e", x"2bc49908fc7cf296");
            when 10262700 => data <= (x"f3dfa8de47486fa0", x"bac63af0a69e0378", x"5051dc9ee9eceef1", x"12869f05577e1be5", x"e12d14af2a1316b8", x"506178e21be27c08", x"be7156ffe32438f0", x"b38b8b47ab71139b");
            when 6984499 => data <= (x"11fe1fe1430e7ae6", x"25b131ef9a6d5388", x"26a75ef72ce6c34f", x"8579d9a9312c752b", x"bcb040615f4046c7", x"df19bdd1a7dd3136", x"b15628f195fbeea9", x"809deaedeca00659");
            when 9794084 => data <= (x"89e8e8c5f3c462d5", x"2207e563c0cbc165", x"98e8bbe4987a678d", x"1feacd23739ac79f", x"0b032046fcab53a5", x"b0fd3168d3fae8b1", x"24de820f0c5126b0", x"a0b64600b5439281");
            when 26968334 => data <= (x"fefc2763a8f932cb", x"2eaea9302bbc30a5", x"ea18af10babfde04", x"da8d27e443e26a20", x"29291028267c646d", x"d8df5da4ba5fd5ab", x"9fbfe5a88e9b9652", x"fec39c8ff83a241d");
            when 24643914 => data <= (x"e8a30af6290b1022", x"0ada97787129d70d", x"8e89ed8c344f6c1a", x"ccaa505c03b040cb", x"c05b800fc3020b21", x"7fad5206788d85db", x"2e2cec174e40bca5", x"1d2e6de659bbf89f");
            when 18400342 => data <= (x"d2ddda495f2c02a0", x"d771d2458dcaa291", x"8271bfca3a700abe", x"b7ec6fe59b15f705", x"62db24dafc35cc53", x"84c2c5130155ee6f", x"3775e302478d0f78", x"ca5bb6704e6fcc1f");
            when 25592303 => data <= (x"683cd0bd79f19b05", x"7db063b1a1c07134", x"ef69bc5ddd68f0cd", x"efc0b373b567e947", x"111d125eb0cd0109", x"c3007a79e7d942c2", x"3bcf19dfcc6d73fd", x"0f3999bb02577083");
            when 10584537 => data <= (x"882dab5c6e805cb5", x"1d02cc53a70e7916", x"e589d05b1598ce35", x"0b1147d516f678f7", x"4955b52c3d7df92c", x"3f6fe886a9b20cfe", x"e987baa4bde7fea4", x"2133182a33137dd6");
            when 22117121 => data <= (x"748c411f29c7f6f5", x"70241a395858ddb0", x"602a5b9b7c7cbef4", x"b4da2e3f6c9bb45b", x"63694cea2fc9eab5", x"c5d7448746916b49", x"b3bb676ee4897535", x"797eadd28b53271d");
            when 29360110 => data <= (x"fbb4a9a1197d1987", x"4f01a129d4e7df6f", x"b45ae0f1ac2310b0", x"2632c192a0a4f8c5", x"2f4d420826d1d9ab", x"89bce73229072e04", x"6e5deda2eb1d291d", x"fcc5ad29551eae5c");
            when 30137648 => data <= (x"bbdc998b468af3f1", x"8628a53587f089ac", x"b135f759402fc182", x"e5a53f3970936eb4", x"ff64e0ad9ed25400", x"41c5843cbd56f35b", x"d36e37f66b84b28f", x"7e9e295adc63df14");
            when 20365803 => data <= (x"451c4163625096e6", x"02ebf7bc0244a991", x"e67d5faf1a4de77e", x"37395cb2fb2236ee", x"77900861ea26f13d", x"852a88f93290a68d", x"dca93ea80b544c4a", x"910f6eb15d80b186");
            when 8999765 => data <= (x"59e91d80fe6cd0ad", x"289d658d395a540f", x"c287e7b21f67b429", x"5f78f8b02f519b91", x"f3537a200bccf3ad", x"71e6b53339d01999", x"6069f3fcc3abca9c", x"4809763b2babc549");
            when 17165459 => data <= (x"1e380e7ad2db0a56", x"303d1bd8139eb557", x"1ca1d0edd6795bc5", x"8a53591d1d7f7031", x"f4ccb1fdcaaf0271", x"ecaaec8d7d5b292f", x"64884dea3d2bad1c", x"5331443fd1d1a5d6");
            when 12838674 => data <= (x"ebe0b1c0c5d7be7a", x"9cc5bc32524378ad", x"06fbaabd558e79a5", x"84adb360835b6b0a", x"1314e80fb4492b3c", x"bebb9e08e7a41233", x"0383b03a88aa56b3", x"99349765518b5561");
            when 26990807 => data <= (x"a0dccc74f0db5760", x"f3ac47687d2a7095", x"94bbc5f1e2fc9c81", x"72431fa85f33c497", x"75ec9e7d95f0b915", x"86b68cc066adecf5", x"b00e4c5c4527135d", x"a61adaf102cea822");
            when 1147331 => data <= (x"ec24e4dfb43ec28d", x"48fc3606accee559", x"a8607dfe7bfe4ac5", x"7c2542e67f726884", x"115b4d95e1b96d06", x"09beebe814213972", x"5de5c37bccf0b07b", x"34cfd366cbeec625");
            when 27934568 => data <= (x"92b94d15f5221c0a", x"62e91ca18f8e6f7d", x"46d544056f315403", x"dd2c6d4a93b2f704", x"0955ee91336f1dd4", x"8673fe2d7f233803", x"b79f33ea9206f0a5", x"e1c661baaadaa1b7");
            when 5677994 => data <= (x"38d4cecbf721ffc0", x"9c2cdd84c79dbc41", x"9d5e9587f63f6fea", x"6413ac01a0e1b66e", x"16750905f382855d", x"bf58dec90d6e4957", x"f314da5ef71bdc02", x"12d9edf265da86c8");
            when 32202233 => data <= (x"15cd070108a66458", x"59f110d2e0b75608", x"945091fec1319244", x"f1f4d9edceef8425", x"ca15a6ddfb9ac012", x"c3515c967790f7b0", x"cc716504783b6040", x"62cdc66d546cace4");
            when 14621205 => data <= (x"cae7d2176a50790c", x"3bef4672a198adb8", x"cab271e4422e38a2", x"51f02f6366af04d1", x"f905fd43bf70dfda", x"d6de71af137094d2", x"3042a79b5f76ef0b", x"fa6d04d2fee429de");
            when 17149034 => data <= (x"4fef1d5725109092", x"04d835f3c16206a7", x"eb16688f5647c38a", x"6468e4afdba70bd8", x"9076f30b03700d7c", x"0229efe608fb7af4", x"87869bfec888f623", x"206b94423718a25a");
            when 20403280 => data <= (x"52b2b9339b0dd171", x"45492bd20dcc2f40", x"3b48770eb62b7f02", x"fa1aa908d15e8258", x"bc3359442d23f2a8", x"7d13b92f249b705a", x"88272700e866ae52", x"acde71db348f4ca6");
            when 22695935 => data <= (x"52ad71735ea11de8", x"f6972f93e6a41c88", x"6923326b49e239df", x"8ae0e79ef023f96d", x"ac7ea489594588ea", x"47ecb640627ad12a", x"a4416e6cd12b9ceb", x"1900095525fed18f");
            when 31555839 => data <= (x"b945a20af1ef2d42", x"c0da13c33d238df8", x"b74305725d1b8496", x"18048741799366a5", x"2d726bfa827dd5f1", x"61f5059e2a31aebe", x"8a594e195861a61c", x"7d93acdfa1ebb74d");
            when 9348579 => data <= (x"a570c448da72f301", x"616ed69278163341", x"e2964910b77aed6e", x"5d8e62b6981e9e5e", x"80a2662f0bb6f069", x"c258de9ef668e08a", x"803c3e2168e3c6c6", x"c5d99fe3121944f2");
            when 31127845 => data <= (x"eeb5b5bc8d9d011f", x"3ad25abf4ea28dd1", x"a4b53e1aa249f0df", x"7e3787f88797ff96", x"cd1c43193c7fb53f", x"45619434519c0660", x"aa5b547042a2ed5e", x"2b798be3ba5de501");
            when 3628730 => data <= (x"624c0ba2a26e665f", x"90f6da669da2e169", x"fb2d109603a0f328", x"893a15b94a194a03", x"29796447574b1a97", x"07bbfbc29b9c0e96", x"19dc78726c8f99c9", x"e49821c13e820d4a");
            when 6066997 => data <= (x"44b1858c45da2ed4", x"c81cd58c634c4040", x"b3cb6e7b34203c6a", x"6dfec6ef4e014236", x"fb5d0ce787e0f6ce", x"5c4e5bf11ccb83e0", x"5fd9238b6cf6e9cc", x"aa660a5e3152cb4e");
            when 6071946 => data <= (x"7556bbfd305159f2", x"bcc6103f3a91fb26", x"b03ec2e184f9b719", x"e74f4af0cdeefa07", x"9c03dd4ba0ba19bc", x"60ee3f99cb3aad2f", x"ac2c350b56a1faab", x"fcf21f6279fb9a68");
            when 907045 => data <= (x"dfd5a2a14c61a169", x"17f068c7304cd67e", x"37b5136d300aa7aa", x"a4bc576971dc64d8", x"e3da60dec9fd4f4d", x"613bffe8defda221", x"a1442c53e78c7b27", x"df71189a1c84bacb");
            when 8799251 => data <= (x"57a4c443caa11466", x"0a185696583b5567", x"829ebb6d66874d6d", x"58feb32e101ee25a", x"ba5470b562631639", x"739eb7fcd54c558c", x"232003fa83a353ce", x"b1b420bee37afcc0");
            when 21242395 => data <= (x"b1bddc857b48fe2a", x"f9f28f44542de94e", x"e468c086e8d9b3d5", x"6b8bb5ecae325245", x"6ee2c4f21d874257", x"c83d475917bda1e2", x"4b95994ff0f2107e", x"0e5f528768d2cd2f");
            when 28187756 => data <= (x"dc49b0c1043e99a7", x"72098ccc3e87c482", x"bbbb3295723f7896", x"142febf690548d3b", x"1223655ccdb0127d", x"1eeca16af7bdd31e", x"e6b4e01fcb0aa0c9", x"e51b2af74e446e72");
            when 11152050 => data <= (x"699e4fa61dbcd84c", x"04b51b008c2387c0", x"67edf23697355ea8", x"df178ea1fad72228", x"4bc39e625e288f2a", x"dadbe5c9092960b9", x"1e136376148eb306", x"0bbef2dccf98d62d");
            when 21672413 => data <= (x"6c1bfc28765a7f6c", x"b46538480caccd3e", x"61e2a9ac3b6c9670", x"749e97bb9c047608", x"b07aa9890ef8a2d8", x"52fe03e5bc3e4658", x"74127f38349d59e4", x"7be110ea5033b9d3");
            when 28913777 => data <= (x"831293042c1416fb", x"35ee8f5fde95f9c6", x"7d54d9279731c646", x"86e0d8edceaa56e4", x"436d79d9c64e72ce", x"8d91ade5e83c4a87", x"91b9abd7ebca662e", x"8309a58ef3a7891e");
            when 11118018 => data <= (x"5730f4616599aa39", x"935e06c55db4791c", x"e86a98fc5d598bd4", x"84241cf2f73c499d", x"e6621f6b5137bfd2", x"094fa170196f40e8", x"0c6e782943f45ec8", x"e2b4b3ac9d92a933");
            when 16947447 => data <= (x"bd7949f08d81027f", x"bd0e75845e25e970", x"1480a8e07bbd9353", x"ab7a0b1722622531", x"90c916dba0135b0c", x"4e181dda3b5cd7ac", x"e5bdca80c765b557", x"b93f7ad5ba6a3f21");
            when 6081045 => data <= (x"8cbf47b087c0b820", x"0704f0f524dee2ed", x"84179da37684526b", x"aab84ac819b2f56f", x"7db4b784bb2fd648", x"25018903adbec965", x"5c01a56b2004f929", x"7e2e74445256ca4b");
            when 20006677 => data <= (x"429fe77e6346a21a", x"b900ac78b3d24206", x"faa3bdad667de0eb", x"91ea8d96fa002bc7", x"0ffb06f946c6892f", x"b8cba34868c53b63", x"45603079a21f7c8b", x"e204daac7f2796d5");
            when 30315132 => data <= (x"4fd876e08cf23b38", x"6f1ff4b7e1962547", x"d9095b4ea2679a8e", x"c2dffaa34e8b0cf7", x"a6af0023c75eb143", x"1516750a97dc3af4", x"f58deb1b2451f923", x"18d3530e55c595a0");
            when 20617860 => data <= (x"3bf1d4551cda1c92", x"5f4f797c1576f156", x"8c35727ab4a4d412", x"7202c3da187ee017", x"4b58aa6729c6ad41", x"14661b3d76c393b4", x"1bafde05388cfa1a", x"1c6654709e10e7e4");
            when 5735111 => data <= (x"4c5a5cbfd5ea4758", x"5ee340e45de7a9e4", x"40faefc4c3e4ae77", x"4a8fdb0ae87d9837", x"9b6a70a7ad4e64a5", x"b4513af9bb845c89", x"b57fff210cfdd9c2", x"f987c37dbbf0e642");
            when 15856168 => data <= (x"572c8bfc2578be9f", x"4b012f8377e0204a", x"62d1da2a39a9e856", x"230722cddfcab3df", x"53fbac1aaf286922", x"fe5f177afa63c586", x"f6491bb1ad4e9b83", x"d38ebd64715926be");
            when 5324944 => data <= (x"74426e12cfeb03aa", x"ed6c128ad2e9eb74", x"c1fa452ada81e089", x"e1ca4c10b8edb3ce", x"43d2e3d2489da8a2", x"3a26ca7952448b56", x"b1079ff219a6933b", x"bb4d0d168dfbfc2b");
            when 28330428 => data <= (x"f4063b359ce8eed4", x"02f1077e1f1cbc01", x"f6706e9fc59d0494", x"1a93f10d511ec67f", x"f4a4a41c224a90e1", x"7bc3e1a3f4f07c44", x"df3e772eb424ffc8", x"612ea4de18882254");
            when 5256859 => data <= (x"0db558e564725ca3", x"bbf64b3109dd8446", x"2c924edfffeb8f9e", x"2cb4cdf2a22c21f8", x"9c62dbd4638706db", x"e32ad3f7f5e3041b", x"6c8b8e48a529b9d6", x"7b2d37c037d87601");
            when 31338249 => data <= (x"a8d38451a898eeeb", x"684f51fa1feb6f1d", x"fd69fc6875ee87dd", x"5a6effd22703c29a", x"2e3e419e625f5ef5", x"cb6ae7ba62049ddf", x"f87e71bacab59b05", x"7f32234a17c5d67e");
            when 8780700 => data <= (x"cfd1611595b531ab", x"e08edb82b39ff84e", x"43629a7215bbc385", x"39f0fb4b936981fd", x"76e86a0a2d52715c", x"f2545709c8c5ff6d", x"8eaba98e7727ae2d", x"513ae245311694cc");
            when 15098594 => data <= (x"eed7b736fd2b1cc6", x"e4e9cd8ccd3841f4", x"8b78c2867ffd8b5d", x"260f0b81f6f25a87", x"570d474b0957ff1e", x"3aa74cc18b45b49e", x"d17efb84d7005761", x"055b69997c429fcb");
            when 19965769 => data <= (x"1a9285e6dc95b089", x"8949f2ccca68bbae", x"2da9b88b7042cff0", x"7eb9efffac99e85e", x"0a7a460e6d99ad94", x"6a9ba2459005fee7", x"f34c7144980a6294", x"fb05214d93e579a1");
            when 31045408 => data <= (x"4ee805de48d33b92", x"acbdc530677d3833", x"a24cf4e98d48d51f", x"a24fa37e859635f8", x"41d8fba799982f53", x"302cd738f48e5bbc", x"f8a403c9d960e5e7", x"19c7c324bf9da6b5");
            when 11653512 => data <= (x"bb1075d11e6f7084", x"9dfc272934ab7118", x"700b7ffdde627c57", x"7343bfc1539864a2", x"f114633522878a4f", x"6964f4779b0ee134", x"7b29ae0fe7625fd2", x"de521e4e4bbb87c3");
            when 22029067 => data <= (x"ee34481c0f8c76b2", x"daaaeeb6bbfeb7d4", x"c15893f6c869f9a3", x"7dd60cc589bf3728", x"dbb98644ac147805", x"65ba570bf087a2fa", x"2e0fc6925ad435a8", x"e3a368e9a09ce7fb");
            when 29705322 => data <= (x"39db3670fb1d6b54", x"01346bcb0b63361d", x"d80d652a0e2cc1bd", x"a98383f1557d3ba9", x"1298f63087f8cb6c", x"7148e0ca50689a9f", x"245ce667a5a25cd9", x"79df4a2ed84e4212");
            when 21031669 => data <= (x"2d31f9650e9ce60a", x"43ed883ca31e8560", x"842c7dd633f43e50", x"c9341019be19f753", x"d672464f450dde85", x"be07974935cc45ea", x"a7eda603f62f9b92", x"5447efa55535a967");
            when 29795669 => data <= (x"c8b295f45aa7027a", x"2c5760d3d0a23a4e", x"aa3059dce9cdc902", x"8287dbd3d7a1744c", x"37586654b091d054", x"23fdc049effd5e9f", x"f87c9a958bf59dd4", x"d671173fccff1178");
            when 32023572 => data <= (x"30fb8b50a5ef1cfc", x"8200d83891307b5e", x"70f047d3097a0665", x"dcdae914f176d40b", x"30c662158bb11858", x"5aaae38c78471124", x"9898cc21d24514cb", x"60c208f528878920");
            when 23500373 => data <= (x"dd542e6d96beba25", x"04a05df24ec7d817", x"50c28b074cea5726", x"e5bd4388ca33db95", x"ff9c8e6b5864fd32", x"3d9af55366562443", x"d516c3f17725099f", x"30c56ad752ac0ba1");
            when 29747228 => data <= (x"7714fe492341e8ba", x"1fd963a296e1f015", x"6ef5fadb1c4c69eb", x"7cf08ac2bad7263c", x"4591e7ea143461d1", x"511e30c8a4bc81d7", x"87411c91b0d4e969", x"41717532dd4e41e7");
            when 7128926 => data <= (x"fe92e367f815e494", x"b1608d7fea023c88", x"a358eef21e0bc896", x"9c3a25a59c583353", x"367f591a55b0fbf7", x"cdb3225f8c08ec14", x"ca2b9ba0f85d8353", x"25c90f5ba87a24a5");
            when 5994702 => data <= (x"139f6b793efd7ddc", x"9d0ae174363f83fb", x"9c8df145e80fe638", x"5ade562f552b0c7c", x"435b388b0f92941c", x"4e47c6209388b6ce", x"e755a3a0edc827be", x"706608a70639bbfc");
            when 17111435 => data <= (x"dc0cdd82f0c43271", x"3835dd5cfd899ec9", x"12cfe9aa9b5af379", x"a0c3696c565ee7e8", x"6cce85245e1d436d", x"1cddea6fd34b0913", x"82842574f10ef0f7", x"7ec6646dd86184f1");
            when 9161655 => data <= (x"2798da7a514747ff", x"c6aa61a18c033e4d", x"5649849ef8e97c45", x"e92a22ccef95b237", x"04ae753abb369d8b", x"e1c8388933f82c5e", x"ae22b0a56e76fbbb", x"fed739c8da0e1a27");
            when 31797627 => data <= (x"c9402136150c2e21", x"afef5871983e2b44", x"86b6b1ab45cba382", x"3f62d1c65484dc71", x"bf448ee1b852fead", x"1b05bc75e63fbe80", x"8d542c7477c3748f", x"5675ba3bb0cd64ca");
            when 7633190 => data <= (x"c81a4f910a6f7217", x"66b11d9bace914aa", x"ce13737cb2c90130", x"066402742e2328d7", x"81a4a213a3a11182", x"e2a3b3177e4d825d", x"4df56644394a5e78", x"1363b2820a318699");
            when 2188445 => data <= (x"b91737132b5dff37", x"e11e96a3cde52206", x"2d6a6a95d5844097", x"78c700facf5b2528", x"5e632f70b80e617a", x"dc1302966715feaa", x"4c510e0e3164d4e9", x"d2c6030a23c22aae");
            when 10905226 => data <= (x"3745f16d2685c141", x"c5450d6ff85001c6", x"bad4c04cf9105e47", x"354345b77dde82c1", x"6fe2c1380a3abe90", x"2b02bb51db878907", x"17daa0d4a3f72a70", x"635c35a57cd36257");
            when 25374332 => data <= (x"1cf130c1a1c94fdb", x"611aeafb1b7cb8f6", x"c1736b127f18c0e1", x"81a288e96a8fb8ed", x"402795dbb7a97005", x"c80d262fabab0b3e", x"59d4883e7377f4c8", x"0abfb2ae541dda28");
            when 21478701 => data <= (x"7239421cf39b2b47", x"208b6b6f43ed4bbc", x"e04dab627ba1a66c", x"ba449406160adf96", x"641d8b45e049ab60", x"b18465449fbc4109", x"fd364e890522e9ae", x"9ede2fc01990da9b");
            when 30950623 => data <= (x"bdeec82c7091ec1a", x"c57fb1d90d5e1cc2", x"df272b97499908e3", x"65132b904e2dde63", x"593d7a3554825203", x"20d92e151d79904c", x"4975bc3e32d75609", x"c8d6edada15a4dc6");
            when 15894854 => data <= (x"0209e17b60729323", x"f961b6dd479dc76b", x"4f5e0537665e161a", x"8b28bff6d17c30c8", x"9b6581d53a5c49b6", x"c6810a84042c1cc3", x"6265ea09dbc6db79", x"3cd7a812f03548ff");
            when 19723224 => data <= (x"12a19113b6638d9c", x"f10089536d05d319", x"5f0c93a0748b086c", x"6f7545bc297ac04f", x"9ff4ac2d35701b57", x"2764b2c35515c84f", x"31e774bc5e383ecf", x"3c55905873545d77");
            when 10918643 => data <= (x"ad20be45e0c5590a", x"5e46fe74617114e3", x"aab6bc735f5cadd0", x"19dee982cbe0620d", x"067a5add3fe1862f", x"d75f3622ac484049", x"54dca38df6f7058a", x"678a558da9b0155a");
            when 6729999 => data <= (x"63449c7641d1b415", x"43cd5a8d881e3139", x"a14883b04dc230c7", x"30b4326482c9a810", x"3ef29cecf7492f56", x"d4e0fecbc56c5dab", x"d169b2eef94d6a9a", x"e8b8b70f98033618");
            when 26149035 => data <= (x"7e2fa9e3767d1095", x"66a70839cdcfe7e2", x"434760a26f7ddbff", x"f72d5e75028f803a", x"0f3753f927546e53", x"92ef18fc0d84a276", x"03e09a29b24263e9", x"0673b1482476ece3");
            when 1157202 => data <= (x"cd94968bee046958", x"2464bb7e0417393e", x"15c2c53d9a4cf4b0", x"671f0fdf44c07108", x"bc5447b6ba6c5ddb", x"156330f1d43c569a", x"479496cf429a121e", x"508b744f395de413");
            when 14651229 => data <= (x"23fcf11a3e24002d", x"da2e12a3b65f79d5", x"e80da1a7f1cb7698", x"1c771a92251b0f66", x"168f0ac26ff51ed9", x"259042c10a70a2ae", x"e39fccead3fd763a", x"a30cd67895605e94");
            when 20170261 => data <= (x"d70b75fdff30f10a", x"aa92a1bb189e7107", x"a82939cfc5f9884a", x"911284e1ab4d48f4", x"a58b500cd1c04af8", x"ee5914f362eab7e9", x"ceb8dd2088130460", x"65ef29ada99e4c50");
            when 16883929 => data <= (x"2f22f6834861bcdf", x"67d23c73d395817a", x"6297b5a03df80c27", x"d04578d88ead620a", x"a7caf0762e57178e", x"52e37a6e59b092e1", x"4afaa3fe052c9f42", x"b648aa3ced1dc34a");
            when 31670103 => data <= (x"a65136dedc28759a", x"c3bb10a25662d4f6", x"dc27a35d61733571", x"3a5bc0c4e0bca5d7", x"f7bed44b67c0bd14", x"ddedbe1a7e88a7e8", x"c4ee05996c43762e", x"5cc1245fc18c505b");
            when 29697105 => data <= (x"9a14374be90bee46", x"44fedfab81bb4721", x"d720a516eed594a8", x"eca9c2833acf9191", x"5f96eaefb4dd7f30", x"70d6916e4cff9577", x"44555a1cf7d1ba91", x"cefb085818d26b9b");
            when 9403454 => data <= (x"b51db536841be37d", x"0b8651727b5d777d", x"68213a9c832effab", x"c54174efad967cfc", x"f449e08899952039", x"8775871b4a38d1d2", x"b0ce5cb10bc3048b", x"241d623714af3113");
            when 11699096 => data <= (x"94bc2b40b339341c", x"acc11e73f33a9e70", x"12c84260269f97c1", x"a5ee21a29cbf77e0", x"08bc7829834cdcdb", x"ba825622b0e28f17", x"49eaa1e5c0bd95df", x"007b4c2513ceb49f");
            when 14259126 => data <= (x"2510f2329318f674", x"2a658bbc0437e1a5", x"2a183cf8d4a0cb4c", x"5727c03310162563", x"6a17b700d4ffb103", x"45d1b19df6335aa6", x"ac76cc6be997b72d", x"6384abebab1f13aa");
            when 393161 => data <= (x"ec8bc6003be6f865", x"21ff062d674cc075", x"2622b516e6f43eda", x"56f159555506f972", x"daccdf4fca7b2eba", x"0e0fcaa3d2dec137", x"dc430d30c18d66b3", x"de90a7a8f99548f5");
            when 24547971 => data <= (x"ca4e75b862e59edc", x"a37bf5970888aaba", x"788813ddcdef056a", x"6133c9e36d28bba4", x"7e34bad10b28f123", x"56a995b9d9750563", x"81bf97c03423acc9", x"07aea9a66cd12e17");
            when 10801287 => data <= (x"8a35de2125e6b806", x"b2c28e21454c2eec", x"2c54d33a607ee6b4", x"9b4f88a6bc8f57f7", x"422d6f4166e444be", x"bd7441648d9d6f9e", x"9afe3d2894710e12", x"dade3f0abd90bec8");
            when 17883851 => data <= (x"9cd90fa4884b6113", x"1008ce684eaf6cb5", x"d861ba4a0b57ba5c", x"cd6737bc2270ecfe", x"08c2064fef4462cc", x"96ffadf08fc97d23", x"52cf0a8dd259ecea", x"5cb8c1122b013cda");
            when 26301911 => data <= (x"722ffd55b3c6822f", x"d4ba806326e00f18", x"70815c2a24399ad5", x"b3442a7b4b2ccb11", x"d6617a972390dce1", x"a0b04c5d15085362", x"4fce4a3ab782fca8", x"4dd366270ef63dbf");
            when 4478210 => data <= (x"28d25134c8d6be7b", x"dc33bd244841d058", x"e2141f34e836a92a", x"be6bdec665cdc97f", x"093703d75110b971", x"e1322117f75e3777", x"cb91b37e0c61a0d5", x"bab84ab712ba7de5");
            when 20855804 => data <= (x"67962851ec530f5a", x"3858029702c29a81", x"1af64de2ca13411f", x"555864627a315d94", x"0cd2e404445fc900", x"736ad48bbe1f65bc", x"aaffaa894113bea8", x"7195fb60327f9899");
            when 28315006 => data <= (x"affd2650aa34c480", x"eef3a3f25054435e", x"0ecae645802f6668", x"444b48666639b4e7", x"8cdb761f7ae46b8b", x"7613123915084195", x"42bd40ae0173e6c3", x"11b85314625f9666");
            when 2356944 => data <= (x"2dd35948f8f400a0", x"c479fc4b73f1671b", x"942ade2fe5a54ae5", x"e320c479b87366c7", x"9e420a1b2e053553", x"9cbae6320b7ce9e1", x"843193681a02286a", x"29fdb7c1743c0f8e");
            when 25606404 => data <= (x"f0020384cc288a72", x"5cced4ec6af40c04", x"a129a0e6a0dbe824", x"965f843a0169b2dd", x"0c1ba5353aac8c66", x"85ec91b72435ee1e", x"2199a61efa5116c5", x"5929984c2ced63bb");
            when 22015209 => data <= (x"44a972ee0c1d16ee", x"4d9cf516d46aad1e", x"98c4706dc9638268", x"3ba9206b284d278d", x"44ceb34b12f44a21", x"f7c5893e2883b072", x"4d76986aa4805c73", x"3e16564045c3b7dd");
            when 12974711 => data <= (x"b0558f474c640aea", x"2c77a1ccb895e488", x"0f63cac5c56d12cc", x"d89c45cf4f00ca75", x"a1b2afba013badef", x"8efa80142945d5b8", x"677e59ec2af6d80b", x"e8f37fee91354dd2");
            when 21991356 => data <= (x"3426a904e166363a", x"c19d1f4b67af8c16", x"958f64c00cf282c9", x"4b2f794f134243b7", x"261deb5d5f219e20", x"3bf35e802c0937a4", x"ad647353667efb73", x"abcc7af664b8a9a1");
            when 1014061 => data <= (x"9250c1801421abe9", x"f8be44dd2a873f7c", x"38daa70770f4a888", x"787052175eca4915", x"6d105cc42f221d91", x"d80a20db870378f4", x"76c3e8633c51441d", x"d67786b7933587c6");
            when 8145796 => data <= (x"293d96ea062596b0", x"5f5ef394a87ee60c", x"77328f0d099578bf", x"3b216b19c2c7e7ad", x"dbf0866afdfcd801", x"b25ffa353362d54f", x"9aa7f71c5b7b7351", x"33b557270aa263f8");
            when 4802343 => data <= (x"e0204e2c5ccd90c3", x"96ab637a053bad39", x"fbcf5490fe7ac3b1", x"82ce478f62fafe0b", x"6240d71f9c869537", x"21bf4a222545d065", x"c7074c74cd7277aa", x"5450ff96d46e2f8c");
            when 19336308 => data <= (x"a3f80f9601e7434b", x"f8253746f5be2bae", x"d6c0476d522f7cb3", x"2fad471e6cc3cb7d", x"0335cbcc1bc29f62", x"f1f499b85b696f68", x"e6effaa19969ed4b", x"9984fa99454923d2");
            when 5069668 => data <= (x"77188deb3f1edfad", x"0326966465e92e4a", x"8c25d6cae0fbc791", x"60bc5b74b97b06fe", x"025b128e53653aa2", x"a1b672b86145ba01", x"ce67d23f5c43374a", x"ad34785c9cdc90dd");
            when 28184733 => data <= (x"82c8d8da14fd1e76", x"6021f8ca94a6a627", x"3d80e6dda48a6ead", x"25ba34307287ae20", x"5eb7c0cd6c4874c4", x"361229592a83118a", x"3c502c9866d7f6a3", x"bb60bac43f971116");
            when 8255352 => data <= (x"d3e0bdf511e5832d", x"6cd02501e6c3aaff", x"45078a65624b1108", x"bef945cd4342a7e0", x"122d86845c667e00", x"7e14899431766634", x"e3e8f4077c54272c", x"1c9b167977a73439");
            when 21630558 => data <= (x"2ca8428395acd831", x"fbc5316cb9221074", x"61e3e77e2b90cfc6", x"bdc18ca258a45351", x"d4e4c32a4aab5050", x"c956c5ba2e46b554", x"e669feaaa96809d4", x"aafd3e397e5abc75");
            when 7036298 => data <= (x"9e79232b53c4cc98", x"78643b4e470e4af6", x"baef7d9ec47694a2", x"ddb105e3175bdaa9", x"1c66beddfb903192", x"e1cf6dbb0967c14b", x"e447646e91dff8cd", x"c790b1d2c698d26a");
            when 30699866 => data <= (x"47a9b1873f879b8e", x"bdc828c4e6b86eaf", x"ff1cf584ce292aa7", x"79e6a2521152ac04", x"6156df9b2e8776c5", x"5a886164aae743bf", x"dd1ed58cd9e58976", x"3b18aa6edbf24afd");
            when 453396 => data <= (x"5c4b423590c1ea15", x"668042b217d78e38", x"ef162376dbd93bf1", x"fa5f393ad9066f54", x"d29333132c0c337f", x"aa41bc4c73a57086", x"1837b51a95b2f4a1", x"274a24bb54a05ebe");
            when 8916153 => data <= (x"b53e8e1a383f5520", x"b5751b9f42ed9a35", x"4443a7909f923b40", x"9ffb99ad0cc53cb4", x"e0f076576a381216", x"5a8f4a100b8bcf30", x"43509262b9b62d7d", x"9bfbeb532352c0b4");
            when 14485032 => data <= (x"9ed73974fb58b75f", x"9b38de3a76519b32", x"e27a515b1fac0048", x"cdec86a96523b731", x"923faacaa5adacd2", x"68ab74c9999b308b", x"f2bb872d5679f38a", x"ce8e3e093a09014c");
            when 21622553 => data <= (x"718432390697b417", x"01a1d32e0f9fb03d", x"848dc911e4c71072", x"3a8d8ddd2a940ac5", x"0788861eb941d16d", x"162f7514b6df698d", x"7b8b9145ab818a40", x"c589206b61a81782");
            when 13316337 => data <= (x"a4758fa16c215ea9", x"743da6ed84cc3483", x"7c4aced6c322a755", x"041ef8b4b4ec6328", x"5788b22acefaa54b", x"682da367d71db2cb", x"0084cf30d61d3bba", x"cf7f3db68d34ff37");
            when 10578861 => data <= (x"6ad6e97500231703", x"bf892d59a183b95d", x"8e5608ecc9925638", x"558a357a939ea41f", x"120fb9836856cae5", x"0829b1465c75e214", x"3dcf5a2016afe6fd", x"5e704e08735971f4");
            when 32086944 => data <= (x"751dbfa5e6e90a0b", x"ff24ec6d18b68034", x"564f74fc344a5d7e", x"f7ddc1fae39438c1", x"094b54917ce9c486", x"8381c83ede5a7d1f", x"990b8a44eb4630f9", x"239e9ca1fbd73cf8");
            when 25511937 => data <= (x"bdaa8ac8176c0960", x"8308faf5a6621022", x"941dc58878ec3ff4", x"f63855415e9fd0de", x"13cdb0c9128db89f", x"fba0ace9ed859296", x"8e5571f242ff9546", x"3b726512d41d0b48");
            when 29503318 => data <= (x"0e63b38fc00ecd8f", x"c1607bec06ffd63c", x"54a6ff882ed7ccfe", x"5836e19b4404cd6f", x"6cecf18ea6417661", x"fc2fcf41b780aca2", x"31f6cffb2fddbf26", x"8f5767cb5dfd9e69");
            when 2364586 => data <= (x"1d29992ecc6b7b68", x"1cd589c8c6480dd8", x"bd77675a55bd6e0e", x"b985b717a078c670", x"12851e914dbc8f8f", x"9428aa823034985d", x"b687cdaa91fed4bb", x"8c49d04813bfbc26");
            when 26026260 => data <= (x"728f29fea85f05f3", x"bd71c86624e591aa", x"70f3e6d465f7250d", x"340db9ef19cef007", x"295187b693988f8d", x"f6e2ecfe6a6e6a16", x"87500c01a7df81e8", x"598c6f5d53478bd8");
            when 27799595 => data <= (x"f3d578b06045cf8f", x"880e2e3a77bf5214", x"86e1e382f1430f98", x"e67319b07883d857", x"84411f57163b50c1", x"a6cf8bb607832124", x"e15070cf952fd2dc", x"bb79449dae956332");
            when 1656772 => data <= (x"618ad216bd95db66", x"5e76cf37bba47593", x"4ec4502d00f1ab73", x"8bf9b04c95a1e7db", x"46e71a6b2a6a64a9", x"e661372a170f9472", x"76cd49ffe28c4a08", x"9f9ca40a29f3e5d4");
            when 30117951 => data <= (x"3c43701118ca2c53", x"793bf834ebff0067", x"7fb015cabca63a42", x"79556564b16fd899", x"313892538e24ba21", x"5b7ba224feff1078", x"f1407bcbb8eee86f", x"b5eab4eb19c55823");
            when 5650633 => data <= (x"95527fc8c54b0cb4", x"bd2eec68346bca74", x"94bdbac39024399b", x"babb039f4698a9c7", x"68becd7cbd053b79", x"943f1b0c80d7b9d6", x"61772021a1da7332", x"7565087cc7f4d405");
            when 6858786 => data <= (x"84b76b3a33435763", x"f68ac5157b106da6", x"9e694477ec53d7d9", x"8d7456db2a27e147", x"09304fc65025a49f", x"d2cb840522e201fe", x"104cb597d3908a8f", x"8e2ff9978022c9d9");
            when 3864950 => data <= (x"4ffc9ab5b7fd65c0", x"9ce6e17266820058", x"9cbd998ffa7b0e4c", x"1b8b01e2b47a08ae", x"81f447f367af0e3d", x"e3564a5e01354ca4", x"8fd44f79361d90a6", x"deff24bff06978a5");
            when 32921047 => data <= (x"05c9460ecd3c66cc", x"8985a53b63c9664d", x"bd1b6874e27dbfca", x"b9399448f6cfe006", x"795ec53ea827dd66", x"93d61cca43dc9d19", x"4fed9e6badf6c85c", x"4f936010a70699bd");
            when 26387286 => data <= (x"99af512f90f59302", x"1b660f0d131cd5ca", x"6a5cbba95d568e6c", x"876c30873d93e672", x"50d966d33b12147f", x"d965a382c92cb479", x"4259e75e0c2a0832", x"6509c0957a936934");
            when 9378699 => data <= (x"d659d7d5d3eaf744", x"9095d54d5c1f0487", x"03905b3f223ab9a4", x"58c5a82b8082f6eb", x"bc2a09fd71d20917", x"6cfdee0d3f13afff", x"b014231d05fcbb59", x"cbad4d74a74ab248");
            when 12229301 => data <= (x"bf256099d0edad09", x"7476a840c5214810", x"4f250dbf716f8ceb", x"7213fd7b00b60663", x"b8ef8448a691272c", x"0143e533f483163d", x"28d302dee5a5a323", x"2a697f22c1d975e8");
            when 32315529 => data <= (x"3de6c20bfc917f88", x"f9fcbe5c1bf264cc", x"1d81d6cefa85e4ef", x"92df9254a59153df", x"eb1cfb56759687aa", x"958b06c17175e3a9", x"553d19e806713626", x"c8831cfef76c6d4b");
            when 10611788 => data <= (x"3ec1866f2d7539c2", x"e537410fead41c25", x"000d038ce178ff0c", x"9af757635cda6e11", x"92c6337164e2298e", x"c9359392b0597660", x"bf3a0f91a4e15960", x"cd182cd9e29fe5cd");
            when 9587365 => data <= (x"a44cfea6d79a66f0", x"5fe4154ab826fd19", x"20ca550ae48881c5", x"7a18e302b96e0a08", x"12a55115f953b215", x"0ac5715f5381497f", x"b106047af581d457", x"efe42094ec1aa83a");
            when 5413357 => data <= (x"44e569bc93909f73", x"518a46463e9176fe", x"ab322d08265e7e1b", x"9df3b491b388bfd0", x"95f35338e822a750", x"6de91048124cea59", x"730c7bd3f01348fe", x"117d1c84b95e1b44");
            when 23773908 => data <= (x"1c6838155fcd5e15", x"39680140a4c70454", x"cd412829e7350605", x"af94247944c0d460", x"9ddf668c5c7c8bed", x"27d7a681a6f89d92", x"39f801223e9a851f", x"c5fdaa5d9cc906e1");
            when 28326603 => data <= (x"2a7e3058a44ec60e", x"7d01e19ba65024f8", x"8e35811658dd6acf", x"5e91ddaf45d814f6", x"a5848bc13e7b891b", x"542fc0e961a53005", x"a530ee2c7f791334", x"60e34b14ab88bfb0");
            when 13116282 => data <= (x"211ab540a3b24f01", x"fba84a777fe3f994", x"39e485fcad8d70cd", x"5312b36600d9ecdc", x"781c491ecea32539", x"cdbe72409597676c", x"92650525287f13b9", x"0a37c46e307352f7");
            when 8591856 => data <= (x"d0876ddca1422c0b", x"93ce800312b627a5", x"0e484c0b56eaaee2", x"726e28d908351d34", x"d799ac5cf1fa511e", x"9f134c62aab1b833", x"3654f6592fe9a86e", x"1eb40e1798f96d4c");
            when 33142079 => data <= (x"944186c34b0d4d6c", x"10cb7020f8e2b0e7", x"58cb847f09e539e0", x"33e62bd8ad224cad", x"27b86a90e7019c12", x"7cd049483895bf5b", x"9f549a96d9d3aaa8", x"5612a5a3409ff57c");
            when 1317678 => data <= (x"7d2ec1eeb2e935f0", x"c721a06f8fc57f4a", x"68c2b2dbeab3a218", x"73000be43166d508", x"c46dc07495a8982d", x"611a35990bccefc0", x"4274228d194ac2a4", x"853448f88a0f2c3f");
            when 10938313 => data <= (x"4bc8dedbbc29e381", x"2ae0296316950596", x"8511dc24101004b5", x"713f1ab67398908a", x"bc3393f1b3872d1a", x"147e99de0fc2fd44", x"defa3946a1b593d7", x"aff9d7e44b6d0c0a");
            when 3323249 => data <= (x"8c95e191292c1b9f", x"ad23f8e47d93073b", x"326e7ecf70d18461", x"51fc33321a7fdcda", x"63e63e6a12e118c6", x"08217a6b93062dea", x"fc379a25cba65253", x"ba62f6060fe6dd1d");
            when 14945254 => data <= (x"b319277a81bf2d61", x"64e4decc264d871f", x"769647c91df9c604", x"9094d7341d9bd63c", x"eee0bb447b35bd18", x"30d4d1936ab51b00", x"7b991a0ad3b170c9", x"847088a3ea0aa471");
            when 20517196 => data <= (x"205cb04dc53a1df8", x"f72929fd68490005", x"2c6bd30f9a5a6bb3", x"dd77da86ee1bb961", x"6ca735b1ec64acba", x"383f55bd3acf9a8a", x"5426cce3408bc6e4", x"1de1f16719833aab");
            when 8503493 => data <= (x"1c29434962d2e794", x"87768384f1f17b26", x"26c99d3733a6cb93", x"29a1491237ca8c50", x"a3cb5fca976d5602", x"f23d362cb5d3d78b", x"281f2438feba2b10", x"ccd956542f2dc688");
            when 11963029 => data <= (x"26157b52dee35bf5", x"ded05277235a9dab", x"6605ae699c6ed294", x"6a1a4f646a74c7fb", x"75a94dc1ae9ec31c", x"040ac89edb6be23c", x"aedf83f0a0f84d3b", x"0c27756805326eb1");
            when 30852347 => data <= (x"6cd8e1f247d341f8", x"ee4b2d66ac855cdc", x"fe3e904981c94518", x"cfdfddeefdcedd0d", x"06fabc5880a85ea7", x"ddf2b37bc9da0e05", x"5391137490a3ff2a", x"838b6453ee008792");
            when 15202408 => data <= (x"1f1940fa3e739656", x"8647c606c909e5f2", x"6cb1754a2bbc66db", x"756f65d5a340d2f2", x"6d800844bf767f3d", x"b3ff32ed62038475", x"a0eae3171f4c3dce", x"fcb2a2336e1024fc");
            when 17054359 => data <= (x"1b32616fe7bc320a", x"6a4804d88631047c", x"a1c65daccb66bc94", x"819124339e4feadd", x"bc904f6cf33551c2", x"b14afa990642e5e8", x"7e19b052c43b451f", x"8daf78a45f28b215");
            when 32686087 => data <= (x"90c4e0b48a39beaa", x"84cdab682e73c691", x"690bfc655e2b0e66", x"3de4ad69443cd5ee", x"a86fd9a5aa278e78", x"9509b0faada501f9", x"4221be64e65fb59d", x"1df8f97253619bdd");
            when 9586325 => data <= (x"97237ea868624c7c", x"6c13ca32b9aec39a", x"d83422b921840d89", x"651aad3aa1af0a12", x"9992ba0e4a7771f4", x"d399b6936c015583", x"94479fdf99ec3df7", x"2c22197a7787e6f2");
            when 7607215 => data <= (x"058402cbd29f76bf", x"ebdff4bbf968191f", x"7fc362ee47ed7c17", x"83b341b2602171fe", x"6d84f88291ecc9a4", x"2060fe5e49e38e93", x"73025d46a31332f5", x"9a013dc8703f1f4c");
            when 11411279 => data <= (x"13aca322f76e7534", x"5b6da8e4adec86b0", x"f51f70868c9ab545", x"cfa3bddca8bae0db", x"82345f940f02197a", x"7d06016feba81375", x"f9af992c52c523db", x"c34e10e9bddcd927");
            when 33346987 => data <= (x"d66c50ba6f6cf672", x"09b8c33d9809c5e4", x"b89c285555c1e71b", x"07982a1abae2108b", x"24e4af36eeac0472", x"a4873116adfa73b3", x"b6e7a3baf17a8689", x"14a40b5a542535f3");
            when 3735467 => data <= (x"cca2612b62d3f0f0", x"58fdc1eaac8f8223", x"50544d8f73666ac0", x"7f14843f2ec026e6", x"3c0f58af926b13cc", x"c90984be38e889aa", x"8f45306d34f9019f", x"49017032d9f208df");
            when 8361890 => data <= (x"4e7492656e961408", x"446ea0b55b54a33e", x"1b163833c7129762", x"34fc127b0d492cde", x"4e0d2d804e04d479", x"5f8b47a6f4f91e01", x"7901a1d0898b0ff2", x"1ddae6f6b778cb96");
            when 30424682 => data <= (x"623bd1a4efe380e4", x"bd8eb013198c162e", x"2dae2bfa7a410045", x"8ad17d7d35dcc0e8", x"1d12e73485f9e7fa", x"00a54485f4fea29e", x"3073bace2923ae1c", x"9fc30a4020527e26");
            when 6494551 => data <= (x"1c5ac25875291a65", x"2de025276e802d27", x"57f6062c45ce9c2c", x"7aced53f6f30b23a", x"75aab8a9f555208e", x"2e1b7d21b69f88fa", x"bec17e00c6521260", x"df54e50e5d08ebbd");
            when 2658201 => data <= (x"c3e64426d40ab4eb", x"adefb1e698c6426d", x"310326fe80937dcf", x"09dddabed6a32598", x"14a9d703c8849cfb", x"1f75cc9052f40871", x"3537228ef5423ca3", x"9b03d220a6648385");
            when 16771563 => data <= (x"a9b3964f85cc9736", x"205dff733940971c", x"df564f75f8bc3751", x"fa432f5f2618e7e5", x"52ae55afee34cff5", x"a87f203d4a48d8c2", x"e64a2638ccc10afe", x"68d130313d86d861");
            when 15443667 => data <= (x"f6b6fb2ee4168626", x"f946e4e62c79045a", x"c52faa9480ef0682", x"401a9492a2c406f5", x"f36ce2ea4780c1fd", x"16ef64adec57ea5c", x"9e31cf0839fd1075", x"4d4d4214fa531994");
            when 26326077 => data <= (x"1f03946d2ff9d728", x"645ac102f9ebe10c", x"21f5e52d4306ee7c", x"b5d457a18eefe424", x"7608a322347a3d7a", x"58648f95d07b5272", x"e95a15e9bca54954", x"daca595837143226");
            when 16387052 => data <= (x"3f2637dfc7e3973e", x"e59fa0765378673c", x"93f737565c86c7c6", x"aec0b6b2515ab9e7", x"4524c5f367a85d7b", x"8e6b84dc585c6a39", x"b39fd34f1706a5a8", x"46576bed325c8cf7");
            when 11360311 => data <= (x"e20c2f973a90ee61", x"72acdfeb072d1663", x"84b2f89d2f354c5e", x"8765895da1b2c335", x"e6c223f0fe5f2fb1", x"c93583f3467ec656", x"2ee70316ff3f5d23", x"99f8318f744ff6ce");
            when 33121857 => data <= (x"63e7054a7b070944", x"f80b1175c350ac67", x"de0914fbc70c44c4", x"ae3eb33672d0858a", x"8a7286ce989e2beb", x"e913cfc846983b2a", x"f0302137957576aa", x"2e9378ae60821959");
            when 8065521 => data <= (x"d6ebb884298c0e83", x"e7086f742ad46093", x"60973382e2604e8a", x"d4dfad1e47edc588", x"ab8d1a2f849389cb", x"d8d7bc4395d7384c", x"ec6e7d931df5869c", x"ad718386a88431eb");
            when 31800307 => data <= (x"8340f4c317e1b661", x"aa66bb3864185caa", x"a7f6a4ba244fc1e4", x"94580df4080229c1", x"49a36f44a8a12dc3", x"b5b8883be0cf525a", x"9a120be436efca8b", x"b8abad4d1cbf13f0");
            when 18188804 => data <= (x"703462de1b60755e", x"085a02853d719933", x"2a4b24a9659e0406", x"5ff0a843246c8326", x"9ede213fec799ab8", x"5b0223fbcbb2d303", x"25d17eaaa26d13a7", x"8f94c97ea4075d18");
            when 22996385 => data <= (x"eb8d155939b069b4", x"38f427316c0776c1", x"440403fce2688507", x"29fbc58285b96e16", x"6dd49dd520a0aa60", x"1b12334cd36e85e2", x"a85865dad4d47f50", x"7a667976b1c1928b");
            when 20459727 => data <= (x"9fea9805bf4b5581", x"5f51b1146a95aec7", x"4b746ccf107df9a9", x"174eeb2e835fbf86", x"ae2b12bed3aa8da7", x"e4e25f3cb184efd6", x"1e1436c84033c5d6", x"58c242f9212e4e75");
            when 2482084 => data <= (x"122ac21256a218b6", x"f2a580c92650550f", x"cd3cc7666ab119ab", x"d9a9fd08dd4d6986", x"68456ad7d90f4adc", x"fcd6783be0d4b55a", x"c3c0d45b2e61826c", x"457596ca06023ad6");
            when 5480524 => data <= (x"d7cb158694217acb", x"1ca478985f5a212c", x"056a46ea74b9edc8", x"3dcb29d29d7b6bf7", x"2f063dcfc17bcf1b", x"2a0bbe91da10d7f6", x"24bc05bfe6b43e72", x"0303341e69215454");
            when 2288922 => data <= (x"48e28627de3d1792", x"2bd458a346f0f6a6", x"ab998a11bb68464a", x"b353bc4f0f4bda37", x"bd584d40de49f77f", x"502dc76524babe1d", x"966b12505da7c8c2", x"740b5b277ec8c299");
            when 33155998 => data <= (x"de2e306eff17a2e6", x"349116ad7b230aae", x"169792197b5e3b2a", x"f2f5a5940ad52ca8", x"8b0d00a0b03faf13", x"761d5c457f9de4cb", x"5acedcc598ed6cd9", x"2f6b0e4f250ef7e4");
            when 33117639 => data <= (x"2bb6637df88abb91", x"46821a8f33ba165b", x"55b0d7ae62d560c8", x"3ba3dadd610ceb82", x"87fa5a0378a9f003", x"54967af793c58795", x"9b558134859a4dba", x"3b067f914620651e");
            when 19781204 => data <= (x"7ffbc8ac5aae555a", x"e7e53138ee8aac87", x"032f6c8f8636c281", x"389aefb1bedf0ccc", x"626a8823294a3950", x"84060afab0231964", x"1496c145fbf9faf5", x"0279c483507861f9");
            when 14147138 => data <= (x"08cc9208d67d167a", x"180705fcc0b1cdfa", x"fa481a0117570950", x"da7be00c28b40f69", x"3d065e7b3a868c4a", x"ceaa506417f23bd3", x"9cb6ccc5a4712c39", x"5e63850251cce985");
            when 16297583 => data <= (x"1cd8509f1a81b21b", x"33d46db3a328c836", x"c73d044228642fa5", x"dca3082420fcfef0", x"27bccbfc9259f3eb", x"df096fc9001150bb", x"9d816008e378ff09", x"eafe34d7810dc2ea");
            when 26815022 => data <= (x"476644ac36cda0a5", x"09dc57b5fad46efc", x"696e4b9a3fcdd6de", x"bb532cfbeac32f03", x"6490aa990dda2a03", x"6304cf8bd5269b81", x"1fa11986140e81bc", x"7af854b6621b90bf");
            when 8362817 => data <= (x"46f148d853d91ff9", x"6ff53d7a542b85ee", x"74c212de4c31ee16", x"017daecda64d7a1f", x"e9f6b4cb296f6d15", x"db098346ee5a4509", x"94ed90e117808b5b", x"d1d2fa1288c4ce7f");
            when 22981595 => data <= (x"009291af0f783bd8", x"64244c9181474d89", x"a296c767e9159e21", x"b9d34d6e6e811561", x"a7015354bf1c25d6", x"7eed3d66178dabdb", x"6a416df24522273d", x"97a8f2fc321f174d");
            when 2320892 => data <= (x"b23267b9c7c1cf5a", x"7916034016b67cf3", x"736082baeb4a1159", x"98fea051278bce3d", x"db531d6460050f73", x"60c933b94bd3d2b2", x"a62d46d74548e3b9", x"2be20b7caf0e3846");
            when 29521205 => data <= (x"16a1a49e527c837b", x"a8b85c01624f2184", x"629c0fa8fea9518f", x"65ccb773ebc2f120", x"1ee94436c198c034", x"19210579e897471b", x"086d22da43de84cb", x"bf7629e94da3e896");
            when 16813803 => data <= (x"3c47dcbd3be04008", x"362ab9295ea5415e", x"1d59b4b3488177ef", x"877965c06046fb95", x"e3f7a0144967bbd2", x"39fbcc3a677d02d4", x"1bf40b0073419fe7", x"2f765021d4f0b690");
            when 22964834 => data <= (x"a1df505a0cf169b1", x"5708f84a37ec4f32", x"1731a6daa2f44e97", x"653cba3bac7adee6", x"b3e10d79e748e87a", x"4263cf272881e3b4", x"7f504a53ad9e3069", x"3fa81fc222e8f4fd");
            when 16022983 => data <= (x"bbbde43eaa7eef84", x"541e5af4160c2543", x"2e16d53357d40b35", x"80e63bd8175c8d16", x"332bef7a3d240540", x"e366c099a0195663", x"8b8c6ad42c069259", x"9043502db87970a5");
            when 16040126 => data <= (x"3495fc970c92c9f3", x"ebd95346ae2d7907", x"5af675eba4649b3c", x"a8c8cc9ee26eb76b", x"fcf8f0bf13a70ab7", x"53524d9140f2e004", x"8e88ec9ecb5bac0f", x"5609d98e2adb58bc");
            when 9653726 => data <= (x"180ca78106666256", x"e7b3ec05f6d078d4", x"b51ceb06ac824699", x"18dbceaaed1ed31b", x"564d573f206ecb42", x"7f639b9c156431d8", x"32cd2e3fcc48fc6f", x"2d937e62547a0aca");
            when 13641049 => data <= (x"67111f2047190d2c", x"27b2acface859c6a", x"d78410df1691f654", x"98140f74e527d758", x"533379ee1023f735", x"1741880069037dad", x"72d51540cfbc2619", x"e14a156277da4b31");
            when 5447452 => data <= (x"f87c4a49c2524935", x"bd09a214c1c2809b", x"4fe19c818085c4c0", x"8d979840a656986a", x"4bcd769e988d3720", x"21c579d93effb422", x"f6a2c15b66ac2afe", x"f994762a4fa64719");
            when 14701049 => data <= (x"d80cb9477d3e6d1b", x"ba88a12375954960", x"0143f194554bfa13", x"f2aa863acdc2e89b", x"ae18be56dc9cfa0c", x"5b6436a1f050724b", x"7c03be45fbfcb25a", x"edf1c9f83b09bca8");
            when 32504986 => data <= (x"da8ab7ff95e7c1ba", x"0ee596f2d4914f14", x"7dee86eb18b1e61e", x"62cc2b93deff9c0d", x"1d4d5a140356835d", x"cce1363a94448691", x"d50f50395115250d", x"cae911363c2ac694");
            when 9581380 => data <= (x"e164f6d25f8e3ce0", x"7afa4568bd9be4e8", x"b97cf6b5e3d73674", x"a156358e7330b886", x"411f0d542035af86", x"41d8f9f6ffeda981", x"acd26f718022afd5", x"9d61eb915a2f7617");
            when 3176490 => data <= (x"3aaa3aea036233ce", x"5eada66fdcb82654", x"e3a8842e988ece92", x"7aa305960828a68b", x"8b106a14e68f3667", x"8d39e4ba492b2660", x"da51445da44522f2", x"40489615556d761b");
            when 4485992 => data <= (x"d11f4f1b1e4ac2ba", x"35675afcb65afe54", x"bf2c7e37c797166d", x"993e7e041d1443fb", x"d24996cbd33f072f", x"ddd6d03f62ef1cca", x"d7224febd4ab8a75", x"ef997ddf17b25a38");
            when 5868642 => data <= (x"7c6f95a38fb334bf", x"d5c5c9875100ac96", x"73c4c9e08793d213", x"82bb2342e5f46db4", x"398f69d883c039ee", x"6067eeef8668faa6", x"bb42da151e54e1c7", x"8b2b127a051a7706");
            when 30466970 => data <= (x"8d1e0c2fcee183a8", x"1668b667226fb984", x"519171f205a1c444", x"6912238d87435522", x"085156cb58a532db", x"47b8c28cf6c0ed52", x"e64711a9a7f0eb35", x"3fb4c2b382a15d4e");
            when 6069345 => data <= (x"ab32d06da4f806cc", x"edda4ff89d4b5b7f", x"2a51e6b8224a3578", x"71413f4425ba2a27", x"dd08ac30fada35d3", x"f8cf0883c15d07c5", x"608f327970e83b22", x"b7681c0393e667d5");
            when 22611203 => data <= (x"674c1a5c399529c6", x"cfd93e3fc8e3b92a", x"9c3eb7a60d0b9e9e", x"13e5df66ab0b179a", x"6511b2e886d9c6d8", x"86336482f66ad39f", x"51c81421301a4761", x"7329e684c7178960");
            when 11774802 => data <= (x"cb56cd6d94cf396c", x"e201e369cbfd0914", x"43cc5d0d7b72fdec", x"8514993781c12233", x"018b36676cd854a7", x"be7a67a03dc99cdc", x"9574cf2d3f375eb8", x"e67bb2b37c4d04ed");
            when 32962034 => data <= (x"80f766886da6c2b8", x"bbec96a1f058bc63", x"4cae6fd097f4e47a", x"ecbb493b1e94abfe", x"0043fd99b617f5bb", x"d6c047b92ff6b9cd", x"42a624913dfda6d9", x"1a6d13fcde4b2fc8");
            when 31950585 => data <= (x"e60e7c9bd41e4b06", x"a839944331e88b47", x"b56e6b20f4bd5f55", x"1127ba894b7d6483", x"5525ed99c0b1f755", x"381660ff87c5274a", x"07c09d9d1ee38215", x"4bd3a5f1fb71537b");
            when 5355154 => data <= (x"b6691c24312b4b7b", x"c0a32d401a94e4f0", x"29e6a9fc088c28c4", x"bd2f9266c77b5998", x"29ecbe5e596ffd82", x"59468e9559ba2551", x"28015150d5a197d6", x"a51517f320e39aa7");
            when 15364803 => data <= (x"7b89486ff73becd5", x"26e6288fcde2ff4f", x"ef5ce3627ccdbd16", x"77eb978760e65709", x"2b7f9c3d3d912a1b", x"d8327c020ad02d85", x"f5bd9f4b8e87f4a4", x"edef08243b486ad3");
            when 6953616 => data <= (x"18ff37f5e1f700d8", x"3f4835f2d6a69266", x"a8641f2d676646e8", x"f9c0e07b2bb13be0", x"de6b3da4094543c3", x"f67ed4062113fe82", x"3a24c927179c36de", x"c12f047585123162");
            when 14165330 => data <= (x"451a97c46b4e6534", x"144e41e34bbe6f4e", x"5f598e8b24fe2e01", x"dc2baca6655c13ab", x"d023eaff6acb37e5", x"ce089542088c02f2", x"3aaa14346ccafe50", x"313367ed3d70857b");
            when 25866300 => data <= (x"b028cda5a939df5c", x"dce5c6d42b4e96ae", x"8753151c000b04a9", x"0f44cbe1cde49628", x"f8936d55848f97e9", x"295820af6606045c", x"18e6ca49bfc6f210", x"a5b7f631b7d3b7ae");
            when 20747197 => data <= (x"787e054b34c8f483", x"5cc38c392d534b91", x"d10676c178ee1c78", x"46025d15dd5ed11c", x"62a0085fc3c7e705", x"ad4c985122edd199", x"151ee1606474e04a", x"c5f73d8c42d9750c");
            when 13002509 => data <= (x"f655d6da2e365100", x"589aebf154971567", x"c32321ca5cff3503", x"3b58821437b9063f", x"07607a3aa1475068", x"a6880ad70daf6bdc", x"77bcc2c86b809f8e", x"6feb23c71d8d790e");
            when 3061367 => data <= (x"59f436cac2dde775", x"77a78739afcff1e7", x"078f47e1959cff23", x"480f4d9aa4e5484a", x"05ab007388e14d99", x"4c4bf70523d0b58e", x"2e98eac5ef689763", x"0b3c5025ce99344f");
            when 26296192 => data <= (x"054489a5fb628066", x"2dc4be44d12cbd50", x"01d54c897df29f5a", x"039d35d802b570d7", x"b4c881778e0e362a", x"1e5cf002a2315a12", x"f6ed8ce6f4fd025d", x"111495a99128bda4");
            when 15305997 => data <= (x"46eebcbc2218eec8", x"880d790d4bbaa409", x"fab3a4fbb1f02208", x"29fc49f6791e5a2f", x"a0d1db09c2844723", x"9cac578cff605b26", x"d03b598745416b39", x"64b542915b230ba4");
            when 12961862 => data <= (x"071532b0c02ef0f5", x"44381668273ae552", x"f7d643793f7445e9", x"0b8181f3e24f0822", x"ec00849ffffe9de9", x"5045ef7abb9e2553", x"3ae4b1a80ba46a3f", x"1036711a225549cc");
            when 31520035 => data <= (x"5455359351abb507", x"b9a2fb65837b7496", x"a741a99b888ffb57", x"30a8515e633c05fc", x"6dddfca47ea136eb", x"53794f1e677d146a", x"76e59d45551dd026", x"529d4dc9be122e06");
            when 22294805 => data <= (x"fca7c55ae6a51292", x"f099117d6f37b13c", x"00a30e572f123cfa", x"733087f7b50d6c9a", x"0afd6074ab28ac88", x"033d763fb6978593", x"4d1bac6bc6d013c0", x"17d9974a567c99f9");
            when 9848320 => data <= (x"622a1dee3b4bdfb2", x"a82b019c9aa15e40", x"e4bb138aee64b880", x"54b7096d11bf0994", x"7a3e92358b1347ad", x"3abf9be9a83d656b", x"64b3e43f088218f7", x"f21f5b4aa67c0f63");
            when 14600222 => data <= (x"73209b5d47b2185c", x"0468acc4a063ec66", x"68d0894743dd9286", x"f61be02c8fed3b41", x"bb7db62fdfb08e60", x"f70d26e4f0918c79", x"56b7615a5c87521d", x"39056c6cfab6d199");
            when 22101125 => data <= (x"9c0ae43b6065c340", x"58d354938427a113", x"98e4954cb3723f26", x"32b3cc570cc67406", x"48b6a36a712705af", x"f45413c6048520c3", x"0a2d5388ead12150", x"57011c57c576c315");
            when 31529768 => data <= (x"900ed6604cf4fd43", x"64c200ee4227c83e", x"bded95a0d7ff30b8", x"3b59753458b2f42d", x"f56615456f10d93d", x"6d922876150c4090", x"032d81444cc5bd77", x"6411e92d4b8216e3");
            when 8745971 => data <= (x"8e0246b69ae45bc3", x"2c44ecf1e8b065ec", x"f8c3b9ab143829d2", x"43b7a1c8efac3ca1", x"ea37aa7f779230c9", x"bff571c130a28f08", x"0e72bded1d7d9872", x"cc87b58a2e49244b");
            when 30570972 => data <= (x"5ba94094f7082043", x"e46a77e04d6d8061", x"a98d8e57376694c8", x"a01aa83bdbb73f58", x"0e8a27296c0ca155", x"8bbfcd2a8be0d3d3", x"8429d1159583805f", x"28d08099f6273c4e");
            when 18720844 => data <= (x"01776623798efda4", x"b49d2b25af244377", x"1dd49528a0bc06e1", x"b5728922815c12b5", x"1cc564d9a66455a6", x"b2243760c2786ce7", x"21b91b4394cd621f", x"6f28e169b0a0b96f");
            when 18893968 => data <= (x"9f89825f24863dc6", x"63cbf1ec9871eee1", x"908e3ca67f6ccf91", x"3e837c8a500a1b3e", x"ad70f674ed2aa312", x"56ba58fc606d1b79", x"3058039eb276097f", x"69a9d49f000a4486");
            when 32203846 => data <= (x"02bb31994a56b66c", x"f2961791e25c85b7", x"bcd4652f7ef26b8b", x"665baed68fef3f86", x"c43edfb5dd56ffcd", x"f7a0b5ac9dd6f365", x"f662e5841d6f18c9", x"ddfff4c83f6e5516");
            when 18684949 => data <= (x"bf0c10d5d85d9c6a", x"d963211ffaad70c1", x"92ad5027753500b7", x"b61f0463cc67b2be", x"b9d3bf5df6c65cf1", x"bd3bda1e1cf6dfb5", x"9f0805b37338f113", x"3a18f8d7f345bd44");
            when 22685278 => data <= (x"2c990e30c973f811", x"649f8e6a49e40137", x"97309f01dd6b8007", x"1ea0f85cd92c1325", x"57df3eb27d481a1d", x"80fe342783ea75ac", x"149037c99d09874c", x"17c943fdc67b3a13");
            when 19023833 => data <= (x"f5733d8955c61279", x"615f2b5c5d49c5cc", x"dd35f117fdb51d64", x"1ba124371ff5b80c", x"419a7144891663dc", x"1f69d24c24b88d13", x"c4c4904d8ca64ffa", x"a9172116e1dc5496");
            when 25205909 => data <= (x"9cf74d6cee3c5d3c", x"96e20058ae06bb8d", x"6869d9ffaddaaa1b", x"a05dc7fa94efe52d", x"18f1346a3da36148", x"813fb174a506c289", x"b49fb681e25ba540", x"a4ffbc4adfa862f7");
            when 18665875 => data <= (x"8c9d82d26b8ec8b8", x"e72024b54eb4d0b5", x"186b35fbbdf07de6", x"1885967d1f053d3c", x"f41d3ae6f2c3b65a", x"e3cb3ca6bdda85c2", x"86c9a032e62aac10", x"900d0a3317cfd6b0");
            when 10231775 => data <= (x"631f43c8b5631f5a", x"e6a1f789e7a451db", x"0a326b285457583d", x"f67a31b2da06ebb5", x"598cb681ad2966c6", x"6497135cc98367ef", x"b474e065e43351e3", x"2726eb48ee418972");
            when 16877471 => data <= (x"6a3733b90c4964e5", x"b882f25002af090a", x"adbdfd64bde236d9", x"124d1da676a2a5d9", x"848507cac1a672c1", x"d7dd6d5a40f312da", x"231b365c72fab677", x"d3ee19b429628414");
            when 4862601 => data <= (x"9b7d01afdcd4fdfc", x"5cd5b51bdd960ac4", x"25125767bfb44601", x"1d057cf2f777b2a7", x"f967a0c20059603d", x"136b0329beed8041", x"0ffddbf100e010ff", x"e0da94fa0d6bf994");
            when 30129303 => data <= (x"bb11298c8eecee8f", x"0778298cf3099ace", x"ed93eb2a1ce9ecf1", x"9a4495f7487b062b", x"2c0ae59a8679df10", x"f4faaa822e3a82f0", x"e70b4ca0285daedd", x"52b199ba2c0fe383");
            when 24219960 => data <= (x"332c236c88c1bd44", x"705ed2e339118ef6", x"b79b1e7146590078", x"6eaa2d0c5f30c18c", x"f9cfaa3fc6bf3ccb", x"357092aaad5ca21b", x"8c5447b8f7af9b07", x"a22ea5e08d106ddb");
            when 9996271 => data <= (x"26b28e37b53512c3", x"76e08ab0d1d5c215", x"4c1d7f32fd0083eb", x"ff528f79574ad35b", x"0248deed41afd923", x"d86453b7c3611296", x"9902c24132ef629c", x"e6ee5cec01e01ef2");
            when 10191411 => data <= (x"9136206556c973f8", x"d2d94b0efc4b6c31", x"6d4bf375fde1d6dc", x"26cb41b12cca7252", x"2d30e166628ff27b", x"23152b421694cefb", x"b1f5be878890bae1", x"d9857b8a8402aafe");
            when 7690840 => data <= (x"77dd35ff78633de5", x"7dbf95ad93d55cac", x"d1c3ac0ab402afcb", x"3509c609f70e0c13", x"d45ded8eb10f9e1e", x"d837f449d127193c", x"3495fa2fbd239ca2", x"242f9f30df9938e2");
            when 8974409 => data <= (x"427860d428315e59", x"ee9d835236c3d16d", x"423d1773ec85641b", x"c49fe2b3aa596ee9", x"31a0b81e895961ce", x"c6eaef9807226eb3", x"755e723327a7882a", x"2f3d7fa581102ada");
            when 27261273 => data <= (x"8cf72aef8ad6116b", x"85b79a8c5c0ba7dd", x"20cffdd2a11f83ed", x"e1b870592f8fa271", x"72df67365f4b28e6", x"c3b7e9b70a303fa9", x"cae08a047b9e570e", x"fc3625cb74077393");
            when 33492912 => data <= (x"c0f71eb14a5d9b5b", x"95c84b1b412bd96b", x"93def8fde8cb3e3a", x"ef6d6b8b2bbfb86d", x"8b12cd549bf0e3f3", x"11a608c8cf81d1fe", x"1391ee047df9047b", x"91e65eada3b905be");
            when 10362194 => data <= (x"2c34925c0b0ab482", x"53a5d6cf299b37ae", x"7a24a9c940ce645d", x"3feef2d932a874e8", x"7b61c8200fe8176f", x"1495cb909f7762f6", x"8514b3ada930e286", x"07361f0015e98804");
            when 13133150 => data <= (x"4cf3e22fd9825c1c", x"92ac2161b52545ec", x"d1629295f0ea587a", x"5be4c3fb52f7f6a9", x"637d2a4b86e4e5f4", x"cf24329178b13889", x"52f97557755ed5a5", x"2021fd50092c0489");
            when 1208223 => data <= (x"5ba953091ba29fcc", x"848655a3840c6037", x"63af01bb52a8a826", x"6d67243e2d6d48dd", x"5b0a3f26010bb922", x"f339237fdf03daa8", x"957b1509fd2d9d51", x"489be0eb2280c1ef");
            when 19706156 => data <= (x"4845702e6ca3dee5", x"6d6d81493afb33dd", x"830f03b962dd7a99", x"3337e25a417f8a57", x"9871878d68a82d68", x"aebcccace74d77a5", x"116ca120e0ce330c", x"c2cdb74eb4dad4a4");
            when 18981856 => data <= (x"40fbca5fd9981b19", x"940a58a0f53bb458", x"7656232f2f17862c", x"640f3ac155159cbc", x"be2c8759969ae4e5", x"98b55491db833cb9", x"b35e2c5148af5988", x"2b7d18c6e63a1485");
            when 1301364 => data <= (x"4841428c2d8c88eb", x"4bbbf700e8ae686b", x"0016e2ddee25ad82", x"358a781dec90095a", x"87304e13e4879dd9", x"1ae714828629a537", x"6fbc93ef8290df67", x"a9db7be4504cce91");
            when 21857697 => data <= (x"9b8d257d80f8b4f4", x"dae87439725407fb", x"d6c3039a71fdd886", x"a8419f45f469b0f1", x"c0e9c497506554af", x"a9f3c67d62c56024", x"15f96a5ec833a30d", x"8812ed25c407475c");
            when 18945969 => data <= (x"77d2b5fb0fce1992", x"32115ed4379d572e", x"2ffaaa82d723334d", x"f010ca5248ee24cc", x"6c28bcde2ec8b282", x"38eacfd579eab2ef", x"973404cdb15ce1bb", x"87e0bed1d3058542");
            when 23702665 => data <= (x"b04d07443457d74f", x"cc7d514b49876e68", x"58bce780292bca8d", x"eade3403702b0f07", x"e8560a1c7e090889", x"50670e1a8b801f19", x"aca4a2b7169b9f71", x"905d92aff739a15c");
            when 10009419 => data <= (x"9c4285f05154177a", x"780d4a62c074605d", x"932fc26e4e9d5e23", x"214277270371f4ab", x"2d027d1afa61bad3", x"51307b0433568117", x"4fec1d7f581157b3", x"eef06a6136806c92");
            when 18160960 => data <= (x"5fee7be00c2b33c4", x"76113ad6172cc89a", x"8d9d4a2ab565ea3e", x"ef076da85c2a1cd4", x"af85c2dcb01d690b", x"f0cb29205452fa69", x"1141433f3c17ecdd", x"ecd13bf9db413f67");
            when 8834958 => data <= (x"84bcbfc7d4bf9ee7", x"cdd6dacb457c5eb8", x"1cebd50e6970c550", x"f7c238e27e3b241c", x"6f1960e7d21c6b2a", x"c72936f34b7eded8", x"9a8bcc5d462e3bfb", x"525ac195f18d52f1");
            when 23691034 => data <= (x"d26d132f57fe5150", x"671310960fa7d87b", x"dc3953e71942fbd3", x"d4ac045e4999084f", x"eda1ddeb98fdaad4", x"af6e7231cd13b17c", x"4d3d258922ae5c81", x"142bcd47d06156fe");
            when 6046082 => data <= (x"672f2606bbb6a030", x"2541bd78b6a27344", x"16e3b20db2d15ec1", x"2c39dfceeb736728", x"bb492acdadd7fe89", x"5bdebc63f4785b26", x"b996db0f737dc2aa", x"75008847a534b2a4");
            when 6549553 => data <= (x"1cbb225c0b1f3288", x"030f0cf660468b05", x"3b37ca290af34931", x"49336944034f6c62", x"3debe034100ffd08", x"2e109d200dea32a4", x"ff9f530bfec850ea", x"6015be903d675d59");
            when 18061991 => data <= (x"d3dda3e1f46eb988", x"3cfa06f855860d85", x"f712f66e5ebfe2c6", x"09c723b55f48f238", x"6307d0c2e0e32410", x"c1e720797905bcf3", x"3cc5b6e4c38a757f", x"7f1e79432b815fef");
            when 21882069 => data <= (x"eded8eded13db673", x"afc55cc7908bf2b8", x"a2fc7da5d62c7b18", x"92cb79f412d4ad86", x"71aae5513ff3f1d3", x"880838d78a5770de", x"8c2c43ae441424f6", x"2720438cb12fde9e");
            when 28952705 => data <= (x"be92d2c39a6f4c23", x"4d3c3fd0d5b7141f", x"94e6b36d3b547220", x"e4a6c8cfb54b96b3", x"fd4f8703a8e884c8", x"32befed9976b2ac5", x"6ec91f2085274bd1", x"8c14cdf5bc304990");
            when 4409975 => data <= (x"470c3b08e8360b35", x"b5748a7b53d36d7d", x"8715b1ed68841c02", x"7a41e6a0c563cba3", x"471e5913cc969711", x"9d5e9fb5aef5b4b1", x"e90901a07cf32c3d", x"aaf7300b5e296de9");
            when 6124916 => data <= (x"e08128d5e1f62a87", x"6267f02270e6ab56", x"5e7fe5d5d17982aa", x"b0876f5d4b258288", x"7c3d92bd17c7f852", x"990f5416e22acd15", x"868a8059fdfd7772", x"73bee95827ec560e");
            when 29058977 => data <= (x"829a8ffced49d558", x"c62bb4028066130e", x"de40c7af899fe525", x"1dd4b80fe6bfff27", x"5a4e4bd2df262df0", x"c9bd1ba20954e053", x"9fc8507f2ac32022", x"5ef86d44c10fce63");
            when 13398162 => data <= (x"b0242702ec8fa171", x"6c5c43a4024e2e4b", x"758bfa34da2d6a6f", x"9097b99471281d24", x"f36b3d7f2f7ecf70", x"319ba8ac6950f88c", x"3105318a19fe7018", x"ad7c6b2fa85d9613");
            when 1505094 => data <= (x"83fe173ec83d7dbc", x"1ba333ae9fdd1c08", x"44cfdb833620ef4a", x"ac006a232cfd3763", x"769dc8beaddc45b5", x"12173a34fbd227db", x"71046d4fb3d59f3e", x"8b08c889d4cacfeb");
            when 11775566 => data <= (x"9102bb39498a91f4", x"ff51e2045280c418", x"0c106eeef5b70796", x"9ac4dd1712596ddc", x"cde77d226e070402", x"5e151e6608ecd0b7", x"e8f009588b924173", x"348e372caeb84074");
            when 25857670 => data <= (x"45d4e9566fddc8a8", x"5e6a0e9a8b61c2fe", x"ffb995df55e50b33", x"e0c517321eaa8ca0", x"a09c8c3a7bc6d826", x"2ed37b1c3bccfdab", x"ac3a775aba484498", x"56a3b41febc56704");
            when 9573450 => data <= (x"3aee4f6b6ccf4804", x"819054aef925c5af", x"8d6560facc4078a7", x"0ec82f2a41233341", x"9185fc07ba61d556", x"786c7ffe964cb39e", x"38399b69f6766f15", x"a5bbcc6edc66855e");
            when 9782911 => data <= (x"5361d2854151b62a", x"a1ad8c39fce3d5bf", x"e70eb78cb2e79a9d", x"ead14efff9fe286c", x"5e52420c83ec0270", x"09a44343e06c51ac", x"4389c0eff110e2b4", x"b5a5e42421c1a8dc");
            when 9226238 => data <= (x"87b63f0b79368931", x"abda55aa64cbda52", x"691275515b09e01c", x"fa5a182d4ab22f8d", x"9d0528ae464f4d93", x"08266a526c88c03b", x"7a93560210624ddc", x"a2829c643b7dfb12");
            when 429456 => data <= (x"c119d5f24a420503", x"fd2f3bd13fd9d0a4", x"ecfca6a532a56ea5", x"b1903e9361c68529", x"791a22e29e9f8390", x"369a7c1b5f338d86", x"f0c03275cd3340f8", x"5f213bcc3f4b43f5");
            when 23589068 => data <= (x"e240d997380ce14b", x"b23f379914bd65d4", x"8c6a11da7f245d43", x"20bef81dc41b368d", x"e665310745f2f1dd", x"8efc73dbbefd1ca5", x"1e7d07c21701d02d", x"b026cf7ec1aeb40e");
            when 9105565 => data <= (x"ec1a4c6c191966d7", x"1a5b4023d9445ac7", x"df021198197575a8", x"4dc74e78fa561134", x"afff4748faa61d07", x"7da6605b520d3b02", x"357ca68796c2cb4c", x"741656a17735cd41");
            when 31210728 => data <= (x"c0932f7c16a2ab23", x"ad31a42cecd9872a", x"a43aa061366bbae2", x"2b23cf4a0b987015", x"5dd7490ebb4cbf88", x"b7076c30be751ffc", x"40e802ee6508d92d", x"e13b41f40b1245bb");
            when 20556537 => data <= (x"7a1156f8db766e5c", x"13bfb04049b5c556", x"8bc3bd6834c86436", x"abbd8abd8da94d13", x"7f585801e1cf139c", x"7b9985f34a2dd2fe", x"ca8d5cb7b082ea18", x"32a3eaad1212b8ee");
            when 5484478 => data <= (x"2b6ab296dc729df6", x"2deef6eee256bc71", x"8a691e29cf454e09", x"e8559cb5f346812b", x"b3e6b4fcbdaf156e", x"2736a868f71bf0b0", x"2a5332f92022e57f", x"4d956fc84c89c338");
            when 32417053 => data <= (x"4aef6ec0fd2234b8", x"a738d281502ac33a", x"d522a56cb56c5030", x"f2a105fca15b7f10", x"afaa6f734b92158b", x"469b26666e05db74", x"0610702d3d9c1a02", x"caef44cdf6d410f1");
            when 740838 => data <= (x"3fb29cb73dd6f789", x"36026c80616a5e70", x"0baf3522e31af175", x"6d53209c4f41a1fe", x"a67f15c68af544bc", x"bdf6f9c3d4455a2b", x"8723b30a42ea3aa1", x"c81216519a4d0f43");
            when 8090230 => data <= (x"0e89a6568823a674", x"a3af6332f8541e94", x"976b399315c7fcf0", x"4029f51322031ae9", x"05b7551121438c5d", x"56441f2177322774", x"b43b412c8dbc2c7e", x"c27b06c90b0d0fc7");
            when 11150229 => data <= (x"e656b38962d943c9", x"3f8a5f406b949552", x"7d6517140c33837f", x"a739d55ae113a714", x"6f17869ea1024021", x"c7976bd96c0dab5f", x"2dc06e358fdd4690", x"0b8230b249b240fe");
            when 3471719 => data <= (x"76c7774b30c9b215", x"9777f9efc47aa84d", x"9513b2e999cf9d9a", x"54f6c1ae6a3ade7a", x"63cc6e517f657fa5", x"07aa7e4b9ff7d20c", x"ccbe1bd5889f10a3", x"f55f5602f495e0e8");
            when 21501362 => data <= (x"b54092f46554325e", x"f0ff7ea2dda11d1d", x"9cf155fb1ede0c76", x"debf6540ca57dfe1", x"87e5d7bb02059220", x"bc1d45ed3812f1b3", x"b4c4a978ddfa8a64", x"d716576726daa97c");
            when 33608452 => data <= (x"9e8f82b7dbdecd4c", x"f10ca9119a393bba", x"0e687581125410e7", x"27d0e6817c55fce7", x"72d82344733746f6", x"f51c6c0c57f8d14b", x"2bf6bbfad3ddf783", x"c2951276478f3d6a");
            when 33082176 => data <= (x"042cd21c0f64b8b5", x"8135d0536d76a0b7", x"37b7ca57e1dfb941", x"9377a0f45d2a7475", x"f00650f50d5d8432", x"81e1fa563c77a194", x"ceecceaf73139d07", x"1607408b86c398ff");
            when 22732074 => data <= (x"a9aef9cca3058d01", x"9915d06d3aad3879", x"e69af7357c9160c6", x"f2e47d8bcd49b565", x"7b853666b916e163", x"ba526ff5ce2f5be0", x"7b15fb140da4ba3a", x"bc7ef310738117be");
            when 32611218 => data <= (x"1f798773942757c6", x"9d35ba3f1e915e26", x"5c59ba02ea883217", x"ff9d79d70ff22474", x"7af7ec14e9e344b3", x"361e25c94690d07e", x"8cceb4a8224927b1", x"d800ebfa482c6f64");
            when 13114921 => data <= (x"ce847d481cf30de2", x"d3bbf8d1391e9be6", x"e981244e60350974", x"bca1c88b4d24eb09", x"00210e9a9df4dcec", x"e6b5acc71ec1a144", x"74a4405b4009f78a", x"174c9a72189d9b62");
            when 18765118 => data <= (x"9986f56402f2da62", x"d5501897bcb476a7", x"90c0070fae868e09", x"21446c45f5f8c523", x"be3a2e08faede33d", x"9651c28e2b22ebb5", x"a4714a9ddd4d3890", x"f8e56b147c6de48b");
            when 16649431 => data <= (x"4434506b4f5cb97a", x"9b1ac8ae8378331f", x"70540a6a86e4c6e0", x"80cbf9b22616dea6", x"d64f8d8289812482", x"96f84df0559049b2", x"3e376d710ae2c43d", x"51d46f3a1aeeaaaf");
            when 4950710 => data <= (x"3266d0095b9300db", x"23fd5ddb754d5a18", x"8b8db4ce92a1115a", x"86f4e0b4819f0789", x"d157251b5182b887", x"d38cd3d1c74cc90d", x"40788d72d8b4674d", x"1894df4e7c42519d");
            when 7724852 => data <= (x"f7c4d159fea17dd1", x"6645daff0f24392f", x"6c1b7f5535634ec0", x"d637aa6a95b0aee5", x"90acfab51a3f624a", x"d8a61a00c6768295", x"d10d0b76bd49ab69", x"190fee26b940a038");
            when 5787543 => data <= (x"3e6f36a82c200e8c", x"da5c8f85378b9574", x"3dc0db1a32a6b072", x"dba2910479204e55", x"5f27af64a064c894", x"95cea327f27acb64", x"9bc01759270a5acb", x"fe0de4abe38b6bbe");
            when 18451598 => data <= (x"32dc10c516d44729", x"9ac143e73371f816", x"a3145139fde1875a", x"184f7598682bc8d5", x"e6b714000bb6e016", x"28c7e98a946ff444", x"d2e08a0d903c7750", x"0dbb486a6c9822f0");
            when 3086776 => data <= (x"4c27357e4111955b", x"a6091fbedada6b81", x"a77c829646518964", x"28f46dbbc6234011", x"146ba00cf46a9860", x"a5867830fafaed6d", x"fd49cbcc80967413", x"fcb50c11f0086c4a");
            when 28466467 => data <= (x"b498524c4234cca0", x"fdd51fe851773913", x"a1acb457460aff61", x"31edc3c3799f0e79", x"882ff22dcc023932", x"a692caea41403e3e", x"162db75fde81233b", x"bc14054131b6c026");
            when 25644122 => data <= (x"f6c4ec67a0dab04c", x"d3a2acee7c3408c0", x"83cfbfe2539250f2", x"e4838aa4fb2d38c3", x"3b2d9578f0dc6fda", x"77359a5ab53aba58", x"022eaadb2b79518a", x"5e5e175ee1037705");
            when 10521079 => data <= (x"ef85c119653f2aa5", x"3de5c81214f371b3", x"de631777c8484a41", x"bbfe71e090ad9de4", x"2f444af00845f786", x"dd93b214b04de097", x"556522b27baf032d", x"0d95bde8fcefc4cb");
            when 31370833 => data <= (x"d8c04bdf9f8d5831", x"d966072343432a15", x"927c8cdebb25f17d", x"c2f5aa05ac121504", x"2d33db3d9c299721", x"244d5cf97a74480a", x"6e44533d6c171557", x"06757546f659be19");
            when 9399107 => data <= (x"8f8ee9ec33a2a35b", x"bd1a0bdc73858997", x"775779e02ea4d50c", x"82d7e0cadd8c0593", x"bbc3b7c9860d01e7", x"2db2b1003ccbf195", x"6d5c3092040d4fd7", x"2c77638f10c4c56a");
            when 28065357 => data <= (x"88f7d64fb1c97ce5", x"39de1b66c8aa18ad", x"ae42693f6c3441f4", x"98c80dfbc85a9135", x"b5b95d84466439e8", x"2e1dffea52cc4127", x"82b71221b5d81f1d", x"7b38d6bb08585edd");
            when 20131248 => data <= (x"5ac29e74f43dfedc", x"ab28e685b4e3643f", x"a2cb1260c1e8bf10", x"80eb8f573894ee5d", x"9cc1b5ea3a91b11a", x"29a6585e904f39b2", x"f2960fea2b9f7888", x"2f314b38b82c7726");
            when 4284653 => data <= (x"a931414949b3a252", x"25b76a1fd5f2cfe9", x"cda1d12287ec8f27", x"c69d701adb116db8", x"ba2667398c72e004", x"1e131c2116b4d741", x"e58eaf80ad45bc20", x"6232dc485e23f56c");
            when 25220319 => data <= (x"d7d4402adb8f380a", x"f5b5afdec95b2cfa", x"8b4e8c9703211520", x"ea6240a1ad0df82f", x"b939dd9cbcbecd3a", x"829a17efdc54d12f", x"b27b41e6cca6eb13", x"12ecd3eda5ec96a5");
            when 11652835 => data <= (x"d9f97c2687224485", x"0e59af8ac588b07c", x"55d4cd004f09c90c", x"e0f766de23bbc0ab", x"4236507dc0758a0a", x"7aedacb8a32055f9", x"083534f3e5e44687", x"b0afe4dd6555ad7c");
            when 28158701 => data <= (x"4f5c4f204a4c255c", x"337dc3eee615190a", x"9ddb49626b198f15", x"1596fbee9143ad85", x"1ab239e67d894a27", x"941c733b44646182", x"1d075c385c0d2676", x"8aabf89710850e2b");
            when 2036737 => data <= (x"04281f6aa9fdb9e0", x"c7762604169b2e02", x"4b3f0806dea0b910", x"be8c2e39cd35ef4c", x"c95df374eb386c1c", x"b5be6d173b965a51", x"b27ed205e035e963", x"91cda718ac5c2d7d");
            when 15827288 => data <= (x"8e8f8abda1b980ce", x"1b8f7a05f3723a90", x"feb080f65ace5dc0", x"923f3c6665aa26ba", x"50c70e357bf9dcf2", x"f8a7adc1ac0fbd5c", x"d7098067f356c9d2", x"05f4620f54f2b41c");
            when 32610448 => data <= (x"71239c5e93976715", x"5eedbe5893140044", x"68d08d7c3828f399", x"a075bae2e360180e", x"3b811533ac811a93", x"666e81184bdaaaea", x"94f2b2e62b9cace5", x"b01d5617d6c89058");
            when 20068364 => data <= (x"529879a5dafa4aab", x"568f8a3953f418b2", x"813cf5dec7abeea8", x"fc639d9e0ae09c8e", x"21166a2294a4a193", x"d1ee942484e30604", x"ca2b3850643e401e", x"f10cb66409d4b802");
            when 13549574 => data <= (x"d6a973290e662cda", x"96b20c096371f780", x"2781352c8637c4e2", x"4d0c46151e286c41", x"ef374f555bf98aad", x"505b0b867e536297", x"af9a0fd8389af1ef", x"508c9d5b07199c36");
            when 30388713 => data <= (x"613d52a0a3ee6211", x"01a033cced031f39", x"63b81ab3876f7fe9", x"be2c108430586c05", x"8a4101574cd88bf3", x"014aa5fb205a8398", x"1d5c5fb31e9d013a", x"74a71fb4d7b0dc20");
            when 29378107 => data <= (x"04cc44ef937a41fe", x"6639e1f61b2b20bd", x"84ef0a6af8f4a18e", x"66a2cba4310beddc", x"bc7e80aec3c52146", x"2f344824bfd5ac08", x"57656bca951815da", x"46dbe91b719804fa");
            when 20181797 => data <= (x"19a546e331d0ae91", x"5ad9a7079f3d5a3e", x"1ff109af48a96b03", x"b524b65af920dae8", x"4618f0a6b682ede0", x"1668132854df85db", x"df4d60a68890d819", x"719c065aa7117c0c");
            when 23849681 => data <= (x"d96b91dd11a865da", x"cf8bec13123f4d72", x"2524b422ca498d99", x"4adad63e0b2993e0", x"1d25b48954898de5", x"5fed1e2786c3041d", x"997a6049c4b1fbf7", x"dc0dc602dd092fd7");
            when 5931569 => data <= (x"c59b7d4e66771c22", x"9390be11a3f8f381", x"4282a5e29ecada93", x"e51bbff37c5a5960", x"3de52f6ba4db1d5b", x"ce4f9c9b21196053", x"cf90ec3c6a3ce46c", x"6bd9d2e806a74a01");
            when 16322771 => data <= (x"1ccc71459c414e1c", x"3aba730310f6f68d", x"d3e828a2f28744d0", x"a2e7479a032d11e4", x"a856a1a7a7f08101", x"d9b614abd13da300", x"f83901e546cee73a", x"4ecc6028cbdaa8a9");
            when 18843087 => data <= (x"608ced778e35ef26", x"af65f46744437958", x"95a5a959fb4840f7", x"cba46fb71e8e3fc9", x"7f308344041bfd6a", x"05a34d29a74b548f", x"db899034803304d2", x"f7d345bef0781397");
            when 23648461 => data <= (x"0c718eb4168733b6", x"b31a3d7535869444", x"cdc38ddd41ad3cf0", x"068d463c742dba1f", x"4ced9f3d946f422d", x"d2e55a44fafc109c", x"f0b650cb26e917dd", x"20c141c1c0fd808f");
            when 5883254 => data <= (x"420cb8a11ddfa6c4", x"f12f2d890aae66e0", x"eb03604616717401", x"170333fc45108b56", x"58b3094c81ac5fd4", x"607b4e5d646ab077", x"204be80e815ce2b8", x"09d813d850e176fc");
            when 6778638 => data <= (x"0d86f003f313633e", x"5abdb19fa36107ea", x"19e4838fec74c3e1", x"0950bc7017344cfe", x"495c7db30a5b887a", x"d9841e624f047e49", x"26b313011614e2ea", x"6ca784de863a4be1");
            when 10594432 => data <= (x"eb364f12fbbcab06", x"a89e0aad7e2158a4", x"accbedbf6db5cd56", x"ca88b707d7b36b89", x"3a0274c4df0985a1", x"f26a66e4f74819c5", x"6c3eaf0d3f858be3", x"edfb549a0c0ca91e");
            when 22272787 => data <= (x"129b1da782caa916", x"31243e98e2c23941", x"2032db9b80b1deb6", x"c2cb4d8181c34a3e", x"20d898f045913032", x"3e4970e9a8e15879", x"7040c11d4cac7996", x"ed109d5a364f03d8");
            when 30980063 => data <= (x"d68b7e20d97f751e", x"5f8fc1dc6fb22939", x"2f6ee60f7b2ed7c3", x"dc098696fd021c16", x"76bd39623806b369", x"57c2d5f200f2c554", x"42deb84e771930e8", x"1ec0adbc599bbedd");
            when 20773515 => data <= (x"43feb27451975726", x"ce29fe32995540c2", x"05b4e7806835e29a", x"b50448310959e4f4", x"2c35b19e85d33289", x"f2544168698f2c7b", x"72b5e9f401495305", x"bbaeaa450fc957f3");
            when 30333997 => data <= (x"c664e16d6a6b4bc4", x"82ade546fe8137a9", x"5f3d2800f5ddb307", x"89ae2566a74241e8", x"5db26f6181985b0b", x"530e8d1291f3a9be", x"8d18dc934611d119", x"2fab777c2bd567e6");
            when 22521149 => data <= (x"05e57cd42c8861d9", x"5f0a4278d21e2256", x"f68419c4c736d773", x"a04896dbd33c0423", x"291eebcaed6df3ba", x"33cc3445f36368b7", x"48059a7c911186e1", x"ea7637e09d2e64f2");
            when 14175901 => data <= (x"1a9dce09b46f1119", x"12a78012af10b61a", x"ce200f0d6db55531", x"674ca07929950e59", x"8f492bb82147133d", x"a72545eafc17ccea", x"4ef53aee5a85a9b8", x"6d527a47e2813e58");
            when 18501640 => data <= (x"a531a07903f2f605", x"37633fe7ac4b86a6", x"5f96f09720032f86", x"69ef4669c239eb74", x"e43c5f4c7396f39f", x"bcb680e566c4785a", x"101ff5624958e809", x"364bed6e626604d5");
            when 5818869 => data <= (x"30ea40c12ecb6fd3", x"0ecdc637bf581762", x"e368b92b88273fd7", x"c9acf4efd5181488", x"38bc9df684814350", x"def163cabc75bace", x"47e99bf3e8678ac4", x"ee2a50a19031fc9b");
            when 8302167 => data <= (x"cc37660cd7d5f591", x"262b17fe2e16abe6", x"d3b80a273336dac9", x"98545db8fa0f7b87", x"e582591ffb64be74", x"9bd7aca4aae9b2ad", x"69e3582dffba5677", x"5188baa9f3685579");
            when 1336483 => data <= (x"09ab9c7b41f04d6b", x"410d815a0bc635ab", x"2254ae15b4d82972", x"d56603892af2dbf7", x"ca3303a47685b854", x"4a5047e6edfa1a48", x"9daf565690f93c50", x"77a7f0ea7a6a3663");
            when 25435353 => data <= (x"a845454dc440ca56", x"eb5b7434f1e8fdb4", x"b6507908f0e63d55", x"923add21cc1d4eb3", x"b0b42beb3b3f0445", x"e5d2786b9ecadd84", x"7063ebb020cb222a", x"4ff1bb3c33c39642");
            when 21393124 => data <= (x"bea3234d9cb6cad4", x"b8e4be2174a6be95", x"48556c69d6a4fddf", x"6f6dac3e73be9ef5", x"7d9543206f1ff0b9", x"c9f43508e46b404e", x"ca4860a869b21182", x"33b8854c7050fa55");
            when 11571580 => data <= (x"7067f8ae26863935", x"bfca04bc8a21a928", x"13ca78a28a9ac24d", x"8b0095ab5cd58a34", x"9403b51300fbb398", x"90da50e9b34532f7", x"f75d0089888203fd", x"39ad63192bc39872");
            when 22522967 => data <= (x"a41b7e0e033e6bb8", x"cd7e04e6681d1ead", x"20cb4de2895fa2d6", x"0136fdc6d46c8207", x"392c9386d01ac52f", x"76afebfc75b81280", x"a031cd4ce00594b1", x"c517d7ef0246c7e0");
            when 22417959 => data <= (x"1fd816178591108a", x"594b8b4412b65e57", x"492152d92f6d8593", x"f4c790bf345c6cba", x"35a2b414ea8f066a", x"4e9a615a2a7f2eac", x"1de280bbcacf9b95", x"707ee3750eb2fc52");
            when 20424282 => data <= (x"6c56c458fbb116ab", x"35fe3f6fcdd96d03", x"025ecf321a99824c", x"59228203b23777b9", x"ef70bdbdd6e8191c", x"81246e96f37f980f", x"d82d34e1c9d87e69", x"6e8fa17db3d67e36");
            when 10400610 => data <= (x"24a713f08931b948", x"36b8bf88bbc7305d", x"d7b15d3a654a8f30", x"beaccadc9cace99b", x"ba2417f6b6310bee", x"52adb71524eed1aa", x"4b6df335eee26348", x"48b7c163c40dd5d5");
            when 33051641 => data <= (x"aa9bb54d89d0f796", x"4bc205093cc694ba", x"03212dc470a93497", x"a198d9ff827c0b30", x"d9b64078834f6329", x"4c128028887ab41d", x"4ca1d317eb436d26", x"1959b7a8015d28cf");
            when 23695531 => data <= (x"476a33ffd8f2d8f3", x"74bc78245c6b8934", x"a914f8adcce2ecb5", x"97b2a633aefa8d4f", x"63dc20b9e9a78077", x"8e3e275d0b666ec6", x"b76b05961efdb374", x"a9c5f4df4a8752aa");
            when 18248999 => data <= (x"39c858ca161a6e37", x"3ce1fb0d1f61cd0e", x"8537a1ab6105bf3f", x"cac1f7dda6085484", x"6fb0b2098f5c0434", x"18d8f4ff37b0f1ba", x"0dad2a14302ef776", x"909caa59639fdbd5");
            when 23578169 => data <= (x"8ea4759b56357e07", x"4531c389c1ec94eb", x"2c4f19baf51742da", x"fd9708c27eca0e02", x"9afaf450c23c20dd", x"d49ce7cecb13739b", x"525c7bc4008060ad", x"b4a68322ab0a0bc5");
            when 21379088 => data <= (x"9c35cf99a5b03263", x"04f38fb3d728856b", x"b0c1108c805c20d6", x"f2c38d2b9e8adb19", x"7aa5a1bd3d70952d", x"e9104c02c28c33a6", x"d0b024c82d1dd00b", x"b085747769f29d48");
            when 15375257 => data <= (x"29bdf4df4043637f", x"8fb2b6c96b762882", x"e52d3c4c2fd003ab", x"bda0472d57c00e87", x"ccc9ac0b34be4c9b", x"e43dc0466be4d331", x"5b15df9938d57072", x"0c02eac9ba3ea23f");
            when 32055519 => data <= (x"f4c2a43ecd56276d", x"f4218714e4ce6a85", x"905932a5d4170c02", x"0dcc17ba60ca79fb", x"ac211f18aa363e1f", x"c6541780cc10bf6a", x"b976d22b22f4dfdc", x"83c138ce0f49458a");
            when 33753258 => data <= (x"69cab759bb6a99aa", x"b2e6b519329d84db", x"8ee03a1a5ad56dcf", x"898d092f895d7522", x"20568232ade3edd3", x"ef0586113cda5f94", x"4cd3ef0077619d81", x"647a645bb106c9b2");
            when 13988497 => data <= (x"12101fff4f3add6f", x"4fc4811c113bface", x"11c6fbe4f3b26b8d", x"80f86ff4a1c31bc7", x"7db02fbe30e3a9cf", x"7e7ac4969a5f9668", x"cd44f7ffed9405a8", x"eb88b6de04d2f66a");
            when 20325560 => data <= (x"22e585aaeac1d1b7", x"8aac9b87f0141bae", x"a805e678bf617f8a", x"fe696a9337830fdd", x"7a494dab0e28f71e", x"85afc4954be3a5f6", x"fb7ff23ba7f9e4f5", x"7fea5dd97b541d25");
            when 21094730 => data <= (x"1411277f1d5dcb77", x"13b641545a2bd837", x"d8e9e719b4f141e2", x"bb5092ecab4feacf", x"425d59d11bba39a3", x"b272258d6cbbb158", x"93de1129d4054dda", x"1937a7359731ceaa");
            when 23590231 => data <= (x"9be46e5898d1a451", x"b0c6effcbad09b8b", x"6e8a8464003a9ab1", x"1369d6ba610f4182", x"6a7c089a43f0fb33", x"97504c31426bb892", x"dc14498c562a29f7", x"5951cde7c43ae74f");
            when 976295 => data <= (x"37b03db047547ea0", x"b9b71367a7d9117b", x"feb24e2e491cef1d", x"41030ee64eae7769", x"1a7cd2c7811e57eb", x"3b2cf5e271b3e43b", x"ab0425743e85d506", x"aeb827b87b151d08");
            when 14808744 => data <= (x"71e52835625dc882", x"020f08f0910f2dd8", x"581dace4eeb1641d", x"f8ca0b1b3c5a7291", x"cb6af5e35a2d3715", x"a80bfb105e7be8a9", x"4b73b33e29ffa89b", x"5463ea3bfa051e34");
            when 21384151 => data <= (x"899003db6bc19629", x"6e12041ce98ee1db", x"1fc84329ceca62d3", x"f8b9a8d05147ae7e", x"f5670c1be434587b", x"5fb6cd50a011bc6d", x"fad6691d3a03d9f0", x"505dc75f945c09d6");
            when 20023200 => data <= (x"d8b3b151b2926601", x"c8ea784ac4769263", x"01a7e80269428e9b", x"034dcf27997cf2a7", x"4c69fce08e9f427b", x"a9d434e453b492a8", x"953971b724694c53", x"0b862a53b598ddae");
            when 886162 => data <= (x"218e4145e1e347b5", x"af0b54e385f93ee8", x"83580472edfbac9a", x"0f9e9f0f5b06c7b1", x"88d27ec856c9ffb2", x"f0e90080ecaff1ff", x"588248e36438ca92", x"9f3aae7a6eb6870f");
            when 528735 => data <= (x"43d0846219637522", x"924b437f942e660f", x"792c3f753e85f2ea", x"c0236bb0d6eb599a", x"eac83653d512c1ee", x"74eb5f8a799f06ea", x"506b50ad34e50eba", x"b8e156fa4525045d");
            when 8273754 => data <= (x"60b6a950892805bd", x"5c71125278e1a307", x"6660cf4f288b61cd", x"77f58b185b64706b", x"56274a8e8cc3ba91", x"92ce04758efd22aa", x"9b1c04acb39d4f1e", x"874be41776778d3e");
            when 1982558 => data <= (x"eaa898bf7e18b7c3", x"e46e0d0b9f5e9611", x"f9e31e8ecd094ee1", x"0227c91306798eba", x"dbdd7a33db37982e", x"2a366ba8c8dc0539", x"620e0276bea70d6d", x"4a95125878bc1b25");
            when 11682801 => data <= (x"db47c7e061d7ac3a", x"77c62c2a2d8e8aa7", x"84b7b8c45a63b64a", x"0215449525e8b081", x"a23408b77306b70f", x"b2a1c938d0fdd7bd", x"bc66ded1c7b23687", x"ad0c83c0ae980b8e");
            when 23816850 => data <= (x"43000cf190b3f10d", x"f56acd0e9e61ac41", x"836cfd1565e525f6", x"0400e0f55e388922", x"ed8ad1b00fb809a5", x"9c4f98fb8fd1698f", x"41b810a7be94c830", x"3c82214b0bbe28e7");
            when 16613993 => data <= (x"475009562fbc2829", x"7d507a5cb3f197e9", x"89aafa55e43bfab3", x"79e74924abf57a08", x"eeb5a90e36113924", x"bcfa14ed282acc4f", x"f37f52886836b799", x"7275529b3688f0d2");
            when 8084104 => data <= (x"47b4f5081be48754", x"11bb72308f1595d5", x"fff327997d63ce8e", x"5b94a3d62394161f", x"1584e62d2f022784", x"11d99f7ff07cca4d", x"635b26821c97fd6d", x"06db5ec53025a7c6");
            when 25601431 => data <= (x"63c3cf7dd10ba4fa", x"459c1d00f009c5ab", x"225a448f19e0c549", x"fc07df4854888e84", x"7f156f3ac19d4bfe", x"a5a31909dc5f051c", x"44ee464046ae2e8f", x"ee004185059e59dd");
            when 17584363 => data <= (x"4ebbd613edaa13b1", x"d829c26796f5ed5c", x"a0c63384ee03d8c1", x"db3eb957fa6c4071", x"5c3a46fdf8326b97", x"f94175bef7ebbf0b", x"9f459d3404c8790d", x"ff2257e2513a5343");
            when 25105513 => data <= (x"6804ca0f265fccd3", x"3a4d53b5ccc1f0ae", x"767f96f8d1c9af07", x"dda766aea785c7f8", x"87a43d07b6b0dddb", x"c345f022cabe5469", x"a6263dc3240147e4", x"5676ac1681ef6ce4");
            when 1472054 => data <= (x"5ea3d8a68e111b28", x"549cff9dc40936e5", x"c7be2791d3938606", x"0d76b154a06d4d8a", x"4ef010305d0b8cc7", x"e252cc33a292714e", x"7f027ce11eee58ab", x"8b17a60fdbdfb169");
            when 4953163 => data <= (x"e87e9a1633aa75e6", x"22cb39af620cfccf", x"8324a26b1f7ed858", x"5ffd027888336ae4", x"31de76faa0fb4799", x"dafcdb70c6ca5a95", x"d91298ddfe4d44a9", x"82c948a5d8eec4e5");
            when 24451056 => data <= (x"516c21f6f4896746", x"17bdbf67542d30aa", x"02f280983082e46d", x"dc2bb7c0dcf9ada0", x"45527f94b9c452f5", x"04c6a595c0cf1070", x"0f09d2dc69dc50b1", x"0f84b3bd495721b6");
            when 11922338 => data <= (x"006cfc9e9b2fc011", x"417630939bca0804", x"e11c3fe9293351ee", x"3aee6ff87579efeb", x"8a3a8759324fba21", x"0d666323c9fd7a85", x"399b8db519ec8b8f", x"1417d6b2fa2f2f2b");
            when 11403290 => data <= (x"9143066a59a3658f", x"1f617a4febdf02ee", x"b4843d82ca7eb07a", x"e02d6510c8edcb60", x"ffd057ca8aa516c6", x"9af575a1d80da251", x"dc95d02a4368e034", x"cee2cfea0b32f3b6");
            when 9660856 => data <= (x"36aec2dfa7d29049", x"9a0c5104916ff9ee", x"30865c52609f67fc", x"3b75ac8396f2a2ea", x"161f699d7c224dbc", x"87e1dd41c3b1e4e8", x"124f6ea3fc393045", x"3c3da0a50564b660");
            when 11685473 => data <= (x"725ca06569cf8a0e", x"960100cc9d910a15", x"dc1d5576e671549f", x"7cd8dc69dd38a52f", x"429964e2e9c0e59d", x"17a98428c3d442db", x"141728c87daefbd3", x"85ebd558f492d569");
            when 19086882 => data <= (x"b6efdcf207804a23", x"ef9c704ef67679e8", x"41526ab6ce257777", x"03e711decc638cfb", x"155caa7a6eec1951", x"678d33395dbd7875", x"6055fd18166ea14c", x"99247d2bbc7a8fbb");
            when 25984198 => data <= (x"19ca8a39e326d320", x"9f923116b32162d1", x"662c546bfe3fcf85", x"48a0db1ecfaefbf9", x"1b60fe22ca5ff4c8", x"be2ade2b096abc2f", x"d463c62d2acc6dd5", x"91cae28800786197");
            when 29922839 => data <= (x"8dc1b13b25a21909", x"9eef92a53301f233", x"f8d6cec6ef0393de", x"860bfc3a85cfcd73", x"c366f7c5cd486624", x"a9931cc44a33f2d6", x"03cd63deea22a9ab", x"210303923f464259");
            when 19922219 => data <= (x"06cd48adad10d2a1", x"41a27567dc8508bc", x"623af6182bf7f066", x"3335d607a3afd0c3", x"60b9c5901e447340", x"7f35f3eac60d727e", x"a16647cdcae04f0b", x"24c4ded739e6573a");
            when 30752631 => data <= (x"690f93456954a3cf", x"3c839b56f20524a8", x"ac4148aa11a11e03", x"bf8b2fb15cb95068", x"d72df9a3020a1fe6", x"2dde115e9118f25d", x"abace6a8aab02c8a", x"17c3e54fdd48a2ee");
            when 24307099 => data <= (x"3236b7cf281ffddb", x"6764e9083bf9a703", x"cbbc83c987db6133", x"9849d68f867fac7b", x"12660b65897d863c", x"dd2f22424dcc6fb5", x"a12bca2c07a63d0b", x"5f5c50d864962f2a");
            when 26113991 => data <= (x"5eaa17a87c401683", x"2f744fc75450c0f5", x"a8869670481d1033", x"bf17ecd800e1218d", x"74d9038e57ff2bc5", x"9e63a99e13600a18", x"80941b90b910e653", x"c2e989c23aaaeb21");
            when 12302394 => data <= (x"d5c2433b92599d36", x"7095f662f1819211", x"17f16211360198e3", x"52a67b58a2cc1a05", x"6a4333771d3f5589", x"b5ff89f0f1bb5a5e", x"1fd7cf2cc5a73154", x"8d901280dff51ec6");
            when 26352459 => data <= (x"1b6c576a78fb9277", x"13e6a2d14dbc98bd", x"ec6840e9c3370d93", x"96a7f02a99067253", x"6f511b41dfd90a3f", x"f2ee6b22ad4901cc", x"31a6ecef53fedd5c", x"9f0c609771040998");
            when 2731229 => data <= (x"7bb3d5e0369bdced", x"c0ec02135f3a3731", x"b1a1bfec562dc1a0", x"a52d157de4ce5f91", x"9e7085e232bb3558", x"216bc84c91992dd3", x"f56d0bfa5bcf083b", x"0f3c91940e3c8924");
            when 21235994 => data <= (x"b78055a165461959", x"a92e0c24ac54835b", x"3640f06e4a8da737", x"5a167adad437e05c", x"64f95e9e654dbc6a", x"d8c8155a65ddb5f3", x"acd12249ff88e7bf", x"7bf667d0e95ad25f");
            when 1001032 => data <= (x"c082fbc860070f2c", x"318bbfb00ca3dbd4", x"f06430e560990cc5", x"24d966022df1934b", x"8cafd49c0744ba2b", x"eb1f625bf5ccae55", x"5b20dbdc8c7deaf7", x"2bdd6cbada50c306");
            when 15251319 => data <= (x"1070591507f97004", x"a49ed6762abdf3db", x"2fe98f6296bbe906", x"061c99911e8a45ae", x"8f99e33f2f5e98e8", x"a366e394dd02230a", x"df3e05cc6e2620b6", x"153af68336afaddf");
            when 3481160 => data <= (x"a8e9f54ecabd7534", x"e31a6aae26b61517", x"af49daddebcc31bc", x"3d4a977dcb797d59", x"d8f4df5136b67c77", x"30635b66b451ada7", x"7e512d2aee740c50", x"711de86288093ad6");
            when 21457768 => data <= (x"d325e22235fde637", x"92eee0ab854cccf6", x"8ba4270ed7034915", x"281007df63fa96df", x"37ad787fef8ed66d", x"5273654630b7a668", x"0bb28abc1c360b74", x"5ae93c70067c0a04");
            when 23462223 => data <= (x"7d553527eb791616", x"4f54c3e8bb37534a", x"c204890cd82604d5", x"5de8141cd5458c69", x"31358f79b5e1a43c", x"84497da8ec785fb8", x"7b1fc1b06fd65892", x"d62240a873a0a4b5");
            when 16629845 => data <= (x"4f0f21774f0b050f", x"5bda3cae1aa59d4d", x"0b563c44e9154b1f", x"6b73dd3e00d53155", x"f02a5e8ff92826a2", x"2e3f8b2c705c3c5f", x"61b346d849e4b372", x"085dc1a741b85823");
            when 20254082 => data <= (x"5af682b944ea6afd", x"b89c632b13c812a3", x"ba4a759eaee4de51", x"b295d07a96e25a59", x"728c2ba50aaac4d8", x"f69bfe596f7bb811", x"a3e7ab46033923a4", x"1fbb3ed93089fece");
            when 2227057 => data <= (x"bb1db549ae358228", x"a48477975e99445a", x"847b046de5741e89", x"b7b50a3c7a8075b5", x"a844efb0d526db8f", x"90a0dbd845885728", x"2c67661779e9a545", x"c74e807e34478c9b");
            when 19881872 => data <= (x"73e887df42cf1ea5", x"a909a250e301c23b", x"9646b79b73662d39", x"73fa63d3d3e1c783", x"bd26148e5c9ec618", x"6807dd8c5b23beb4", x"b067e62a423148c1", x"8fb57dd208aff14e");
            when 5879060 => data <= (x"a3b3212ecb5e0355", x"3847a89ef1db742f", x"0af85927689bfb16", x"f909d5d80c55183f", x"b253b527f8cb050d", x"a59569d802dc6fbf", x"218d9be64d9ee4df", x"cf473ba32cf342b2");
            when 32847533 => data <= (x"a15525b8f4a1d741", x"816f4d936396a9c6", x"9a102b1b56334192", x"672e888a3eac8f33", x"13f026dc5270c22a", x"ccb38f85748df068", x"e3f0c0a0f46bb011", x"ba95df2264a63dfa");
            when 23821623 => data <= (x"3e44786c6d212b54", x"8698439ecd957a86", x"dd0497b0dc747fc6", x"c51e918ef5de351c", x"6a8519ca980fbc5e", x"1043fd7600c97cfb", x"db34572e8b3e7ba1", x"adc3eeb4d7f08254");
            when 8783143 => data <= (x"c28b378b34dd0e5e", x"c07143d7327515a0", x"0013595f22da3b5a", x"0ce63465472e82aa", x"4daffe1bb4a08dcd", x"28a70819f6391f0c", x"1d5e466781da5ff5", x"f00848c6e868e1be");
            when 26106636 => data <= (x"5e6e45dc3f722ea0", x"e802d795a605927c", x"32561bde3b61ac80", x"189e44c02c5a017e", x"d2256823857d7c63", x"3852b913d037c19f", x"da53243c50987d58", x"8c2ee1763f24e5b6");
            when 9716948 => data <= (x"d5f5bfe53a17ac64", x"50144b28fcf2c6a0", x"22b5998e1507a118", x"54757aec3b6d2bb0", x"bbadfaf6a0155361", x"baab04310e90c41c", x"3c157b186f5e4e0e", x"daa898e353b959ae");
            when 1816186 => data <= (x"d70241a91e138695", x"944311857622c2ff", x"5cfa509601053cbc", x"eebb3a68d558fa65", x"fffbb52f4c235d5d", x"0bd6e9a5586de228", x"60c08be78acf4c09", x"01d6cca2101b27ce");
            when 20124533 => data <= (x"d8573ddb157273d3", x"9ba97596376313ea", x"c60721c4d4f4c741", x"50c2d3e8ae0794f5", x"c8dbd7c285b8d1e2", x"ed17b95dca0c7388", x"e39b0cd16bb451e5", x"4b754a35c2f1c50b");
            when 12168488 => data <= (x"df2f5003fdc6e85e", x"7f6b4a2486f81ecf", x"e07afdd6d2ec94ca", x"5acc522b102cff82", x"71e41618294d95f2", x"b686584c2e635277", x"c5d739e87d76eb79", x"ddf972d2120df155");
            when 26677646 => data <= (x"8c1268e85d88e545", x"33fc1c121a039def", x"f7524b14a18cbf95", x"ffbcaaa9bc634199", x"56d9eb2083964c1a", x"be4a5489ce8d6edf", x"83e9d341d4f908bc", x"9e9e8d902558b5f5");
            when 12939553 => data <= (x"f0f7ad9eb091e390", x"a7a65adf8915679b", x"4bbfdb9b6e5a0c94", x"887a7e58eedf223c", x"a0d7ae9df36ecc11", x"48f5d84b57662a4c", x"80d2ad24abf38a2b", x"ca3ab64b743cec1d");
            when 10287774 => data <= (x"fc711104f0e13937", x"e02ab15bc7ecb2fb", x"390c1bda9668970e", x"c6c752812da5efe2", x"c5d13ad51dd3cfb3", x"e5565852492412fe", x"1f8d349afb8eb3a7", x"fe56e5cef06259e5");
            when 28186079 => data <= (x"2b7cb18e5c344bfa", x"a04dda41827db4e7", x"502129b3bbcfa420", x"27e89db97d236cba", x"df7dc59d9cc113be", x"61acb85af02cf422", x"9439011003fe152b", x"44f0f5039530b251");
            when 8851620 => data <= (x"088067aab8e4e9e0", x"86c7a14b83cacb32", x"54fb049b14acd8e8", x"71c3d0a33bbeaca4", x"f5dbb0898bec513b", x"c0499a486c2630cf", x"bb50408da753c0bc", x"cfb96dbefba4da09");
            when 16660346 => data <= (x"07d68e815f9847c3", x"04751036e4178b6e", x"bf20d5b90d13b80c", x"ac5271d02766913d", x"1195a6d91750eeef", x"857c790a39aa4ef9", x"6f2fcab6c18b37cd", x"637e3fe6aef23cf2");
            when 5152578 => data <= (x"7f160ed5f2259b13", x"f316e619c08ef3ad", x"50778f7474abb53c", x"b16e9fa7d8b20973", x"d4ef78bffd0795d0", x"a784c8fc02bbcff4", x"aee19563d92d823d", x"13a4b9815ba8b1da");
            when 2582314 => data <= (x"539e1feeb74cbc45", x"cff2f0a0b397cf9a", x"76aa8412f1d6a352", x"b50568ffeb830f48", x"8d7fcda3e3c39adc", x"7cf461043d5c2b6c", x"2f8f039f342bf13a", x"60efb621e5259e3f");
            when 31678687 => data <= (x"01d7b6d8cf01d8d4", x"d4520c4c6c2f4c6c", x"7fcc93d4568923f8", x"8272a360439baa89", x"70116ed1e51c3b73", x"ee1e2f467e4bb85e", x"f23ac9590c92f069", x"ae90c7b0fc96008f");
            when 33303801 => data <= (x"969ad4481ed8a8f1", x"a02dd2c2d8702676", x"0446397e1793694b", x"fb38a9d0296e512f", x"ad861470b3e2ed65", x"1b638f158e4646ad", x"10a990d22716d832", x"48fe8423b8740d8a");
            when 22198126 => data <= (x"380dd0d47ad3092e", x"00646ff3e1a8e99e", x"b6b4c2618621c3c0", x"80a332f835539181", x"77e01f251876f976", x"572c0a828f2b863a", x"7e1097dabab44aae", x"6597c161e8b8866c");
            when 28015043 => data <= (x"fb68483c5f83526d", x"31169bf0721ba6cc", x"0232f482202fd540", x"8d766009996b3479", x"0fc834dbfcff2713", x"bc8e0d7d9888add8", x"eeba45e5f95f35f2", x"c28fd04ec887187f");
            when 20941391 => data <= (x"115c940ea6f4ec83", x"a6ebce8c9864520f", x"beed7d67d639a8d6", x"1004408573cdb7a0", x"58c4cf8745b8dd7e", x"b979d7c7448b8556", x"01ad89faee9e5df6", x"c6dca044cadc5a88");
            when 18765038 => data <= (x"847487cafbd966a6", x"3c96d08f3b682e9b", x"03cddcc521da6835", x"696d8e44037bfde5", x"dfbe62516eb4e689", x"379262891fd004ce", x"a1e3510b788ca00d", x"2acee58b4366c5bd");
            when 20877486 => data <= (x"012a2da2ca301136", x"6bba72daf40aa512", x"da6fccbf257083e0", x"5a2cd65173d0f404", x"ff3d99c7d016ccf7", x"194e13d9de643ab6", x"ee664c4f6bd760d7", x"b1f8b324aac98a2c");
            when 5528907 => data <= (x"efd3934c04e5b9cd", x"e2277683978aab5d", x"b773d88dc71dd457", x"1f1c63ff25d7fd17", x"7cfc2bb1ec66b3be", x"d6ef20fc330e1ed7", x"a28b66aa8e34ba2f", x"db655868c04b4625");
            when 24721356 => data <= (x"413f4a03d046283e", x"97aea2af4d5c8b94", x"d60671ad5409d410", x"6116aed9268fc95b", x"efe0a7e5fc57b9c8", x"5ef4646f4b523723", x"493929379e0657e5", x"67f349b901f5b0ad");
            when 21723591 => data <= (x"486853e676f9c0cc", x"41c9b1df9ac708b2", x"ea9510f69c010e5f", x"dbf13198daa79bfa", x"6b77830da5264928", x"a64ab32407f961de", x"857cd9d885785add", x"66eab4a412515676");
            when 31382869 => data <= (x"f6577de0cebc0af4", x"41ebb53c130e1138", x"9f90b5771eea8b37", x"81f1e8b8b3ec80e2", x"1264353386d9c5c8", x"6911eeaf9aa808f8", x"fdab938a552b9554", x"cfffddb65ac66a1a");
            when 640887 => data <= (x"5ed348fa4def8ddb", x"996c3a828e30ae6c", x"525275cc25dc53b0", x"ba1d946e7ca6b202", x"5d4d06864a76fda0", x"1a8cd3734177da59", x"1f82cf3248ec6022", x"ecc5e61e8b94b32c");
            when 23231607 => data <= (x"944485e0a0749f78", x"a931f4551d3f2343", x"0ae0d72dd963f31d", x"2c1e5de585ce01a4", x"da957cf3b06ef80b", x"72f62fa74d6f1b48", x"7655f184e03d3046", x"cc75e3eb0d676c85");
            when 31947112 => data <= (x"2b3f91305256c2fe", x"e1a4c62af400d65e", x"2ed13c69884273ac", x"1d90b6f43e2504a2", x"c51c50c3237831a9", x"46e0fc153a14b514", x"6aef6925f34cd746", x"d2736e673277c917");
            when 23389083 => data <= (x"bebe1993d2511e6f", x"44c419ebc044b3b4", x"b13cab727f13e36a", x"34510c10008f4665", x"be6b5f54434b6d97", x"82629b836b65513a", x"1ae8ef798a832486", x"f7f063a71683b044");
            when 15066965 => data <= (x"3567a0df5cb64cbe", x"22af0da27aa1cf18", x"148323701c869169", x"920c6c33b6c8fc77", x"8ca7c789a5475135", x"bc3751d365585044", x"fcfdea40dd992ca1", x"910e43f73935d707");
            when 15492625 => data <= (x"f1604e0b56becaac", x"0c76af57c633a6b9", x"44d6a4ec30fd144c", x"0cf2e4eb067321a2", x"cfcbb9548818b57d", x"2a5ed806afd8c4b9", x"e683fd6260872db2", x"5edcb6f753f62748");
            when 22147045 => data <= (x"a399a73a96eb941c", x"415771850117eb3a", x"d9f3dce2eb1a80cd", x"787a79f9fc740e44", x"0b38ce5efed88991", x"03c4b09d515c9668", x"9b204a318fe17073", x"2003fb3fa655c04f");
            when 19600688 => data <= (x"3fb01372d3738212", x"c119861278829ea5", x"dc3e87e9548cbe72", x"7a0c98f6757d77ca", x"cda5d916bce24688", x"f828e35a55c2836a", x"79172fe5b4f39685", x"889b99fe61185d88");
            when 12264205 => data <= (x"9cd0fc7f68aa0629", x"d8b1234b7c1941c2", x"e4f32feae069d6f1", x"fc2d8627c47e9241", x"ec5e0529af25b31d", x"470e749eb1a12c63", x"949f90a6cb2c007d", x"de2e1099f98bd48d");
            when 12684577 => data <= (x"d458f33cc55c1734", x"a20122e9101d4dbf", x"09ef5399f6e3fef2", x"a1a2ec4bce33414c", x"d1434c8a9a1e130c", x"262817ec53022e0a", x"46c5963ff3f54887", x"e3e9abe52b3cd3c9");
            when 18130194 => data <= (x"0ed2fd94898964ea", x"39c55b43dfe51b4a", x"4cf8344e6da88b51", x"cfd8f0092d30e8f7", x"3ecd353f73e5b35a", x"31061294a9c51770", x"be1dbc9c11c7f56f", x"2aaa765fbc967df2");
            when 7360539 => data <= (x"34219ef5bfcbb38f", x"b13fc69e02cd1449", x"5f5685c48f8a959d", x"ba38261babee3f06", x"9e8df298f68ac9f1", x"6718456217c5ab32", x"0edfa79232d39b68", x"b1fe330bb9ce82f3");
            when 18778204 => data <= (x"f32e5beab52b0a4f", x"300c99f58fe0c751", x"5868b91ca4531762", x"0eb67a96584590f9", x"f74f6eb6e2e100f2", x"23d20b26836eaea1", x"a5fbc2f6155eea89", x"786880010fc7d777");
            when 33662092 => data <= (x"0a1f676bb2b1c9ee", x"432c4e2fb6bcb493", x"f97958936390ac7f", x"cb06b20b41ccd647", x"f9ec2bd267db8953", x"4ee97b0d0ae404f3", x"5d5da903a228e474", x"45d51238238a43d8");
            when 23393818 => data <= (x"e55af0d16134012b", x"c7a5ec397548bbdf", x"038f70c9fa0e1185", x"dd9195852a0cff79", x"561416e771cb473b", x"b53e73e367bbc0a8", x"2f88eb84af647da1", x"f39db06d0268cad5");
            when 29449860 => data <= (x"4cae3e4fd51ea793", x"859cefd81dfa1c6d", x"208688a021592174", x"9538fd9e5e52ffe5", x"ac41c602864c85d2", x"96adc2f989ab50dc", x"623519585a232f5b", x"5a1df7b765819b5b");
            when 3414856 => data <= (x"a51d32844004ee39", x"bbad5df00e259120", x"55a3ad903d4a87a4", x"911804d551f2076b", x"bbac3de3bfa13a01", x"9edfc1410fae9332", x"4a5a0fe5e5de088b", x"1db0695dfd4706cb");
            when 15080632 => data <= (x"c8cda8b608dd7c68", x"21fb7ca4f90d78bf", x"8694bfd8b5ee078a", x"9062af8d2138c4ce", x"ab515385b70e25be", x"1deaff18b8d72821", x"9fdc2866b92d29c4", x"1f49ec3fcf708845");
            when 9321286 => data <= (x"5ef911e22d59deeb", x"2be08ba5cb1986ca", x"2bf5648bbed2681e", x"92e5f642aa76fafc", x"af311540f4b57231", x"89021411203fc9d2", x"8353bb559dcdfd21", x"7742fe41ed560a32");
            when 7218137 => data <= (x"1eed9aa4fc882547", x"0b96b89673086564", x"0ecd7c9f629be815", x"aa83964b328f1e6c", x"6bb57ea4af5762d9", x"644a88fd9f33df75", x"f65c72605a811e62", x"3df5d4c8fb047bd7");
            when 16171558 => data <= (x"9473bfbe1dbdb763", x"cc6e623de4992bc8", x"10889ad852186734", x"7c48794c133c00f7", x"76d68a652d5d191f", x"24c70f1a296eedde", x"f0bce073dcb02d50", x"9f431deeb4d71432");
            when 27939275 => data <= (x"ae32cbe8c544f8b6", x"e824b4eacf9431a8", x"d55a82a23f8b4cae", x"42defd0faa2cfc5c", x"8dbc010ca62bae40", x"716bdab3b2174f1f", x"df564e1777c1f369", x"7dcef3251faca923");
            when 18979193 => data <= (x"c39bb92c41682893", x"604c6be5751ddf7b", x"45112487c4ba3f39", x"378ba4ec09c7fab2", x"bdd9a1d0a61a3a7c", x"cdf16d1f72ff7edd", x"be5d6816b35272d0", x"22de3ae7d517cc35");
            when 22942533 => data <= (x"f3f01bc042246c1e", x"1c7e220d97bcde86", x"401f69602a29d102", x"924e1aab8eb99df0", x"abcb9d86afef74eb", x"5cceed4d995eb0c2", x"89c7a8359705abd7", x"29e0d49756870e5d");
            when 9778393 => data <= (x"9fac4666b42aad99", x"52e6da25c1f5ca8f", x"cfb4c872b260a912", x"9090b574c27c781e", x"b46fe089f88f820c", x"d8b408f6c893350b", x"3f27c057b1d8313b", x"526292e0ea160d18");
            when 10455922 => data <= (x"15849b557e8260e2", x"3240a9d21b51324a", x"63aa5115541136c8", x"3a689aa4c9277252", x"9d6cba834a559538", x"d48291b4c9c889f6", x"578e8a84b0346297", x"c59626db6b907787");
            when 11273189 => data <= (x"9943257e050c14d6", x"7cb994f2a9e3bc11", x"21a50d03404146f5", x"ad6441a1752b7a95", x"071bd981d277175b", x"8807590164a0de16", x"1364d492c97dfb6d", x"10b8e3a3cd425f0f");
            when 28878114 => data <= (x"198459e0cafc7e7b", x"48e6915529ea8079", x"2bfd5c75ea2b48fc", x"d4add2e6194dbd39", x"d86a27a25cc9683d", x"03bf68f9d7d06df2", x"7e8b31ef3ffeb461", x"a3d9e76d12dc5ea3");
            when 32843002 => data <= (x"5e0e39a99b5acd19", x"d690806d4142a27b", x"b9886252fce195af", x"e745c0a6e9c80af8", x"a7d3c26561f93920", x"ccb17e12dc48a183", x"215e9f51349a97d7", x"253f77eccb2cc95e");
            when 19375546 => data <= (x"e1a234efaf3e93ba", x"2adc8fe4408e2de1", x"d20eaadcadf2f665", x"9e7a104c79182e70", x"3b4c36958ca870df", x"bdd31d0cd08e2b1e", x"6e0433d108d6ab62", x"c78e536e97d50cf5");
            when 17437491 => data <= (x"1fda091cdd5d3c54", x"e4ecc5f9f9d44572", x"5b4634f47793a5e7", x"d196d791c1813a78", x"05bd967902aaeee0", x"fa400fdde387ac30", x"37b9fcf359eaba4d", x"7f5f541f0273cf7a");
            when 32860975 => data <= (x"3691f4f43e2e31d5", x"639952adc2d88b4b", x"1f5add183af0a476", x"23107171a9e11080", x"44be4104cabef929", x"bb5562d5de9a5e4b", x"db1d68352de73728", x"1fca54a090153c50");
            when 29793016 => data <= (x"20b8b578e49a70a5", x"bbb914685fbbc989", x"a943243823071bcf", x"00fba09fb459a779", x"6eb8a4e8e2c8e284", x"62efa72d9ec81c3e", x"7cbdf3698cc48b46", x"ebaae9a66ab42516");
            when 21752755 => data <= (x"d7214dfffd2588c7", x"55e2a94a34e0d159", x"19753558783eb667", x"243cae1eb26519f3", x"dfa6579692a2a509", x"502ce62983cf3883", x"64e0b89e1d766621", x"cf6e7ec4fcda0c42");
            when 25653672 => data <= (x"fab1e2201977991a", x"1adcaa6d8a745e07", x"73c7e28ca1592c4e", x"c8ab630c3cdb5cd0", x"5de3771236723ab5", x"c56e199a1eb2892a", x"7e9005ee7511a50e", x"f8df1903e89b8f08");
            when 3303986 => data <= (x"a0d2d18eba9dcc58", x"59c2ec75463721cc", x"06352d5da7a9a353", x"7eee18b188364395", x"97f80d8fad4520f8", x"776b9dc91730dd2d", x"6108e667d402dad9", x"f99bc9c3cff04ab5");
            when 22050725 => data <= (x"f602cf2f657632f3", x"c92dc82979e2174f", x"5d033e4584b3b2fb", x"875c966b0e09c998", x"56a2b18a493fe042", x"8426c65748d486ca", x"9e451e5880d8e85f", x"70a3d51fb3d2e276");
            when 4013595 => data <= (x"95f41ac78cef14fb", x"47488382b482e952", x"f00908e1afdb2c1d", x"f308ea99bc48dec9", x"959aa4939b02650b", x"24474224530e3aa8", x"a16c86a64c92347f", x"1ef923f65f1aeab9");
            when 6691854 => data <= (x"93a0251df4cf71ac", x"d16c7395ab91416f", x"3a452bfc5035ba60", x"5d2148cb94ad3403", x"34338e89b71bdb13", x"3e7ffa018d5951a3", x"22089c7444c32d14", x"1b8bfb305ad2d757");
            when 2565911 => data <= (x"3b096eba32ff2dae", x"2a5697d450bacb06", x"5da925db31f5c041", x"b959fbb71d40d7f7", x"6c13f8336610244c", x"e73fe1691a05fc8b", x"76dc54d3ae641534", x"2a1c1acb39d6e0c0");
            when 10960865 => data <= (x"6a9c9ea3eb629d4f", x"559e52c3a2624d58", x"f99abaf65d07f2ca", x"6ad5828e380dcbc2", x"dd2830cdb69ca270", x"70657a79a7c77fd4", x"db11ad3d242f26e0", x"4aa04fd5c3421555");
            when 31499742 => data <= (x"87a336ed835df340", x"c473d804f520874e", x"0c0e5e2235a9b37c", x"03f794f2bc7b2fdc", x"d2d271948c389435", x"6472d29dc757cb10", x"aa47597b96d30538", x"48aaa1e50683512c");
            when 10201188 => data <= (x"43762c7d9383d014", x"ae7c845a6baa4ebd", x"db64e87b14295fa6", x"c2f35764371cd02c", x"b14681f2822a813c", x"234a9627d339774c", x"af8c59422d86ee0e", x"9a8d776a40a13ce3");
            when 12896552 => data <= (x"c5f365b71d980190", x"df90ede02e409d7c", x"d6be25decaa698b2", x"ca177010e913d88e", x"ce9adc5a258f2a21", x"6861069aca03b1c2", x"65d5a78933a7a847", x"fec16874e57dc37b");
            when 30217337 => data <= (x"7d4a103987963b97", x"c2e0bdbb46e3f1bb", x"3bcee3d414deeefa", x"0f9e7d6881faef28", x"7ecd650e96f8f667", x"ded215bc36e328a4", x"c7bf2e8089980b4f", x"b3bc3b4f7de476e8");
            when 16522519 => data <= (x"6f54c838b3c62c60", x"89cd4b050fb1f47f", x"2246fe0c8f3ac9ba", x"357a9a8346004f4a", x"a063385a666cb038", x"d613cde352b1a9f2", x"c86470407772bbb3", x"f2686507cce5ec60");
            when 19760678 => data <= (x"009ade1143023c49", x"c6036fb4a2620bd1", x"f64ab4d14fd8a9fe", x"f12fb9dfe102b241", x"e6c7511973dbbc6c", x"89a740e9c7e11b5e", x"b90b6638fd599c93", x"2d21d29a7bd65b97");
            when 7887304 => data <= (x"d53b2b2eb295ea3b", x"83176bfdeb7b6634", x"24c81c9c55c07a2d", x"5f83a695e713e76f", x"27be7f67e706f594", x"8c7f013703cb432c", x"f38e565032625f1d", x"a562df4f7ce0d5df");
            when 11146908 => data <= (x"a4bd3133f70077f2", x"ce5513ca0c22ad08", x"d3d5529768c2ce32", x"f9ff307b3e52dd8f", x"d8ed0a0377a1b2fe", x"a72952cab63cb18f", x"6773c9fa12a704de", x"f34921792d01a6a7");
            when 9163774 => data <= (x"872815fb824868d7", x"2a879e2dd6168c00", x"f66daddc655ba8c8", x"01294cf9b251d292", x"128451c7133b1eca", x"4d890886a3e08b3b", x"2958fd8c98abae0b", x"0dc0cf63f82dc5b0");
            when 6333695 => data <= (x"58bbda55a18d8ede", x"888370a272255793", x"d6782daa27c9a8d6", x"7e327a3ccc91c263", x"abfd1f3e335cb223", x"9535f076e704ddfd", x"30c40d5c64fecc9c", x"616f8354ffcb6f10");
            when 33393514 => data <= (x"23225427bd5d1e79", x"359b8d6be10b55dd", x"4bf3394f9e0c701f", x"68125005b3824e9f", x"7c250f326aebfccc", x"d6879cf28dcaddd3", x"ac07cf1fbaf00caf", x"0ae965c3d425b9cd");
            when 6183523 => data <= (x"2178a58b4d9dcb92", x"70e80fdc59c6b68b", x"e118866948642e89", x"4a8e95432cf748fe", x"7c70af070953f067", x"24c56c2f2863bbf9", x"03f5c69a29759e5b", x"7a6687d7f70a739f");
            when 10474950 => data <= (x"88659d2f61847306", x"2343e280e2fbabd9", x"6b99931b78843ddd", x"d9c50cccd08cfd9e", x"868b6c1d18e5e2e9", x"cc7c8c3acd099d68", x"8a4cdfa0e024224a", x"c4ae17d5bcfbd0bb");
            when 18716438 => data <= (x"cd4f37a1b60e0bc6", x"946f7bc0f0a83f47", x"249b3872cc183ea7", x"7597fe17bfac8784", x"0ec3f7bca3b24102", x"27596d720b9f951c", x"a46338da02ece577", x"7f237a9eddb66044");
            when 5330391 => data <= (x"b4c1feb197c5cb48", x"93bd673c44c3865f", x"9908d26b4da8e0d4", x"c6ebc104148ef8a1", x"aa3e4da89fc5825f", x"f83a4ce278ec93d8", x"c59ac1cd1f57b37e", x"e2d9895249744434");
            when 27102353 => data <= (x"e9fdfe792b58da96", x"93664d4be60f6e33", x"02fd1889e4e0dc3b", x"a230508cb6c5e23a", x"da89a44f929bf617", x"f9ca5dcb189613d2", x"5b9d6a13c99f2c45", x"7e8ca194f5e03d33");
            when 31725594 => data <= (x"c8e28b79b1f4ce6f", x"78a1992efd2ffbce", x"ea3684ba606e0832", x"7cd32cd6228ae493", x"a294fedd0c4eb1fb", x"aa851b81989c1350", x"0a7609cae5603e0b", x"1b9ffbbc1d2f13d0");
            when 30336732 => data <= (x"bb1b9addc36a14fd", x"5132b15925675af1", x"e7cfc325b5d3a036", x"3024ce8aef069e4b", x"2ed2344cb511d28f", x"e2808a0f15ade9d2", x"a83015eae6596c78", x"778c3298a5433717");
            when 20282588 => data <= (x"98d61d5a5fb97c34", x"123dc08bef3d63ee", x"68d7cc6074da2832", x"b542412eed235baa", x"6d6aa7cfab542495", x"27aaff8b8f2e5a6a", x"355238ddf1be0296", x"60a7b25f9b9a1094");
            when 8297857 => data <= (x"af7c2437ae17d39d", x"29971eed1b7302fb", x"ad2d7945280b2b6f", x"d5c4b348fc632942", x"ac554b23eef231f0", x"abb6138c6fec378b", x"310a8d86a88c67e5", x"c66330db02b5a26e");
            when 14827672 => data <= (x"557f1c6482147094", x"87fd27d8cc624885", x"f0923e89e9b94117", x"ef375976c6b1d60e", x"1eb950d77b929b11", x"f4b27b1d224f8559", x"c42807d5710a5ea2", x"cb0d8958ccce73c8");
            when 27234217 => data <= (x"12606751b92fe10b", x"6205095d11b4c8fa", x"fd6579e3dfa0b1f2", x"b25f2c65523eb145", x"a2619b4cf1fbcfef", x"5d6d98b6f975ce37", x"6f6eca1b767129bf", x"1ed7a0db6a14d0c9");
            when 19749639 => data <= (x"57b04b343e945096", x"ba5c3783299a75ad", x"decef8cebe403a15", x"42615dd67bf15c58", x"b2f3c2b8a83c4738", x"6a00405d179f80df", x"f9e268beb69cb0d8", x"7d7e7952db8e7ec1");
            when 26305567 => data <= (x"515c238d10d0cb5b", x"61c3b3cc04850aee", x"f1eeeb2599dc4bd1", x"6f8b8f7f05dedcac", x"be6f8372700b14b4", x"ccbe61110c57a39e", x"b81b715741584daf", x"337670c4d36d5ff0");
            when 5894862 => data <= (x"360432240e6869aa", x"4c0521fdd5c287ca", x"8c08dd252b687c9a", x"5ddf17456e9d7f18", x"9006ff6c3de2b4a0", x"1e068d7eed3e20d3", x"22969d2d32fa2202", x"758539749c59dc58");
            when 31884042 => data <= (x"4664d2a8ee04bdcd", x"d8d735dba24a7e32", x"10e9f6f0dd0b132a", x"243273ac173923fa", x"84834a29cf975cf7", x"5478ee1b6dacd41e", x"21aaf36f592e485a", x"a6efd24d5c510817");
            when 16765569 => data <= (x"6c65ae5dbad9d6d4", x"3247940160666018", x"e9464c49cfeacdeb", x"a118fa05e66d0e66", x"b6c3d9f20bd83d71", x"525bb0c8b73687de", x"291b845c7e8f4193", x"fb77700e0d9806d5");
            when 19557504 => data <= (x"9f2463f340dab8ae", x"9f5506ef2c1202cb", x"aa4ca21f372c717c", x"c0e11080eec7eb1a", x"7cd7ed7583a7864c", x"cbddf2117b553d6b", x"67f2c6e227f337c0", x"72f85cfa9f2719c6");
            when 10977465 => data <= (x"ab050ca8c3fcc246", x"083b933f783ac527", x"f6bb3e89027bb676", x"3b509ecf19212f19", x"f2975701707b9020", x"9cc01f40b628b2d9", x"bed1ddf0b024b375", x"361a546945556f2a");
            when 20262387 => data <= (x"4c49ef8957b8d357", x"a680380178d9179f", x"7d02db03f969cfd2", x"5e7433621e5dfe67", x"e758111fb6806645", x"f3adce9941ca95fb", x"23c777dc8b877327", x"5a072798870cb0ff");
            when 6250641 => data <= (x"7eebdc85830ca5e0", x"f3f0e3c95b5ae9a8", x"0a809c99926e71a3", x"e3240c030a64536e", x"a3f2ec94476b1d8c", x"c34e3d4bdb45be5b", x"dd51282e04c0cf17", x"f48f0c2512eda127");
            when 6646347 => data <= (x"e39f7dfb15414f91", x"7b89e88944dd4291", x"5db3372f9f77ceb4", x"d567178ece7b4477", x"afafa7515ee55c19", x"11dfd6ee7d78068f", x"30e07e59068e2b89", x"d965df0ab35f2466");
            when 9539016 => data <= (x"10df865dfac762f6", x"cbbc543eba301534", x"76ac6f2f8a397a27", x"9e2f96b3fc222314", x"8edd7d8fbe83e644", x"f4b6b0b7da4c8795", x"4859324b0b7380ac", x"2849065e0d6c925b");
            when 32132800 => data <= (x"6293809738e47e40", x"81c379b6943d110b", x"d5ee09d50b9640c7", x"64382216e29b7c96", x"3015ceabd9c86d69", x"d820497e5b1a87cf", x"c55814e55344669a", x"3c6e52764a0fdaa4");
            when 12683205 => data <= (x"24c01d6569770d49", x"1464e77cfcc3f19a", x"faf39d15da6548be", x"ce940d684cf53c47", x"f814678a646bdc9d", x"6e41735c432eea90", x"417db41034a8efd6", x"d036b0e09e101061");
            when 18240719 => data <= (x"b5cb0dbacb7c71fc", x"f745b182adb00dad", x"c47d4f29e8ba3790", x"35e2eeb7791253a1", x"7a2fd30ba821fc79", x"20af4e8d256666a9", x"801a813320d2fb80", x"b347661ebc8f370a");
            when 30074940 => data <= (x"38744b0b1c4a1fd5", x"3cdc5678eb91a375", x"0aeac5e97dc0aca7", x"50931af538b8508e", x"71540ac5e0d3e612", x"39797c6ce1d856ec", x"7a3ee1fd739f451b", x"8c9d2a1bb839a155");
            when 25216261 => data <= (x"1a92270bd86252e7", x"b8d582e1a2fc714e", x"899465b46a5cda44", x"a68dae8a374c2336", x"9e5232e3e85f08d5", x"c8493c39e5a8dfcf", x"7550aeb601559212", x"7a13ac2182f32674");
            when 18704146 => data <= (x"37e42065a9cf0d4b", x"0612a825b34d1a17", x"1dabdbfe52f2d95c", x"8852d088a9a12a5f", x"5da11c8096330608", x"2f34cab901973f06", x"a2abd0c6ea75d57f", x"8e08837ba6c6bdc4");
            when 19579745 => data <= (x"c2eafc13674100f3", x"600d226d4573d5fd", x"d744cee88e86a2cb", x"9a8d1b67f5138fc7", x"41dcacd1834ec5d3", x"3d84560d02e995d4", x"38cca628373f051c", x"6028bd01111fd484");
            when 18743224 => data <= (x"a86afb4004bd819b", x"46bf8222a05712f3", x"dc996b1c6557b072", x"9a3b356827e5cb02", x"87038d6a610dcf92", x"c7d442bb8b309547", x"e4f458edc140951a", x"f03fec931b1deb99");
            when 12119948 => data <= (x"ce36734cc354e35d", x"5f09c02a9db54d98", x"d24f1a60e23caf22", x"48c77525e2fcc52e", x"707539a528ed79f7", x"d8796f3e499753d4", x"f9ac6c58601b47fb", x"d603f6bfcdb2da5c");
            when 20121947 => data <= (x"2f1e0d4589039547", x"1c0788807f4b2ef0", x"18ee9718815a2925", x"0f8e60f606eca0a9", x"0819bbc36b59bc48", x"956425b62cad0d52", x"b32223fe4d85de28", x"c4f74e6a9256ffa4");
            when 29293503 => data <= (x"4cb4c6b568c0b11b", x"93e44fe960c235ef", x"f9e3e9fd5dbf3c23", x"6e9879e06f3a1da4", x"911b796965181d3d", x"7ad0cc318cd7f825", x"20be8f9d5a6d6741", x"f1a4c3967323e047");
            when 31740391 => data <= (x"4157f0fedc85eb66", x"7a5ccde65740e1b6", x"deecadd22148efdd", x"9a3e4d8fa0d0551a", x"7f9e8271547a269a", x"375b9b5eb837e5d9", x"39178ce9f520f458", x"9cd1f2458d7b50f9");
            when 21600793 => data <= (x"9afea304b9e370b5", x"52e33d767a9174e5", x"99ec30470ac04b0d", x"ebe6b963742f5689", x"b12b79db2ffab3d1", x"937ebb809df67fb0", x"bfde5c930fc574b6", x"3c838a8853ddca0d");
            when 1225163 => data <= (x"812468d56ad10f18", x"4c740b53673912ce", x"954f3a03f382a458", x"6f93e67de09c3446", x"af4174ab80a9ee5c", x"6662067c89ab313b", x"7d77273eef9a3464", x"d48c2cd9b70853ba");
            when 9648489 => data <= (x"c5cddfe9cd91a397", x"1ab8b8292a0cf59f", x"44115abbbf71b9d5", x"d78e879a109641c7", x"e8f91f9a3baff0ac", x"d653cb2cd95c597a", x"7f3d4634b984e88b", x"28dca1ee7e5e5517");
            when 26650982 => data <= (x"cc6be8831abab232", x"cb498fe487de50d8", x"ae7f31c8b8ea324b", x"9ff7f540d941d184", x"2ca965e2b2ceb67c", x"592effd11363a1bb", x"50c90c64f36f0289", x"e19b34cfcd5a3c4f");
            when 6931612 => data <= (x"c8b6c17de9e3e600", x"dc7bee2b7c46112e", x"4cc9bf89760f1aec", x"fe9b5485028028f5", x"739d1fa4079d7ed7", x"c48453298ef625fb", x"673dfab872a70a1c", x"9d9082af45bf1f62");
            when 936214 => data <= (x"8f82ba8a626e7118", x"b6d9fccd730c32e9", x"ba3a1fd38c104111", x"4844e25c6662dc2d", x"843296cf7ed49ef4", x"08db1e9fcc3b5774", x"73f95a1527e556cc", x"4b1018f101b6f8b2");
            when 20366839 => data <= (x"02676c80538152ec", x"92dcd844e6896c44", x"ba2ffbd1f2743e6b", x"be5687302eec7670", x"167b2c13acae9e03", x"a1f51072a76d3af4", x"7d964e6003183b4d", x"c20a37e84a6b8b3d");
            when 13308325 => data <= (x"e71f76ad5563635e", x"11358d942c2135b1", x"c5690cb7f76e1a9f", x"0a2436e8803f623d", x"3cd4a996430e4822", x"7a65d6bf270d0626", x"f223c8dd4b03a3b5", x"d875ad8e56e1fe42");
            when 26727870 => data <= (x"eb1732b25ba8210c", x"80daa57041d4fb84", x"c3bbf39697dc8127", x"5e2f53209ec1a701", x"4191ab9c9e25aa8f", x"ef49779f35f919f1", x"acb6151bc606e856", x"5c18bbbc3ce785d6");
            when 14139671 => data <= (x"7360c08feca7a971", x"94409959a777399b", x"3f7ea2546eabc159", x"3c971f4a9b8b15b0", x"0e45db3682b6f32e", x"fbc970b7be25fc71", x"42459581fa678989", x"bb4980e2f3d000a1");
            when 24358764 => data <= (x"1f529b40f5a01e12", x"9801d9b9280f1574", x"8cac98f3db3a85c6", x"f8ca502912bbdd59", x"cffe1f87ba08b1ab", x"66a1683f016b25e7", x"188dceedd0d7b66e", x"6f2e230c4658298b");
            when 5614577 => data <= (x"942de50d6f5623aa", x"4f5a0a462ff68908", x"d43a09f4cd2e415f", x"d47d1db4882c171a", x"44c0056f8c2d8e8f", x"7793e0baf4ea9df1", x"efcb79291b84da84", x"997f940d7f58fcfd");
            when 17977275 => data <= (x"2d9d7b41f4c119ce", x"9dd5b2e70502d28c", x"6855edee260afff2", x"02d8e8e57831ed24", x"17e0c2d4831a2793", x"06d82977d9dc6060", x"7aee923f09e37352", x"d9495d7f1481a4c5");
            when 25320998 => data <= (x"a825d18e5e6d0af2", x"6b48b2c1e3a4b251", x"ec16701f3340def6", x"c01798bc8d48dcd3", x"274c0412de718ed1", x"49fad2ecf778cc06", x"034073cfc6a2e0ef", x"2c056b52ee4c6f06");
            when 23651143 => data <= (x"7aae22e94195cdf1", x"f5f35e0bc7cc2218", x"576cc54ed7f4964d", x"4a6fe9adbcde5f87", x"1dbf60f12dd4bf9d", x"4a2e1c2d837283c0", x"744e9a4c9ecc320f", x"9a5164e793b326f9");
            when 6203318 => data <= (x"7134f3ff26660f20", x"ebcce78b75ae6db5", x"ea4d5681282b921e", x"d057fe9cb3c58bb5", x"2440d79e898a1d17", x"797d14034c4c1fc3", x"d46e96e6f6b4088f", x"7ec406515e083f9c");
            when 5615831 => data <= (x"f3535059618d6913", x"cd12332cb51d5a72", x"cdad7eb42b6eae0b", x"50b9e9968242b39b", x"a79ff5e71037d565", x"dafa3c3ae6c6d1b3", x"ba58c29616b51b8c", x"c946bcdcd3618c0c");
            when 30193386 => data <= (x"4419111355be355a", x"3adade029df8fb1b", x"b39c8019bb5ebfef", x"c149feff1515fc6b", x"a4af5ccc119e22e8", x"6565cfebd161cee7", x"85900712075df00c", x"9e4fcc9ced96d1f9");
            when 7679950 => data <= (x"70e79699b0638442", x"eea4072b80073ca5", x"9a8552aee541f66c", x"c0387fcfa2fbe7a7", x"a93945fc8dbc0df9", x"14cce5fefe45d7b8", x"ed8fbf0356ed94e6", x"77cab88b36e126e8");
            when 16343006 => data <= (x"8daa0f7d38217367", x"e54e9b983e0c571e", x"c3c5a2e240dc1638", x"b884ededf82277c8", x"7a7721f5dab18d28", x"b17e7ff597cb5974", x"8b0eba3a6fbf46e4", x"463fc4aa6d289c6b");
            when 13123229 => data <= (x"aa9ca58740e5d2b9", x"24e96435ff76a4d3", x"ae0acc54a3f2f629", x"0b920b96616ace76", x"430d99273e346b99", x"447c3f5b91152ac1", x"20acbcfa82c40c3a", x"2b5ad7a19b5af1e5");
            when 12368054 => data <= (x"f9136e0f496bb269", x"772b0ba708087ae1", x"c3711d66ab3cfff8", x"f783130aed010b76", x"46661b85b6b44d85", x"231042cc59d43f5a", x"602ba4cd3cb8eef3", x"d63d8a53f155da70");
            when 17427001 => data <= (x"82f6521aa91c1bb5", x"0db7986068040f16", x"4cdb0f29dbf39eef", x"5c81913d798c6eea", x"91d58dc896921af9", x"d8927658990b9656", x"83b2bbf516cdc525", x"a953b9ddc8185beb");
            when 17586291 => data <= (x"17784cab255cd9c7", x"e8021024c4a2d31f", x"b78575bf72a0540d", x"4550fe732f08d764", x"fc7519749396bf40", x"b76d774f2d4eeb48", x"54598400ccecd7a2", x"9971bf78ce50e315");
            when 9018584 => data <= (x"36d5cdcfaa9b2437", x"a9c28333b292f142", x"0f7b65c842f795ca", x"da62689ab561df95", x"5c01cff48e5c8d81", x"7c2bec561132e797", x"a51291e5c036b5f4", x"6b3d87df5e79aea6");
            when 16419821 => data <= (x"481abf9a6925bcd1", x"0a888d05582cbcca", x"57bbe552f6cbb737", x"05c6ef9c023cf4aa", x"76b2947688847eb8", x"557648ec25b64566", x"50cc830b552b35fc", x"a873e2b07e3b2548");
            when 21433163 => data <= (x"827d8857e8dc09a1", x"34931b56957d453a", x"734a151b1716236e", x"1c1809b88d0137ee", x"2b81a3f2e60633c2", x"18137def72cf74ec", x"ba8c34bce7258535", x"bb4d6c06f62caa4f");
            when 2201967 => data <= (x"3f798fc89fb7ab88", x"f7e17a8282ab1620", x"29fe6b5d222e18f8", x"e6ef5e37719d2d20", x"b79b74486816cd9f", x"2af5423144bf9de7", x"a67f60219b291df5", x"0156880691ab2e11");
            when 32963490 => data <= (x"325c2b7e39a8b31b", x"6aea34ed0c4e8df3", x"36b877d5c7a6125d", x"de0c3b013036590d", x"85f8213604754ccc", x"f3ae32a29b7cce9b", x"4c50f5875249810a", x"d772adc62ef118cc");
            when 26742441 => data <= (x"36d2e62be4934233", x"6ebbc7fbb636a092", x"4da6eef1de0670a5", x"44e07e106e061e9a", x"512899831b1d97bd", x"73af075ac7a5e452", x"4898bc7eb558757d", x"4134bfcd789c3694");
            when 4052545 => data <= (x"33ea73f478db2d1e", x"ef986d32abdb942e", x"2eb99df45d61d876", x"2e1af0e3ec231bfa", x"6738a3bb279eae6a", x"ee52eae406a0bd7e", x"45f038458f0001ea", x"2b15f3e3a5d41434");
            when 28342023 => data <= (x"36b724e44f77e005", x"631ee0a8c6ba6494", x"b05ffd57d5075c5c", x"e7de12ecd97921da", x"84dfb1d2959638f8", x"c6d195f69f55c72a", x"122fa28944e8a976", x"be71c5f73f222f25");
            when 678887 => data <= (x"1e75654e8d37a990", x"122ac69326381aef", x"a4a0d5e645e7b6cf", x"a7bb3bb49a104bc4", x"001e48406d40c051", x"114c1e18df1041d7", x"21ebebe7aac7f495", x"e76458940da67d97");
            when 16918698 => data <= (x"ca50377bb4e5554d", x"2b985c4699938d67", x"f401cf1356ab1f26", x"d89818607425c77e", x"236287ffc0482bb8", x"edf6b75ebdae6ef3", x"dc74eeedc8d50ae5", x"030a782cb627d251");
            when 10882921 => data <= (x"b56d83e101c2e92c", x"17ab6b296fa08f9c", x"f3fc036dde92a9e8", x"19da7f02cd03f950", x"fb1abe5b71898067", x"38fa9538cfd2ade7", x"ed3e158e0cc3f365", x"ba3178654941e931");
            when 3886922 => data <= (x"dc8e4d000fb7e014", x"fcd7c74248d186c0", x"83013705fc23a7a8", x"38d02a63b4a236b8", x"f7b3607774e27ef8", x"5236afe215b9a03e", x"c3f4f66669adcbc1", x"848204171056d60f");
            when 4257220 => data <= (x"a0d237b23b528885", x"24c4db34199feda1", x"9b5ac3a9f5e5da7d", x"8b953845b0acb380", x"9f9f986c6f792f61", x"c8a67e8a75dbd8ad", x"f4e7c63ac590bba8", x"747679a44c565fe4");
            when 929786 => data <= (x"fcca8c69850ccc9a", x"4e62c7877db0f9ce", x"671666d1c0722613", x"3489da04742a849f", x"6cb520d057db64e4", x"82403b3eab15bc6d", x"45c3089d593edddf", x"af0eeb38112617e5");
            when 31626325 => data <= (x"e8dde17b01a1d664", x"f08c508ac3f18241", x"0468e55b83b7f566", x"4810cc7b296d0282", x"ce16a1c2436ffff8", x"66477f2a980a3f9c", x"a57845d7e803b39a", x"90f873828a91f52d");
            when 11367793 => data <= (x"1dc86915eb546401", x"ab53bd48673d30c5", x"4a6cbfff94d1827c", x"913c0150c877a38d", x"a4f138d0f839922c", x"f3b1993aacbefcca", x"850945a8780f03a3", x"c820564abc30cfbb");
            when 18274000 => data <= (x"24e46c8f357dc70b", x"d248791683944b85", x"ec3b00e5cfdb299f", x"bef1ea655c6ef91c", x"b9311cced7fc2b01", x"5dba67e5acc09064", x"ae6c25f51a1734f3", x"c99f4714cfb36ae1");
            when 27132952 => data <= (x"f020feb84796aace", x"ead4b0b853759d3e", x"5dfe8aabaea9836b", x"d25d5ffc53ac7bff", x"66838341b6dd6961", x"b91ad1d4a0c50d40", x"9c996ec20c12bd78", x"864258cfa1659233");
            when 20514287 => data <= (x"400d540061ffb168", x"400769b99e58fb36", x"1f6a35596c91a00c", x"b85c637814cb0864", x"8701d020f5066e2d", x"85e22fe9a61f9b78", x"bd52a92ddf959cc8", x"7eeeef209b75bee0");
            when 20944390 => data <= (x"a02477256cb7e314", x"22e0f502ff64603c", x"c778729ff8af233b", x"e29b833e4c9831d4", x"dacb09f016ea2725", x"78a2ee48d301ba95", x"2a8a87abe415c426", x"659c32f7ad133761");
            when 12419890 => data <= (x"11bac087e770c9f4", x"9b0e00b5929c3653", x"aa3de7553d95f0a2", x"6b65468f3068c652", x"2171904541024833", x"a670d9816d8e70aa", x"a47346fa7564c384", x"6dcea444caf89140");
            when 16669454 => data <= (x"7394dac71fa2845b", x"011a7efd0af3361d", x"8ab8566584c44a0a", x"f7c443a4e9149a08", x"f258b5e4e9854873", x"f5810462bec11be6", x"81c6f8428e613a4b", x"4e3c60fcf9d41f50");
            when 9134608 => data <= (x"0f82213f24d6322b", x"bcbbc23f2385ce9a", x"b10b7444f40af42b", x"70fed08c3669679c", x"cd9e72dcb9e469f5", x"39b23bbcf1a63442", x"3a7e2afc3bc262c3", x"2dae719d3e35eb6f");
            when 13554615 => data <= (x"b8a38bd5bd4ca79c", x"80f7a25561889092", x"1e1c7b6c948dca7e", x"2959467fbd65ce34", x"40a185fccf9509db", x"36fa8c389f0d8da3", x"c1f0c91ef4987a9a", x"96e2492ff9a8fcc8");
            when 1081462 => data <= (x"7565253b6d7710fd", x"d031ae683c512f9e", x"80a1e5fe263d59c2", x"4db8ce662cb82e79", x"c0720bd7dc57ac69", x"ca12187a1a5cee07", x"b86ee2be691e1aeb", x"45899e92e485e0c6");
            when 26158877 => data <= (x"3f2ab269594b3a8d", x"8570ac22bd91722d", x"75af63dc85a3bedf", x"8833fb3001239a9e", x"f4ae61f831b6615f", x"9d946299dc7c9821", x"83f29739c6a818cd", x"ad175174ae7dd6ac");
            when 31884923 => data <= (x"f305f20f4ffb48db", x"48d9e0e0ecd27bc5", x"36b868c329c7d100", x"5577289a5b6d0591", x"a1044fe46c1dd90c", x"d9bf6f896d15d6af", x"b2082533c91db386", x"ad201c0bb75705e6");
            when 22147182 => data <= (x"f1edef1ec22829c3", x"232aa922d6d2187e", x"77b565decf435288", x"9e834403a3ab2cfe", x"bf6c2f1c07871e63", x"3c91d9a533fe0e31", x"8ed8461438f14bfe", x"5db79c2cb2d2baf5");
            when 1302847 => data <= (x"eb5e45e2ab21531e", x"f9cfe10b76d7b69c", x"9a82ffc22344cc31", x"5259af02939a5252", x"1ec34dd2a9728235", x"47b028f4e27cd5ad", x"3f995b92e5c4405e", x"5219a2a6e31ee7e6");
            when 16733681 => data <= (x"db306deb39541e73", x"da48ffdeaf5244b0", x"64040aede71d0f5d", x"da5c39b0050804fa", x"ef7d50af49cea7e3", x"7920c0774541aa19", x"0dd49bcb9df278a7", x"05e85ff8c98bcd59");
            when 6885395 => data <= (x"ce29359361e401e0", x"1cc494e5341e0563", x"94330e19cbe2366d", x"723b6ea71adbb90f", x"975ddd669c70ab93", x"9d95ad9ca5eaecbe", x"9977d01fc4f41ba2", x"c9fb1e73386d9aaa");
            when 2060808 => data <= (x"92dfc2d73dca6234", x"3a4f13831e893fdb", x"5df565e10700fa8d", x"c2fdac4273ac6868", x"8a382a4f88f5c7f0", x"7e90c9d285fe3b2e", x"5502a08c5004e3df", x"265abc089d44258c");
            when 21977267 => data <= (x"5a9120bf8c3d0f70", x"02b9fd1bce776bf5", x"07394a4d791f3683", x"a82aba4e872830ec", x"95373c4170c5db86", x"a849c81c72a926ed", x"0220788ff4f59b88", x"b74301d0565d19b5");
            when 8744166 => data <= (x"ff5c47232c8eb0a5", x"51318e69de7a2bf6", x"79ab69b0e50a9175", x"ab948389ac913930", x"98c18ec2fcdcd404", x"bd771aedca52bf8a", x"960843a2da207cfe", x"34023538f76b9130");
            when 13535500 => data <= (x"ec714a0ab4c155df", x"4d3f5a971f873ef1", x"4f97024c0530893d", x"0d922ab081afcabc", x"f0e328158d372d4e", x"0654266397f377c5", x"e740a3e53586f643", x"6ec2b65a5b5133df");
            when 8979184 => data <= (x"d7db3d1cc619a820", x"dadb314642538b09", x"5a0d5bdb4be17c72", x"962b32126dbdb5ba", x"70c47dbd1d21ba34", x"e250738b1b17de0b", x"186e004f699a530c", x"b1d3ba64ac0d837c");
            when 31648945 => data <= (x"a6d419036549019a", x"978b81896962d771", x"ae7589f94c7f43c3", x"32be445c3c8b3210", x"1de4cd929146b401", x"bdde8d6889f4b3c2", x"e831a3cec69de81f", x"1eb7bdd894550738");
            when 1483858 => data <= (x"e3488f682a15d5e2", x"e06540c5982a29bf", x"8ea2ad9eb4603617", x"5f9533cb7165d497", x"5cea9393fcbd26c2", x"fa7eca02aef25a42", x"51c1f3c7f421b478", x"97c00f4c55413638");
            when 12299901 => data <= (x"07df1480c59c4873", x"3792af7fedff5149", x"4d39c189e9c1b894", x"de4a58e2f46d331c", x"80589e5c7c316a43", x"5fd3ecd16ea24e1f", x"76b8d25bf36625e5", x"d65f5c2af5314ce1");
            when 19177625 => data <= (x"6d1cf450f7aa05da", x"2729e254dc0ff936", x"df01d664dd039fb1", x"6b419b386bfe5006", x"3535ac736bec1151", x"7057c973ff7a0052", x"e8f62ec05ce1e1b1", x"237312c526cd50bf");
            when 16285232 => data <= (x"fab00a84e3c6b71a", x"d9d6ee32ee3cc4b3", x"e97b9d3d95d6ff07", x"9d9cf88f06278332", x"88ba6b1746d6f958", x"c8e5db0b6baa73fb", x"432be2d8cbcad687", x"53f0f9c5747231c9");
            when 3372673 => data <= (x"a6a6dfcea3466248", x"a3a5ea292fdb6828", x"8406147ea8d32779", x"c25e14c087cd982a", x"d2b141432fdee17e", x"d9c80c95ac56f412", x"a15178f9be54d064", x"05e655ac37a41074");
            when 11169268 => data <= (x"b5755dfc89cf8ba1", x"f424c6b288a572b3", x"4fb264baed34dc7b", x"2ad302bcadf065c0", x"80ca7aa75bcc71ec", x"5f6b6d67ca4f9577", x"014a4b3196eced2f", x"7f05a3531304f980");
            when 31997963 => data <= (x"dfa484f222b065a0", x"841ef5753357fd00", x"6a48c656059ec17a", x"3a86522822bd4318", x"73ac80087fc4df94", x"ed3d150117181c41", x"955e80cb87d8b206", x"7388227085711d66");
            when 9530357 => data <= (x"65b6058e489e0aa4", x"0d5e326814ba1cc0", x"ecd37445b6c697cf", x"72b904b08561732c", x"ca8456de2affb15a", x"36342763ada70706", x"1397d6abe576a3c3", x"60499d4fe2c7f2f5");
            when 14965481 => data <= (x"aca85a19ebb831ae", x"3af38b3154aa6d64", x"e75e68a1f835b870", x"3249c6e757c8b4c8", x"ec66c7b7da6f64d3", x"3c1c3241be6ccaf7", x"12004ddaa68493e5", x"cd4a63ec43f3e618");
            when 26913572 => data <= (x"3a905303fe9f8738", x"a3e016cc43814472", x"aa2277d8b1b1745e", x"c5f303cfc7a65b70", x"dca62f61a9c4a610", x"dcd05f2188a3fab0", x"eb218e3544e7b105", x"e2df0e2103347d3c");
            when 10503936 => data <= (x"e9ad2a37f56ac98f", x"6c935a253c333870", x"8a98538724219958", x"9ed4cf2974f99385", x"1a2314d63cb5684e", x"5e740af9599fa607", x"7ebf5257569124cf", x"7f652ecaf777f235");
            when 11050441 => data <= (x"9680f892caf3abb3", x"37da4fbcf61cd09e", x"69ded032e80fa600", x"5602b97af3fae455", x"0b7dccea2ef0b9f1", x"b4c44b7e5e2afa97", x"1fc1f37582afa622", x"a83e3c2e2fa8176d");
            when 6994951 => data <= (x"5ec2606f446f2a69", x"ba048e45b9c56476", x"88b8ed446c42db87", x"6844b320b74590e7", x"9cb6099d6d1b3ff2", x"f380e242d4038099", x"586c05b11cb117db", x"3aac2f32425f600f");
            when 29980467 => data <= (x"b0d0efdde117da9e", x"6a1c307e8495b40e", x"6866672fd42725b0", x"e41d4db0e001de9c", x"72dc983f10827d8c", x"1c18d055c2742c2c", x"841b0268e9a40eb7", x"23db3f37662b9e0f");
            when 3516316 => data <= (x"4e6978391202df1e", x"bf66a6a1b67cccf1", x"17581e3787f54e8c", x"3fad11b03f4b7584", x"cdcdf7d60646e489", x"2d5e35f6bbf75e52", x"76bd7f67342984c0", x"0bd8027a6908df2a");
            when 31696217 => data <= (x"e87ebc978b170a86", x"1b1367dd74ce18fb", x"75e87e7aa59f1b38", x"f896d5063a755d84", x"4bb1c7765c6cc30c", x"e9efab5a44cf0217", x"f133b505bedbc12c", x"19f78e10e20ffbde");
            when 12235028 => data <= (x"6092060e49cf482d", x"3a2a876098d9a9ee", x"a1662c5e4486c4bd", x"02c9d097801a5fcd", x"b461913445057095", x"78ef3eea07a7495a", x"7a956fed126ae1a8", x"dbd33973c1d90eae");
            when 28592352 => data <= (x"8978994432fefd02", x"4730e63c5db6dc64", x"02b0ee1c13dc6fb9", x"99213fb5168c56b6", x"d023124593c3774d", x"b800e8a1bbf6739e", x"95b626b2328d2eb1", x"c40e9831beb59f63");
            when 16583161 => data <= (x"452e36700b4ae42d", x"60b9b6be8bac51bc", x"4dfa6572812eb84e", x"03d8dfa246a9cf76", x"acf4bdc3a47a82f1", x"1ce401f701ebbdf3", x"37310f465a617939", x"58d6ac95cd65f102");
            when 15893579 => data <= (x"915f7c282e27b5f5", x"67d076ab196a23a4", x"60339a279ce81f50", x"50bb029bfc9a2483", x"01710e43e11cedcf", x"d22e99a2d3a824bb", x"1e7c2b2372cfbb32", x"b3d03b9ec3be7922");
            when 1442740 => data <= (x"1a5da8653d48c884", x"21e771b4983330f5", x"46e780cbd07a15ef", x"2e49b3a845ef8024", x"6d9dbf2ea5ff844a", x"1b0c42d2b60bbdd2", x"d153507a7d303f9e", x"2dd28125bbb6bc31");
            when 5513649 => data <= (x"eb61daa700c66157", x"833894e1f2288004", x"3454954c3440094c", x"5107aa55ab5a99fa", x"2b488a997ed6f7f6", x"d171a8df790de89a", x"a9f294073dc2ed82", x"9171fabc83b04869");
            when 8447825 => data <= (x"dbd4695a1fce0cf3", x"284545d92235d96e", x"cd191b71f45a44d9", x"9d6415ff9c308566", x"4e130ff205936771", x"1daf3286700b6750", x"c807151b180903d5", x"1a151552676239ed");
            when 3595943 => data <= (x"7e1ecb3578c2132e", x"eb3a36261c86b035", x"e2742b48ddd9578c", x"1f07045bb672f0f8", x"884029f7562fe922", x"ac4f253817493321", x"ccaa2d6cb3540e46", x"d26e78a96d7e7735");
            when 27740330 => data <= (x"2010fbb55fcb1480", x"222d7ad802f7f687", x"f86f91b91472dd95", x"6728cb2f14ac9124", x"76aed328095b1922", x"94421bd741f3ed75", x"adf41a0566136278", x"54e84ed58dd3295e");
            when 10510980 => data <= (x"74202066e6baea00", x"7402710ca21b667e", x"60d926440afd6246", x"00e9b7f77bb17009", x"c26235edcef30283", x"05cf70b815d09c3d", x"ba0aa754b634eb80", x"0e634cb8e28514d1");
            when 25856088 => data <= (x"3f1001b4500daa33", x"095b244c0a2df4fe", x"5e10ddcb737189e2", x"d8bc5cf58c3f1556", x"fc65597591d03ecf", x"240fc7fdfbab678a", x"545477c79d455f3d", x"8f3e006312a8b8d8");
            when 27843542 => data <= (x"8a95927466595d0c", x"831f3bd4025860dc", x"606eaafe85139fde", x"51521861e96d1478", x"2855ad55be8dd589", x"8e38f3785ffb542f", x"f303cf69d7f5cdd5", x"b0ff3143872b5fe3");
            when 7133994 => data <= (x"f45625f3d52b92e3", x"83ab6efd1246603b", x"d7e84698066bd6de", x"a3ea01af0bfa11b6", x"28b6091f736d7d51", x"024643950badabbb", x"eb89afac95c7a884", x"d40449a3096fd147");
            when 23528370 => data <= (x"91f77aba7a32b4e9", x"9b7a5d0489a3b6d1", x"de49d0cdf229c265", x"ae8a0ffc4346ff33", x"0d651fd220f6f1f4", x"77826c9df460a3fc", x"48681d12dcedd9bf", x"a21f6c8da7aed6a9");
            when 7970044 => data <= (x"47f3cfd8a60d3303", x"b05b94b5d611d51d", x"1d88f1d5e3205433", x"d1e77d021c18b899", x"b56fb9471212ea28", x"1cb8d95e9ca0f560", x"863d7c3cacafcf89", x"c726e96cbb3f173a");
            when 20454888 => data <= (x"34ea07074c04d83d", x"ed6a2443c0611497", x"222748b6cfe5934a", x"0894f27bba303d62", x"9c81137248417e2a", x"9b1fa93f7ed6f943", x"0b441d3aacf65faf", x"b04fb4156d9691f3");
            when 29168356 => data <= (x"3a3f9148ad1319aa", x"2505da3b8769be63", x"a96794e4085571c7", x"0c1f6b46aa534197", x"d4248bea573a046b", x"d5a0210b2941e440", x"234caa5b9ebc2245", x"311bfb379d66cd95");
            when 3006240 => data <= (x"3c8bea18e95aa8be", x"76fe14a15fc63ea8", x"2cbf56680d771d05", x"6cd70312fae1d386", x"027a1401b79a5d64", x"a3cf314f588f4f96", x"9c6afda7f2a48e11", x"87a5a052d5f01fea");
            when 398330 => data <= (x"ec7af992970e79dd", x"f18e0e3f570c79c9", x"90d2bb9d4835c355", x"8ae49b5294ef8507", x"f51f77c9ff5c9e91", x"a5d80ead4aa29a9f", x"d77baf258b0812f3", x"fcd4adc205e5df7c");
            when 27487248 => data <= (x"63a7893a078d61de", x"ae6a116d5ca30597", x"56f2eae9ac017e8b", x"e7eadc5096fc266f", x"ab8ae6bfd7675196", x"289ad8ebbe675b5f", x"ddb9142b7b60cb55", x"5abe497453006bcc");
            when 1996185 => data <= (x"f05b9c1b7f2cda4b", x"7ea3e86267df9faf", x"620e8c6e36410052", x"7661e6b813386e10", x"1d4066e4b421728c", x"17fbc9acfbcdff5e", x"b9f48441bbc121ec", x"b6c72c550b59ea52");
            when 27896589 => data <= (x"df206b8a9706aaff", x"7c4693e5c89d96fe", x"4b4a7696f172f2ca", x"ad464ab5d6a4a816", x"c0567993030f2cd7", x"15c1ba6b8f864438", x"3cdd9111e918ee44", x"87194a14880f794c");
            when 14841077 => data <= (x"6c4486857321b9ac", x"2a313be2361d260f", x"63c079c95cd4f3ad", x"395d806746679100", x"6058cb886946b46a", x"cacb8c0798fa43cb", x"fa2894d9301cad2f", x"ee65cfdd38e4c84f");
            when 1289723 => data <= (x"a6a70cb9e20a9277", x"239b1cb3487c3fe1", x"b614181afbef7556", x"aed2eca15ddc0803", x"834fb198f5234041", x"d83e3f6e17200095", x"a7b22818463f1bc8", x"b0da0b11d031a9fc");
            when 17635677 => data <= (x"26a06bc904809930", x"60006123cac7dd01", x"c03ef73e12c86e33", x"8c727d4ffea5384c", x"81967a935d1c0b3d", x"922f4fba2c246e1a", x"3fc87c8b8ca0a936", x"48c04093cd7e3a62");
            when 13256835 => data <= (x"f0bcb4b68a0459d2", x"43ae1f8becd09fff", x"3127b3ec5ff19479", x"a355029b37fcad34", x"3eeaeb373216e9f4", x"ccf1971db5e86a97", x"6cfcc99b821a5780", x"4aa706d35bb5be8e");
            when 1002375 => data <= (x"dd942eb308a27926", x"41dee2fe9c515ad5", x"e69cf6922302c77a", x"cd779eefdc915a55", x"ef41df0641d4e7e0", x"37df1c7cc780d835", x"b6a5ac9afef29766", x"50ca4f0c92eab37d");
            when 33719934 => data <= (x"1870908bc65e7893", x"087ffc912ac5f875", x"7bd511c9a8d6b00d", x"c0b1f10a9f1d398c", x"04592d14c759d979", x"af0141994e3acc6f", x"cb55b6d872102796", x"1cdcbb1f71eebc9c");
            when 33422062 => data <= (x"608cb35fa09f672c", x"b3e5e2c4d7ae91ca", x"be6b1d4037e56996", x"1d6e8b5307c3a3be", x"ae663b272d0050c7", x"a1d95117d3acf647", x"6f5798eb014718d7", x"6dab59268650231f");
            when 9838518 => data <= (x"175ca4654f53b647", x"45234b784ca4eb87", x"c6daaae5724ddaa5", x"dc2bab81fba9679e", x"4d7adb36c8bc5f6d", x"1f43ab576af38d7c", x"d0050b33052a607f", x"53b767f1d027d270");
            when 23190658 => data <= (x"f9c400056b0644da", x"940d0f09a4922469", x"4d1fa08e4270cdb5", x"4b205a5258d94e66", x"266b7f1a387d0b46", x"ce0ee9b31b3714d8", x"641efa3d5a52aa2d", x"9d76bb18c207e5e7");
            when 13702054 => data <= (x"b94856f92b3a701c", x"cd6e5c99ba5cb81e", x"8543c32167e6f351", x"2ead79a00a34fdd4", x"680b6c60f89a14f6", x"9874d5f203b6e237", x"fa0fe8a60a29c05e", x"3aca4e60fb53525c");
            when 6339675 => data <= (x"ca9cd2668d155e59", x"849b0b333aaf710c", x"7ff43e4f93799e84", x"bd310fa5731b6bfd", x"9dba66dce8cae59b", x"a6e5e4c804315c85", x"a420b28c73a8d53f", x"e1c8d7bf4d37fbf8");
            when 11832350 => data <= (x"5b250ba7975b265f", x"aa9ee917fbbca376", x"b33575e15283969e", x"44e6fd0d21b8741f", x"5d0c83a9143494fd", x"2298cac67fc29272", x"8c58eefe7260f33c", x"1ba0f3483731d621");
            when 8960037 => data <= (x"2c795f96be0b8f28", x"cf1c8a7d7ef8153b", x"f3cc940dd0b558bf", x"2cc0742e329e1f19", x"520c5941d8213c94", x"67eacb2e4b803a7a", x"70360b28605e4256", x"1f1059e7859dd2b1");
            when 30013289 => data <= (x"cbc1d09fcf9db9a3", x"9b5b425584181c07", x"fbfec1d56d872a73", x"7115ec78458f4443", x"7fc65070e1c9ec78", x"74c01f06e5c78b8e", x"48ccd54858142885", x"0431c3a934b5c6c3");
            when 19411786 => data <= (x"89e9e50b2fd62187", x"212ac09e6137fd8c", x"de0e68d7fc20b8ab", x"9647feaf2d18bfad", x"e624482de5e49c68", x"fda3672654b4e0b8", x"565eb715576d0f3c", x"7f0c05a64699c816");
            when 23655759 => data <= (x"788bdc9c7ab58f9f", x"328301fc390b7170", x"111c97cbb122f238", x"26ec503cd71af5cc", x"fbf16d1ab864bfd8", x"4f4bd58d5960672c", x"db821cee7fe8459d", x"a85907c572d97d6d");
            when 9300882 => data <= (x"5fb3fb57192ddeea", x"b1d97316c5f6b628", x"f47479fd62dc5c05", x"b8572c4ed03385ed", x"2146e94f12660f25", x"7182c8abfb4cf420", x"318f8e3c46732e3a", x"4d0f91907ab4fcd3");
            when 9094926 => data <= (x"1374da0f52451f5c", x"7d09313a76e2cc06", x"b07fceb2501f7773", x"277aa5f3ea4ad9fa", x"0ec1e2dd456d1a5d", x"f3012b5b1feb64a0", x"5d422260488ea686", x"7490cce944cdb49f");
            when 24928853 => data <= (x"eec87e3475e44e5c", x"698fa7a99c48a77c", x"8447a08ea99fd7a0", x"bb5800c05668f1e3", x"2759bdc173a68326", x"b295d0efa6f9366d", x"8b9435ee5f78ca5c", x"9556a836c8475de5");
            when 29854286 => data <= (x"58df52620145c356", x"fbe19f1ea8cbc86a", x"9c3dca0a81eb4388", x"5f877be599044d3a", x"9006a89f9b86092b", x"d63bd0757d88958c", x"e6a9ff7831db1aa3", x"92c62d4b3396611e");
            when 3750795 => data <= (x"9871490c471a397e", x"4337da46c936f03b", x"558243cc4c32cbaa", x"d181dde7421acba1", x"b0111bd53febc5bb", x"1ce29c1d94a6beae", x"46448ba6dac8e8e0", x"e4a25ec1f5f5997f");
            when 24102145 => data <= (x"4646277dc6cc9d93", x"4b96925866bcda3f", x"3d7a48d6f0e2be89", x"33412278092ba874", x"3cde81c4d74daf38", x"751611e822b759c5", x"66c43c313f1fa191", x"0f229add5f12c60c");
            when 6638815 => data <= (x"0ba2ed528edddcee", x"128f3fa1aa338527", x"81e60ee3c0e382ce", x"3c5a51ef700548a9", x"d245e926b2416213", x"c581f4a180feff98", x"5d6774ae5709db0f", x"69df239e14599842");
            when 18020838 => data <= (x"c292de1b775308c9", x"d22a66d2ea1df47c", x"5f7b821698eee497", x"c87ca67a0a29fd33", x"0fd24f43d8de0d77", x"75f518c1798e4ecc", x"4415737b6f24c0b5", x"5248b9248898db66");
            when 9403512 => data <= (x"0f133a1f24fcc608", x"80e634ee02b1f259", x"96d464ffb497c74e", x"bd092adf07dba105", x"a0de674acfe6c574", x"9560f6d7846272a7", x"1b484e1e7204fe70", x"4afc969b8f804e7d");
            when 33130902 => data <= (x"b6e850e6ba2fc697", x"2f09f0dc63bd3b08", x"ecf1724f8e2b44a4", x"8bb4e1b25169cdc3", x"463405621674fa22", x"cb9098faf64d42e0", x"02ad49471b9442b5", x"4c5645e27cc6f15b");
            when 2318135 => data <= (x"0e24fb110b67bf56", x"1c1a75fc7e4f0676", x"4e05c76b84f9e6b5", x"81794b32932c6bb4", x"bea649f0c5de147f", x"c4d8c81f7f6c67d9", x"9066de18696af7df", x"9586f32cea06b9ef");
            when 12853040 => data <= (x"468b7ecefd7e30c3", x"dc01b16c69b6243e", x"3cf267c392ec0b58", x"937ac0d23e1110b9", x"7c8a2fa68916d613", x"9d42826d9a80cfeb", x"abefa98f1d76a452", x"f565e5934afd75a2");
            when 28653204 => data <= (x"a2ad949ec89e039d", x"b1d2e184520a7223", x"27694eb70b742281", x"d1873ed069c12fea", x"9a4a1473ec371adc", x"bf261d06dd3ca0c9", x"5e4df12a7fb942d5", x"226a25bc66a41706");
            when 15587799 => data <= (x"27d08d7736b55cea", x"80195d8b5afeb151", x"0c26bc0696442b65", x"9b7d4b1318b4d2c2", x"2f1156cb71ecd4e6", x"6050b0057a0b8eea", x"1b2afa68e001612a", x"74a67a55c15df779");
            when 10093920 => data <= (x"54c1726fd109971e", x"8514aeeb1f4e6ae3", x"140095736a73e65f", x"3bec339199e5a8fe", x"689e5ca7711c4976", x"016dc04251a4a25b", x"6ba37ecf3f4f357f", x"6ebd71302f750f82");
            when 1374454 => data <= (x"6cca41363d06478f", x"e87cef18815327b6", x"b3cf67a3042cf0aa", x"be7bf6c7f4c48d72", x"029063a3bed69c7b", x"b5b783e08055d130", x"faa19c81c3acbd02", x"d35765711fd287dd");
            when 28592410 => data <= (x"b60d18e6684b3fc2", x"1ae37e5f99570dc8", x"94e30625b1e5f45a", x"3e67338cec614fab", x"839e172c8b63f4a9", x"f99235397419af8e", x"626193115b5232c0", x"9c5ae05a20f3b9cb");
            when 32242213 => data <= (x"6aea0d18d4edafde", x"e81665a362faec1e", x"9c99fc9d6100e8a9", x"430fa499219c691a", x"39287f01eeebcdb9", x"5963b7848d514c61", x"57b801f59a830b57", x"9e088940d5ec19b5");
            when 19365263 => data <= (x"80e3576e732fe470", x"82db1076c31e39e8", x"83797ff7c3ba3a11", x"e06c9151e399db53", x"09a28587d20afe3c", x"085550c16374e73d", x"968e667c13ea0dfe", x"ccc84fe0bab95ef3");
            when 14322208 => data <= (x"70c32a89ecdfbb2e", x"95b9bf3e8015a3f2", x"5148e10a1e60a7e4", x"4c6c41fef7cfb44e", x"1b225e56a11f9812", x"222bd4819213007c", x"1ab67c06fbd337f2", x"e9323680f8d6e2c1");
            when 14231958 => data <= (x"a8a49ed97074b311", x"f74d2d4a263b71f8", x"0ef13d74064662d0", x"4b844074721c01dc", x"ba060b528d78a254", x"c39f9ee1e78aa864", x"8e974ef88f6443fc", x"342308055e2da499");
            when 1863763 => data <= (x"e382885976df9289", x"e174f5c489293aea", x"a372b878fbc2ba2d", x"9c1ca9c7c2d37a58", x"9c6a914c1140c2c5", x"66d0c2b3ae8ce937", x"32a7ec7d60a69091", x"be1f98059f176303");
            when 21574757 => data <= (x"4508d60a90ba485e", x"e9ff4fdd43a49d8e", x"735b75b171908e85", x"c3c595778cc53928", x"f9cf0c01a8e276bc", x"c44097a743100b8a", x"aaf5c2fd6452f410", x"8f6b329334d8bf3b");
            when 17691448 => data <= (x"da0aae6171fc3723", x"1f47d72170570732", x"6593aba80753f819", x"2392d033236eae2b", x"5c9798374a4225db", x"a7b8b0b89da9eb93", x"e4db934c9e3c744a", x"93ea848f7f98ae90");
            when 3669293 => data <= (x"fe9e39aaa596755a", x"1f3180543bb5821a", x"fef974bd1724c489", x"4229850fe49f8bf2", x"c26e5ccc2f45ebb9", x"a63f60653ec4f7e9", x"b9fe72b9900a71c9", x"b3501e3bd9637e47");
            when 5885378 => data <= (x"0dd67d7d3be76e2c", x"3cb37d6f4b49e90f", x"857eb665101e049d", x"e84d9894f30455c2", x"f9954e4e3c87da14", x"acfbba18b4ba02e5", x"2b1f1e41b08155c9", x"ec423f199f06c508");
            when 16829851 => data <= (x"e9c3ea6523746ed8", x"2c494d32b737ac37", x"17366fb0f7f315d6", x"fd79386dd464236c", x"fa2d1b22083bb08a", x"319f4c6f7edb3f63", x"1a4ea089ba6810ac", x"a3c3105ab1953b99");
            when 8840791 => data <= (x"8135d97074d6ed3a", x"d9d7eb27fc51d831", x"8350202cb1517bf1", x"ac5de7be57f84586", x"2e2c374d4a6ce04f", x"6ed5c05acf99768b", x"7313ad1705c64f4d", x"b98e25986e3fc317");
            when 23229181 => data <= (x"3ba5b81777703006", x"1f006f453cf8c131", x"69e75d576a8c574d", x"7fcbf743ce7f81ae", x"b0a8ae4aa22ac26f", x"592772cd35de699d", x"bf00cb21948a47f0", x"46de05ab0137481c");
            when 2870483 => data <= (x"5913445d5a76e62d", x"a15cade97be9adbb", x"176906f16936f05c", x"130d9e809a96974c", x"b22c95e9704207f0", x"f637a0bd2642fbd5", x"dc54fba4fa07c323", x"55a9d15afcfb2d24");
            when 22399282 => data <= (x"d67bbb793eb80297", x"2dd68436b14c8eb3", x"5d5fb9ce6e35fc65", x"6e42b624f0bca049", x"9330b288f7ca8440", x"209faf4d6b1f9d64", x"e2fb10ef242f9a83", x"3a6a0dde667966d2");
            when 384707 => data <= (x"0f1fdb4b9e798d58", x"c94bbad4241f7d9f", x"0d3c041c0322386f", x"c5a61b38dfc46fd5", x"c38d1010052a114d", x"34dbcc6c246d9614", x"5ef15bc9f40376c2", x"feeef3841f8f42ea");
            when 9668056 => data <= (x"fc9525dcbfafb490", x"3af841a482d93d57", x"522fd745b8e6843d", x"e2b9566e6e9ee16c", x"cd2d93ea1207d3d1", x"010a47975218f6fb", x"0a5330c3b6e8f490", x"852309e068e59ac1");
            when 21304125 => data <= (x"967820bcc7e1d744", x"62bae286d51905d8", x"b177ed67b7d3f84e", x"2072f07218491e51", x"cf419f8b4b9bbd9c", x"a75520f1e737e21d", x"144f6393dee70a22", x"433b4414d4cc952d");
            when 3586548 => data <= (x"945ace3224349103", x"96a0722428796529", x"493227e0a4102fcc", x"8fd9635f729f79b2", x"4e699fc9d620a510", x"f7fc44da4d303d81", x"08e692087f0ab887", x"239652662ea08289");
            when 11739364 => data <= (x"d00fbaf63b0a5cac", x"cef0e646c174d45a", x"6ef10c9e6d9d05d7", x"a191c7e51d1ebe06", x"72b59cc452bd064a", x"e7b22d1457fc24e9", x"3897c680a0cb70cd", x"091e99f40af305b6");
            when 21728152 => data <= (x"426f5300a881b193", x"5ff287febc1cc58f", x"895e32ee0bd0047d", x"05f9d75c76ba0e68", x"c2f7a2ec19048e7c", x"efc9d5c2b6618b7a", x"d56871a4e0c9b9a6", x"29c8beb285ea76e3");
            when 12164500 => data <= (x"7b518d6d77869c39", x"9769ffe25a173561", x"5c3ba27392327161", x"0c26b26e7196bee1", x"dd962f5d06fda0db", x"94e9eefe72126c30", x"5a3e0ce0a6fa93a8", x"27e8f62d51d9fd58");
            when 23372904 => data <= (x"dfd3c09ef44d6e63", x"d81fcb811c308968", x"637ec93f30c22ae5", x"a6a068185b3f47e1", x"0bc8424776a7200e", x"eb2c6e32d70bac1c", x"251ebc2deec44b3e", x"b1170c7a49e13bdf");
            when 5010409 => data <= (x"7e586f2cad961f07", x"f3b3a595ba0a6977", x"9b1b9f489010dbbc", x"a9e0bf742b379dee", x"127b7c893aefa9c2", x"8996f690e73070b9", x"076b4838bb2b52a2", x"51282b42e70bc2c0");
            when 1032929 => data <= (x"04b08da64403707b", x"0dc9d6587d8fcba6", x"0786b74f5e887198", x"b81c1d0cf0899459", x"4a5075b34984eba9", x"179139b6d6c713cb", x"64293641a92f9950", x"13bf135109f553b5");
            when 7635624 => data <= (x"33a05061a3dfe78a", x"657595dcbc9c1d6a", x"9b9964490719d729", x"7a17a299c02e23b7", x"ca143859f2d05762", x"450f205e859eeef9", x"ae7d12eadf5f1a23", x"aece1ce7c3bf3c11");
            when 10665576 => data <= (x"1f165402790da4ef", x"723131f3f7502ca0", x"b64fece59940ae90", x"b8592eae180c202c", x"487d0d0c01e7ef07", x"5315b2defc94e7ad", x"78cbb8fd032b4fe5", x"4b5960895df85d3c");
            when 14520672 => data <= (x"fdb8c5d6a46b34c5", x"a82184fa68001631", x"d9915d691138ef09", x"93b9458d0fd36e7b", x"1fab143912cceb4a", x"fb2b8fc9671596f9", x"dc6e46212f2b5640", x"4c4d41b5a52ceb75");
            when 4631205 => data <= (x"a34eef242194f63c", x"8b2d59757078bd47", x"e7abf2a417878efd", x"f97face7818b3788", x"1002537c8437f8cc", x"2b7f455c0a7d02bf", x"8282ed4adf5bed77", x"2021aca62ccc4402");
            when 1605258 => data <= (x"cffdf33c6b54b255", x"89a69a5714f1226e", x"33ac61f9ff643105", x"4ece3af975fbece5", x"2d75591e53d8174d", x"31055631dc753840", x"5eba4fa996a8308b", x"e5e426dedd902912");
            when 21400129 => data <= (x"22803092ce80180f", x"50ffb32344f98a8e", x"9be1062c7ba4a87a", x"15b8379349f2c7e0", x"d8299c5a17c32766", x"ef7034b10c43e858", x"059cd317e4170960", x"1a5c8e6cc11781fb");
            when 29120960 => data <= (x"e910e32ec8127230", x"967803bf4d525808", x"d5e900d4bbed563d", x"a3d91e63d48270e3", x"f1e91c23cd4fa6e2", x"f7b5525ff6fdfa76", x"b6110e195beda1cd", x"0be168cd5d058a25");
            when 21601701 => data <= (x"8c8a522469f1a848", x"5c878ca411f48fb3", x"8b3e5f2dbe9dc4b5", x"9dabfad4dd444032", x"27befdb6a323f6ba", x"b6aeb7582599fb52", x"5e4c52f681b633cf", x"fb2c034b3df1926d");
            when 21291019 => data <= (x"d437ebd6bdded976", x"3bd8a09ab8034e51", x"03299f1582d23c35", x"df37a0ea29badfa8", x"ae3eb358cd059979", x"d6f6e58b1eab946c", x"714eb2087ad97f9e", x"ee0d97f62c635337");
            when 4111941 => data <= (x"37c4bc0387950111", x"87fc5f7b25526fb2", x"19edb14babb4fa34", x"2cf04103e9b45993", x"ff9f9a8f0a346db6", x"e910afd9aae5f8d1", x"59d0b3e9e10e5e74", x"d817d7e9985ddd48");
            when 8948378 => data <= (x"439e2762ad2491df", x"766a1a070785ea41", x"336d7f283fed9978", x"6cef5963d23fd981", x"0c7a824358b40c91", x"6f3b95234e4441b5", x"5a9bb4e84d6f4b20", x"212c73ce9ebc1cdd");
            when 12691764 => data <= (x"3a1f7e0439be58be", x"df462805d15da9d0", x"7d53a7cebc3fba9a", x"b62831e161dab5a2", x"947812a1c86ea5a5", x"e1a16511b6b89da1", x"0cdec659eeb260f5", x"4c2c5aa1fc3519a3");
            when 30565465 => data <= (x"8c6f29ce59c7a370", x"117430b835a21117", x"40042b21c9ed6dee", x"0b8b6f887095a065", x"6bbfda24c1e393bc", x"1059491827f298c3", x"8c0748b91e698bc8", x"b3d65e1d4c3ee559");
            when 30718724 => data <= (x"511b0d28ad27b2ca", x"a9abfb6a1e942b30", x"4b7704bdbec5af5e", x"fc44de2d05b67fdd", x"cbed80d206b3c059", x"05b25f6c3e505a95", x"f85df284690ecb23", x"9e8a8ebfc3947bd7");
            when 17567738 => data <= (x"9fb51775b75907b1", x"0761629921e1bc87", x"abdfd082a3690d1e", x"1a4dc382ca4c8f5c", x"dc62fac9fc626fc7", x"c02e8248c6e7c688", x"c3c4b70c4fd8b191", x"edd7c5664d51512d");
            when 781307 => data <= (x"9b386365c315a070", x"0e64ac519f0eb658", x"64d73e5eed207710", x"3cf4170db89a2a97", x"9bb9c26135e7d61d", x"606fad89d2d507cb", x"a9dadf8b88624d14", x"77c7191b31ac8c08");
            when 1084292 => data <= (x"d008a34116196316", x"27b70729c085de6c", x"5cbe23d019e8fa83", x"85cd5d2fdf67e52d", x"1628996e1a9b2bc3", x"5663cc0d0cbaf2a9", x"9426806e9adc4441", x"43bb560966b2c1ce");
            when 8089975 => data <= (x"e7619d98b266d014", x"17fff90042fb82cd", x"06ead10bd1aacecc", x"5e6f23990a602560", x"ff893475069518eb", x"1ef68b3c5cdcd2aa", x"c3fb084d2f826ec1", x"c2e3660c1306b838");
            when 23631348 => data <= (x"a8b8e207eab0af52", x"c4a25df12e38263e", x"7af1be7f17b1b29e", x"c911719e8756917b", x"dab8f5f3b34d7f54", x"7b1714e56f5e1daf", x"d48d3f23c10fa849", x"b91724929f56e8c6");
            when 3064011 => data <= (x"84a1cd73772c620c", x"2f23c54f5510299e", x"ab57afdff8e7833e", x"fea72d0f1db4e5b0", x"4e99b7aa17f9cc57", x"7566812804f3d6bc", x"77af247f257190e1", x"e31bf6449f21dd8e");
            when 15086518 => data <= (x"a207a7c3e6f9e121", x"23c5f3d127a602f4", x"017bae8bf4977542", x"418dc3093754c36c", x"164492c95e73e81a", x"375d1a919b9849d9", x"3cb15892139059ac", x"ffa2895bb6f21214");
            when 28322745 => data <= (x"ffa75f4af17b3965", x"69f8a3b2035cf08e", x"689189f7cc4ada32", x"216d42aefc993b47", x"c0bff125dbe87b01", x"9614b78ef4d86f2d", x"62fabd584fb3a31a", x"b4b8aa5e09bbab8c");
            when 22250090 => data <= (x"b14825ac46bb65b9", x"b41467d4e15cc315", x"cb04c9ea366ae8fd", x"6efce80a61e74e67", x"ead3632d52d979fb", x"07ffb0025c658499", x"0e4118edbf9ada2d", x"ad5db04fff440e0f");
            when 33047036 => data <= (x"3171e59dfff69c16", x"10b387201538fd61", x"7f7d964e6ce44a43", x"4a439fe796018a15", x"aa7ab1b0cf4bee5f", x"a726c2a7314e7ecd", x"8b21e7963a08b752", x"3480cc4263907ae3");
            when 7399098 => data <= (x"cf97d13ead7c664f", x"d3792346ba278b9b", x"e4e3218bb67cb194", x"7f75e63d13d12039", x"ffcbff03cc543f6c", x"12e9c2b16b7a2d97", x"22d0c338f6685760", x"358ff479ce6ffee8");
            when 22289644 => data <= (x"ef5e2a59b62020c5", x"e8a2749cfbdd5de7", x"794873c1e699f045", x"f7d928f93588e3a0", x"e1555929f5637fa0", x"d8e8828121b8cb16", x"5be0561137d2a1ba", x"ed209483945e8c69");
            when 23268449 => data <= (x"a72c6443b17f9921", x"63e91dd8b42bdef7", x"866d582dcbc7323f", x"1d2198d21280f97a", x"c6e2dbad089d0589", x"2de551a09da524e4", x"da365b6d6be1fbcb", x"438a533c8c838850");
            when 24570937 => data <= (x"c46d2fb09373cf67", x"3da92f3515ae526a", x"aebf261e27cf34df", x"f7c4c94c726ac847", x"14a3859e221f2ee4", x"981c085d9830d9a5", x"b284b6632f230ac3", x"deeea704b2f3066f");
            when 26697297 => data <= (x"b700572bc2e89eca", x"942cd9a964c80475", x"8b7666f1ab556bfa", x"f9aa813e514843ac", x"563a7580be4982a2", x"8e4397f2a313c43e", x"38d65f96df53d9ab", x"1b8efe0b497ca1ee");
            when 6035895 => data <= (x"37f6291a3f82cec6", x"69d93e13e89faba9", x"2702b4a0fecbe938", x"3d3638d98f90d57f", x"d304e7ace32391a8", x"4b1975ef440f7113", x"0a4c40a0fc5a5e2b", x"6f813711753ea1a1");
            when 15371015 => data <= (x"e35cc1d30b1ab653", x"de807e3d97eb19dc", x"dc622bce28c3d30d", x"7009e22e22eeb20e", x"bcda66efc742385b", x"d28dae3bd61162f0", x"ae657627d3765baa", x"b436c20561e5a06b");
            when 26108498 => data <= (x"423fd4f538eb6d3a", x"a45228bafd969d40", x"f8a797ee490303a1", x"b85048896f7ad054", x"c9cbb526bb821d40", x"961417667a8b50c0", x"afbd68ec9f532e8b", x"497e9ec96c5f1b2f");
            when 21022339 => data <= (x"52e88fd61edbaa43", x"16341ad9b67ae1f0", x"2a660cd080a7f4e9", x"e4761272ba642bcc", x"36fc2a433d937d7d", x"ebaca41cc6ec5889", x"9154dd4cd02997ac", x"e7a9bb3ce203b35c");
            when 25011797 => data <= (x"06b161a3c5db9193", x"84b9266ce7fe8fa3", x"fa7306861530c688", x"1403a3c2926cbd3e", x"3bee9a173509c989", x"d0f4b3a300bde761", x"07a77a05abbd20d3", x"c7b149f0d0fce152");
            when 736611 => data <= (x"df2d8d9117d00bc7", x"6121addbf0dd8a30", x"92a559b72800c3c2", x"945a49cfc53f4af4", x"5a1c9914de9a5625", x"7719da8f5ae28663", x"e7da86d5c594abbd", x"b744631006c7ee0d");
            when 11787997 => data <= (x"3cac5c5f17612a3b", x"66e152f64562350f", x"20ad1a4082b53ac5", x"ee78a5ae7e02268d", x"92383dd8f761aff8", x"e228fe837fd1cfed", x"a29c4ce7f4bbadad", x"e7233c74c3d296ae");
            when 32482109 => data <= (x"e6718ffa7b4094dd", x"4fb2613ccda37d50", x"e6735b8b6e43e56f", x"3a18b7a716ea0d08", x"25c678da843b1266", x"b498d0862023a001", x"6574c93e78ec431d", x"d9469aeea15db753");
            when 5705889 => data <= (x"05c94b04c3d6b93d", x"8ea2e9676c46ed89", x"908de496357ebd96", x"b65c8be8700f67f3", x"b347ac8b6170a42b", x"d1ba77853ddc1959", x"76acfa6f4f7919b5", x"5220c2e89f994c5d");
            when 10173415 => data <= (x"aaa201c17bacba04", x"564060a54e2140bf", x"d3ee75e9a1504c84", x"eaa528c5374fe396", x"ed839f7078fd8ca5", x"0db6d029430b4923", x"8a20ad20d17403c4", x"4d1fb6988868bb8e");
            when 6106848 => data <= (x"5f2d9c2843187041", x"3a8439920d0682f6", x"fdfcc4b759a828de", x"34d20932c4fecd51", x"94fd30a329050375", x"4db01d49e50b61da", x"c785aa4d57f696e7", x"f5e5947e157e444c");
            when 12942948 => data <= (x"ed71b3c293e14f44", x"fee3fcfe8ee8699c", x"8fa11edb6abfdbfd", x"a86fb898227719ef", x"2915a662efb9a777", x"15611d4e7102451c", x"c60d6ef3669aaa82", x"a1e8320b44f734ab");
            when 7720921 => data <= (x"2caf0d4e22c0f493", x"2b7db8aa14ac3ed2", x"fd2d5f3b677678b0", x"484c4e6b4a9cea45", x"8511c484e4e00551", x"97abbf5b31404670", x"195ca0ac4fe1792f", x"7775312ba5aaeb94");
            when 8507226 => data <= (x"3f09b83ec29888cd", x"bc2402d79e61f2f9", x"df333fb68a6ab171", x"7704be58cb1074b2", x"b1c01f4c94598bf7", x"bea5477dc33ae4dc", x"e2fd96dce684eb90", x"53b6054f1cb59857");
            when 33303648 => data <= (x"754fcdfc552298fe", x"aa10a08cf17a76e4", x"d27934847c3cd972", x"fc26de624eb3dd6c", x"f1c13972abbecae9", x"f5f1ed567b4f61ac", x"9c60ccf571ccfaad", x"2574a653030d223c");
            when 12215382 => data <= (x"f197997ec39aeb2f", x"6e900a19cbd13aea", x"ea24044da1cb964a", x"a049f1fdacdb8ec7", x"78b333aad6b91545", x"431d32ab74ceeb0a", x"1f30dfa848c1db7e", x"393435dd90e19be1");
            when 726677 => data <= (x"4f18ad55f759ab2a", x"9405ba5bc79c2c3d", x"1a951f0279e26c26", x"dc6cc4215bbe0a13", x"2c372e7f56ba945e", x"6a55a7de6d13542c", x"ac2f2938e14d3091", x"f6a3438d0f139681");
            when 20729957 => data <= (x"c8311b71991b238d", x"b39fb51682e391e7", x"dc792c3b1da40442", x"b6bf540f6bb5d816", x"40462b9e7f91647a", x"4490fc358bcb94b5", x"e3fcb20412dc884c", x"1e124a0862e75f7a");
            when 27556183 => data <= (x"0b0ee1a76268a57c", x"b6cca61ba252b579", x"6fd5612bfd669f12", x"24f1c847781f87ec", x"84b94e226304c80a", x"eca2411786b7ce0d", x"118a533287cecde0", x"99cc6e34b0fefcbb");
            when 22183573 => data <= (x"4f24eeaf580d85e5", x"76d8ade10dcb4b7e", x"0592d4bd9b3653ed", x"c97aaff56c67376d", x"289814400ee15e73", x"47c69f26db3f765f", x"0c47b2d7c98ace17", x"ed12002c20665e5b");
            when 27541863 => data <= (x"40743ab9f7df3eec", x"fcd92d0b5d0b56af", x"20f992b98e46382c", x"021458c9b81ce325", x"df7d3c6e85899401", x"e6d41c6a944539f3", x"3f8dbd98d08a7095", x"9e3896bc0002e0ab");
            when 21664002 => data <= (x"1c5f87b62860e444", x"d6f5f5a34b0b82b0", x"b7963685eda689a3", x"ebab97c2ba42b089", x"b57f932cefe26706", x"1e7a50a127625385", x"6859b61007fa7522", x"c3bd9ab08e232f46");
            when 20138036 => data <= (x"d0aa0876d7e602a7", x"3d001f906e231d6f", x"daf47a1a7016e91b", x"8aae8cb21659c5e9", x"ff9aa28ce5936eef", x"949a03b636e36f59", x"32484e3fe84e987a", x"1684460d0eddc7bb");
            when 33150693 => data <= (x"1711c5e6507149c7", x"505930e3914ce988", x"ebfcf0a06b5e2e3a", x"132cd8ab4566484b", x"1860033a2e5e0a20", x"4cc265fc4f4dd4db", x"16771ef722f8e441", x"7e98c9f1d51e67c7");
            when 22352088 => data <= (x"891be1ed9eeca870", x"69dd995aa248867e", x"ae3f49e44042075d", x"748e42d4807bb0bd", x"07323bbd4f104192", x"631670350090b7c9", x"e8b87eb09cb8c983", x"0efb2b87f6b42769");
            when 25887006 => data <= (x"3e202c4d2c90505d", x"c51582c29cc3fd97", x"79ea0e1b1a383023", x"026bb5093c4fe124", x"0ff7763b5a7ea890", x"27538e83227b3312", x"48822f2cf8177a33", x"952d2df991ab8f29");
            when 6833259 => data <= (x"c99c13c6e591e39d", x"7c4be85ee31f2053", x"0dfc884b0d06c973", x"68e17b40f6acf7b5", x"db7415b43241f5f2", x"02fe57073c530cbe", x"d63998f8f817441a", x"3aa9e879bf877822");
            when 26904920 => data <= (x"90eca814807639c6", x"c5017751afcc5355", x"99239f922f0557f7", x"e446f308c6ac2f82", x"32beedfe56330999", x"234a13500008e414", x"607db918a3dace69", x"1f637ff364da05eb");
            when 25609886 => data <= (x"74fee93e8fec5c9a", x"03bf10d0abb20be3", x"660607b3385f6fca", x"b47c1f704c9b726e", x"9cf0734984004363", x"cd5cfb44f3eb8ed4", x"b842fecc3d958a17", x"e43d2c17efafa600");
            when 1987084 => data <= (x"fde2287e6b00c192", x"4bd4378903154732", x"eea82d94431ca7b1", x"08b6ab199efb92ad", x"079ea6d73673ab9d", x"fa66452b0477f570", x"8538b6a3a12d88ef", x"56d8a1855fefc8ff");
            when 24120933 => data <= (x"0707cbd9b6f99a67", x"91e6833a17570177", x"527641dbdbd86538", x"185ac4b3706bf74c", x"93a59335701f0a55", x"b27c8410d52395fd", x"55d3f38246838a7d", x"202f0c89d213c725");
            when 7055821 => data <= (x"bc29ebf62dd49274", x"16750730ad726d43", x"4d466f3f12b05bb5", x"e7dd8d6a7209bb11", x"5f6af4115b928d41", x"5fd84c72a68c39d7", x"e601f040f925aa1f", x"042e8e05fa65cbfe");
            when 20682018 => data <= (x"c7385ca36b7aa683", x"7f4d34de5e2b70a4", x"d31a733f67bf5ef3", x"c7b66a88b4bea7d1", x"3a9863af5416c971", x"cc73eb24915f118b", x"bfc7e534becab0cd", x"deb54b30be3f88c1");
            when 16956240 => data <= (x"5734c352770b681d", x"aad9094459b72e69", x"5758cffa182962b6", x"33a001cfb2a18748", x"7aa38347f21e6a63", x"bcb815a523dcc35a", x"c202180e07cb9a1d", x"e3258fce1010554f");
            when 16821019 => data <= (x"7e2655a9211ff0f3", x"bf7b5636c4310a8f", x"28bd3f9c014fde53", x"fdc5a02bc2c39a55", x"aff70313f3c26416", x"105a9d0b546ae13d", x"fab1bacfd9f8f57a", x"9259c122828a57db");
            when 27203608 => data <= (x"b048213ed83ef9cc", x"a93ee5fdd41bbfaa", x"27d6b361693348a5", x"3d657b27397fd63a", x"609c7d1a21bfb2e0", x"aea034b34dc43ece", x"826688561b5f8a3e", x"4eaa41fa04167354");
            when 7848582 => data <= (x"91ae2dcc63269572", x"595824eed5acea5d", x"9eac8cec3987442e", x"169d4ff4d8278d59", x"b0c5baed7b67b7e1", x"f1d26fbbab3cb093", x"d0179f74baf57141", x"41ee11bf3b688bdb");
            when 11434481 => data <= (x"d7c26e3b29d6ad20", x"10a6aa538ab304d1", x"fb9f62c95cc0a9d8", x"fd5d34f885bf0663", x"e571eacb8ae61c7c", x"a8e8ae5e2c6baf41", x"5d8d2d92df45920f", x"d51fd8983a2ca2dd");
            when 17720393 => data <= (x"fa0599a41a6a1821", x"26a7c9517f3973ef", x"a6269e9049cb153e", x"c62b4659c83df0c2", x"4ea315b1ebff09ce", x"89cd87220d04cbbf", x"040461f7a406b21a", x"669e8c27f8602e18");
            when 33414329 => data <= (x"e25dd0d002292022", x"cd28c4b5da6c289c", x"fcd6c3472f18f65e", x"ad9ae9ec01e7b959", x"c23c18a00820c243", x"5476f6a09c25f474", x"69a3f42881665278", x"00a63c4aa4e3da28");
            when 3258333 => data <= (x"9b1a49a5556e33b9", x"79e737322c132d2d", x"f291736cc3687e82", x"1e19ce54bf985c0d", x"2cbe246cb69e615e", x"371f65e0808da128", x"1d91e6418ea2c100", x"24af1503dd9b0135");
            when 7322917 => data <= (x"940036f3dfd7849f", x"f6ed35d842617d1d", x"faac42bb98bfeb49", x"774570ee56a64836", x"1296f3bfca2aaa9f", x"bdc9b03738035d03", x"24e5268bbf2dcafd", x"fa1165f44f661296");
            when 26157164 => data <= (x"54ab54e8bf3cb813", x"84ba2995a7e60f0e", x"a143344f42029822", x"9aafe720329c202d", x"2c2742b7c9d36275", x"eacdab6864ad8d2c", x"827435a717c7b680", x"9daa63d0a95461fa");
            when 716143 => data <= (x"372a563c517ce5c2", x"403e84f46d816cc1", x"09221534187180a3", x"dd0de4715ecab591", x"e1f5dd808d408b72", x"f13a89060b8325df", x"33bd0b29a5f0580a", x"2eab54347dc57e6d");
            when 550116 => data <= (x"1b03c207459c84ca", x"6933a42f4e1bed55", x"98b116b5c0c32b07", x"867f6db949315959", x"52e7f5a1de469147", x"a560a0f3e3e3eb3f", x"7724b3309ac945f4", x"795e64130346ce80");
            when 21336771 => data <= (x"0aa47a5241e59d62", x"d38b4e4537ada2c2", x"76c7b2da21f120ff", x"25c1ec73b49d5d5d", x"10f5f074920d67ef", x"ace07eae7a43f9ca", x"c0ce0a6d2e6430cf", x"1a31dc1d0f30fb90");
            when 20484047 => data <= (x"0f0c7da30d1d5af6", x"13df50ac040d63a2", x"a18bb12e0af773b2", x"8178a8d80981f1a0", x"a3b22b6e0ba1102f", x"2ecb26c7a2bcdbb7", x"74e18328a91779a8", x"78cc3bd0f177b369");
            when 9015078 => data <= (x"b96617f5dd96704f", x"b4cf677338445d4b", x"aedb81d318468afa", x"042d70a1f5ff7c48", x"b0970b0d9785663c", x"8320bbf5cf3ced32", x"a6390296aa58bedd", x"a01edeeef31bda83");
            when 10551531 => data <= (x"635488b3f326f368", x"cddba7429041603f", x"e7997f8e96bbf0e2", x"c784019483adcd8d", x"f466c4f2c501636f", x"af6012ea6664c318", x"ff4668c93431f178", x"7f48c9baefbc6065");
            when 23307554 => data <= (x"94fbd8acd803e872", x"532de71afd7de786", x"f0b2a45c3876189d", x"e8ea4e6703af8188", x"b4386103ca170523", x"3aca68247e6f10c3", x"f8f92ec823dbdf75", x"e663bc48e4b9a6ca");
            when 12226858 => data <= (x"3c1c4aa4f8e4dc64", x"e900661be36db2b7", x"01cfccfccef2efd8", x"315b575466af7e52", x"51fc240fcd687673", x"964d692d62df5ae7", x"de4234495c00cc59", x"b8a2e6389a19352d");
            when 27411155 => data <= (x"70b6b779138291f4", x"7dde3f303e7c7648", x"1abb4a6996944287", x"8bf680a9ca984907", x"cc335065c314972c", x"590f04844ee0ea7a", x"aff749f7314bd58b", x"f8d2ad60dd05cdeb");
            when 28787905 => data <= (x"3486611ff7e097b3", x"7ebe0fa06b3e503d", x"eab51aa0fc4c126a", x"24a890ecbf84f634", x"d6b8b9e8fa98cbff", x"2aafcb3e8d12495f", x"902facee7f7ad96f", x"8d027d877c7fb9bf");
            when 30162553 => data <= (x"628a35b99d1e2105", x"ea9e343714b111ac", x"73260070a6eea9ce", x"e0dc42b026256ac6", x"0c4a9690583b7706", x"d20f8b290e25fe19", x"af02e37a3accfc6f", x"63efcfc8c6c4379f");
            when 13445267 => data <= (x"647463df0f8d574d", x"7409b54b8050603a", x"89f15fd7f2e329db", x"acf517d9d997f5b7", x"184ff98ee6caa3d3", x"3a985a210e4a38f8", x"4da750c11a197ac7", x"1db9b7d0c6d4636f");
            when 19020615 => data <= (x"335e5cc504e52345", x"e6aba8873e4827b5", x"bf6b766f8c96e067", x"7e3497655ea60e37", x"39f5c277e70c67f4", x"5546340cc261fb34", x"3da95885cef93e27", x"852ffc1fa90eed4a");
            when 24056569 => data <= (x"08639048f3423ce0", x"665e76b2358b7bb9", x"ab58e6ff1f9a1b66", x"fa3f294ca6d2e487", x"8c096988022ada0f", x"88cb899f0324bf26", x"11cfe5fc30c3b4d8", x"1d042ba4279b5fa0");
            when 5032103 => data <= (x"3fe8479f6452806f", x"c80212392ff68c67", x"61b6e4e9776bb851", x"0d6ae32681cc9d52", x"b0ab6c7b05041038", x"9fc7ec41dfac9ea2", x"4d4596dafb7053cf", x"a14a66d8a4a0497d");
            when 19279396 => data <= (x"be018055baf502be", x"17db210eff11390e", x"f799755fd8fe96be", x"70ec8fcefc902ee7", x"3927d83899d10a6f", x"7f4639ba255e0ff5", x"77becb8561acbc70", x"6289c9af9facd3ca");
            when 806500 => data <= (x"c87139c8f8fa42f2", x"d1d5ba7a656caee9", x"f32cceb4c4c93e3b", x"ac24edda4e8dd8ef", x"ff39b4073194c8bb", x"ba6a262a5987d0d8", x"2c414563ed96c9bb", x"fbda46a84571b9db");
            when 21879118 => data <= (x"db5487c74119419c", x"856d3856cbb45707", x"2aab3769613913ba", x"d023552ff5af4bc7", x"0b3dec1873733139", x"ead3b6ed7f607e32", x"d3eb5f43497eeffa", x"0a42210b94ad87cb");
            when 23878164 => data <= (x"5c9dc6a9c03b6a4c", x"80be2293eb5226d1", x"85b2c252e647d274", x"6cf240a67088ebb6", x"782dfad0aefb9853", x"d35108d12bee4d99", x"89d7e2acedafc4fa", x"94c34f3e62f1e3d8");
            when 11209989 => data <= (x"2380be219a069f1d", x"3b9ac968c0751ec4", x"d89b0aad00f02bba", x"554dcd42976bf2b0", x"7d6e27c91eb40b5a", x"8c651bf65b6b61b2", x"7d0f3dd2c8cdda34", x"c2b740adef3fd39d");
            when 32131351 => data <= (x"5bcb8b4d57269b35", x"f8272efc3671c02c", x"67c6db04c6090a65", x"0c9be0fa001b1abb", x"c9dc03cf4f012442", x"93d9d5d28a0b4823", x"301e504f093e361a", x"e33bc3bdea921ec2");
            when 10142814 => data <= (x"8f1bbdc34de0e9a8", x"d14b34dd17dd1928", x"3bb137579c609665", x"5eb10e5aa523ddc5", x"98b7e8f6c7a10d27", x"414386c71c6c0bd2", x"8910603b32886509", x"5f30cedf360a2bc8");
            when 22858022 => data <= (x"45d1ee92489daa68", x"be850728a8923d6c", x"5d20863a7d1bb0b0", x"e94fe4e088562953", x"28cc2bed994300a0", x"0bbd7df968c140a5", x"7e6b3f903d207df4", x"d1b4c032801fa8c0");
            when 16578749 => data <= (x"cda0dd4b3da8dc24", x"4ab645178344f0ba", x"38698564e77724f0", x"cea7d0fbf7503ab7", x"4f523f4bd0a440cc", x"b35a32484231095a", x"c8508886d61d9786", x"cf13061b609e7066");
            when 7894451 => data <= (x"1940b1e5accc816e", x"df70264a9f60ba5e", x"434d6de3184b6d8e", x"7845353335c2e221", x"1a2d655bd88c75ad", x"c5f5140b22ba1726", x"74acacc532c9f200", x"c01a8d6a3206b2ea");
            when 23614815 => data <= (x"53662c707a6c72a0", x"dcf2928099ce365c", x"d817c14ba81f866b", x"1afe9baeae9546dd", x"d385f31a8e2739c7", x"60451ec7d194826c", x"e9714d93ec3da531", x"bd4079788f3e8a52");
            when 24135407 => data <= (x"c106cc890418d782", x"1f5959360fba089c", x"881fe8b403549890", x"d4c509bc13da620b", x"7b7019f2b646e36a", x"9a26566627eb0ee9", x"98cb043bf3946d5e", x"00742bc0078cf8ea");
            when 5622372 => data <= (x"82cb3cb510daf3a5", x"41b18b00c90e3b4f", x"994dbd6e3adf86ec", x"34e272c7de5bca01", x"af6bb90d76910752", x"aa28d5fbee5dcac9", x"00a01416f02808f7", x"99bc163fd8f507ce");
            when 23306747 => data <= (x"fda7f64c15a9a5b9", x"d2f2bd5a16019db4", x"67333312faec434c", x"41d5b3462986648d", x"06648858a76588f3", x"be0f42905279a2d8", x"78085e6eba9ee2ea", x"a8745cfb73d18b73");
            when 8879275 => data <= (x"15103f493031f40a", x"0bd7ca09f2bd962f", x"253b5b5f44f89957", x"f43af7d61c044f14", x"b75745e10fea1edc", x"decd7bddd0810d4e", x"d5dba854d2059230", x"23468eb4bbad5705");
            when 29798404 => data <= (x"d6565f6bdd4faa4d", x"8c4578dd7e4648e4", x"17e3cc8d2bd1c043", x"42382eb341d1b077", x"b00db7c04fef2dc4", x"a3c99f70ac93797b", x"3cacef27ae2788ae", x"5b6a67130d01d29b");
            when 12030857 => data <= (x"56c4177b879fde3b", x"e04a0964100b820e", x"0c415b0d1d0f62e6", x"2ffec67af23d1324", x"adefed1985d8ac93", x"414bd5325e90bdc8", x"0f93f62bad7e558c", x"bef13f8b9f07f579");
            when 26722248 => data <= (x"9583711e9e0f7822", x"ddc23213dd95e646", x"23cd7ac3df8f9301", x"8db9300b6b0d8b29", x"2fe31ef3f944858b", x"9eadd6de60180fb6", x"596737f858a8ea1a", x"f23ee8f7c224fbdb");
            when 26020194 => data <= (x"9840d84f573da237", x"cf8e0c0fff523b4a", x"674875957372ff1a", x"3ab782f87af0584c", x"f0d535a7ecd55407", x"25f21cdf40f74ed2", x"be618c9b274f037d", x"87e2d9cf5e46094b");
            when 2332419 => data <= (x"0d026d2bc1386806", x"18b836d862b3a322", x"5550f0abcc924aa5", x"665f73c386b925c1", x"79521dabdc9411a3", x"0d80b0febd71fccc", x"7b1975f785f98a48", x"1319def1a4bddc9e");
            when 10912400 => data <= (x"6952c30759649091", x"965975655add1263", x"c7e6cd8543a41fff", x"3cfc8407ade127c6", x"97d071a4e313e166", x"06e8ae63e96557c1", x"3dae4574568209e1", x"ab3578dd223e434f");
            when 7447128 => data <= (x"d328638a042654fd", x"f8e260bd0acbb827", x"f5d9dbf14708c74a", x"8f266c1668cec7e1", x"4640748413b65970", x"88749b0628839d57", x"e76211bb9ec6c77f", x"7846ca6c2cb00059");
            when 25416043 => data <= (x"01f8c2b695064225", x"e3cc4d84f3ac750f", x"d33198876783e660", x"9917770dca4af220", x"e3267d5b661fb00b", x"37e6f37c78818bac", x"efcdff3b8d96bbc4", x"99ce6c6c77e3290b");
            when 5472160 => data <= (x"3292ee85d8a7ef3b", x"ef9345bc28c56bbf", x"40ab5fe87d311a36", x"5652c6084bf39b68", x"0de560fbfcd4472b", x"cb9d1604f56ca337", x"4127ae3e6e96f561", x"70951a705ae433b2");
            when 2042111 => data <= (x"7e7b93643eac134d", x"59d2a918ef4d1d68", x"0d79778b1593c295", x"ea61d9c41e0878c3", x"372b47c8e7e2cf6d", x"7c5c0233ecc9cce4", x"ce4d54c5145e24ae", x"2b2a41ec69233341");
            when 20500207 => data <= (x"9db506112b18a89a", x"d6e5d4d1c62d4a77", x"d5c37aa79fce2f8b", x"4071e175c607938f", x"9ae5b2d1391d09bd", x"213c81e5ba575436", x"9d688a5bfbd3738d", x"31cacace0f64a9e4");
            when 10886038 => data <= (x"5c62ddaebd982747", x"ded5a0ee0cbe72fe", x"031167aeab3325e6", x"af961a86b87e2c77", x"70a5fc7aa6c3fb48", x"006414c463011c27", x"4b9145cae6fba519", x"ab4781dcba679e91");
            when 22224290 => data <= (x"1d8da4043ed08f70", x"926b79afc6ead53f", x"795b970194cbbaa2", x"f043418d31774055", x"98e51042dd396a89", x"75dd8b851a0d6373", x"33936e52e5c80ae0", x"0514fe47afae54dd");
            when 30784918 => data <= (x"d79c32cd4dd10f25", x"c59bae640b27e370", x"55f7e78fe60cfa1c", x"e7082267678da3cc", x"c6f027b9f50d2f1d", x"ba3659d1998b532a", x"a40ffac2ac0b9421", x"ac5449957213e2d3");
            when 12161187 => data <= (x"88a5c2315f7a04ed", x"6cd08f58aaaae2b6", x"9b1803ffc7fdefb0", x"f250129f9f72d635", x"11f85a808faddede", x"2b5cada637196011", x"0065937152eee691", x"8c3a7bd8279272a7");
            when 10184894 => data <= (x"c3f6ea446c6ccce6", x"38ecb1fe7eb99f20", x"c9b68b368579584c", x"c037c2b54fdc4cee", x"ed95150098781b17", x"def1c077a12d1248", x"3d957307a777011d", x"01c2957e9806a93d");
            when 30161783 => data <= (x"deb0209b36310c4c", x"0ede9437947aee6c", x"bcbd7b1e3d73ff6e", x"1398cd42de949e7e", x"e9e91e68d2b746cd", x"3a8abcf01d241822", x"25db3189b1b7c1c9", x"cb6463222f367824");
            when 4012996 => data <= (x"01fa0012d66738ee", x"ff7a34db85f78c4b", x"b4dbe682972e63d1", x"13e4614ce3e3438c", x"5332d88b3389386b", x"dc1d161b396c62af", x"36e0b7665289433b", x"68780776c2051dfe");
            when 20971856 => data <= (x"2ba351bbd9835f91", x"a5b1794390aa1fea", x"fb6d9374a91ed059", x"341bce1adf14129d", x"9151f33545773c46", x"8aa9631e617d9054", x"cc0597280f298c2c", x"37dd9edbc4632040");
            when 14874552 => data <= (x"c2ae74b7f3ea1ecd", x"c0bd031becb51d2e", x"5b2a6615cffe8e9b", x"6d0e9a9a8a6bc61c", x"4862ca93e55e71cf", x"544308c8838d2d4f", x"199e9b9e4b6ca131", x"fc308835b01df63a");
            when 25388020 => data <= (x"e4f5dd06290450a1", x"5d790dfa09f4996a", x"54311e4caa3b3bb8", x"928b3de6ec75617f", x"7b75f6390cb6ad2c", x"5e291fb8fc4416f6", x"c2b4de32974144a0", x"68057a15bbd6af70");
            when 6671481 => data <= (x"39d7d7d3c7bf3ece", x"9def3e207a47df1b", x"27f22784332749fa", x"89019beee1ac25f7", x"c8e83c60bf23b421", x"3dc05ce34c6abfb5", x"411f398ba083f457", x"d72d2572aca90983");
            when 20963319 => data <= (x"5ad3d5cd491cd91d", x"786bf14aa1d4203a", x"03b87836ed3e6e77", x"3c0357c499ebdead", x"22be5eb737e9f78a", x"520bc6d5b1f832b6", x"f46cba873d3098e4", x"12ce14f8cd06e096");
            when 32154023 => data <= (x"9dd051a0cd78a36b", x"4c0213b332bc930c", x"2d21a9324decae5e", x"d7de658cee690bc5", x"bb5f29e514c08183", x"f3d7b98b5d436dac", x"d04966d99b7d39f7", x"c71db2a0fbfc7bdb");
            when 26774136 => data <= (x"5b5c21ca2897d125", x"259e7c104dd31c17", x"5f4f46947b6b4808", x"138a7792edbb81ca", x"bf0ab39339c11ecd", x"d8cb1def2e8fda21", x"3bf0e21aa562b54b", x"43827d378dec7c26");
            when 24685574 => data <= (x"7fd75e38cf8ea431", x"46bde0feb36a92ba", x"f8562a4bce48face", x"7466c9464326ff00", x"d64074664b49f542", x"d48637a5a80d3995", x"0d6f8e065b07fe22", x"1443a5da4a63b409");
            when 14365684 => data <= (x"bf5aa73b1575ff5b", x"5163cc1fe7145183", x"c54961c6c7d5fe4b", x"6796c72d6d2d2a7f", x"6a544fdf21665f96", x"ef256b89d8672b68", x"08d3f1f189f644de", x"6117339df615feaa");
            when 20002302 => data <= (x"32fb319ccc39e26f", x"7560d976b6cbf962", x"e48c8d7efa8627ec", x"3af8f83a6a125113", x"a8db4716bdbe2adb", x"d385e2801039dc85", x"4af4980ecf3fc2be", x"316746979f7e4f2e");
            when 23643789 => data <= (x"850cb6b3700e28c4", x"6cac0057ca8e09b9", x"2abd961fdac629d7", x"6627f174bc8d133a", x"77896b405b121942", x"19176a74f7e4e3e7", x"a0bafe1576d1d016", x"48ab50645c4d6128");
            when 27824316 => data <= (x"ab1d30c92d6cb197", x"695fe1b808952672", x"f7a247d13aa789b0", x"5c3c9f2da29fef49", x"0a304c5536bc3f77", x"a646e9f28029bb06", x"5a309b7f59627ca0", x"fb1fdbe0b109ae7d");
            when 6982760 => data <= (x"79a41cf19a46ca65", x"616de1632e9c82bd", x"4971363bd146d43d", x"fdba948f2786bf0d", x"185b6658647820c8", x"950e2bde20981e54", x"a01cd38399aa0092", x"2c4dcaee3ba36424");
            when 24206833 => data <= (x"0a817e700c8d3e9c", x"ece1bbcc26e59e5d", x"c9cc5455b295413f", x"14794852e28a7229", x"1d25765820510118", x"6eda73d325d6ceb5", x"eaab21c3386b8305", x"8d39bfdc1d4f8508");
            when 3663577 => data <= (x"ed13354b16f707d4", x"99ee7012385dae21", x"aeda419ddc15b4bd", x"c7fb81f602a62129", x"e6fce5d13e4f0688", x"17df03c5fbfaf4a7", x"1d218a38276b4c56", x"9f7383ce86e5e449");
            when 16845207 => data <= (x"7f75a195d916f6c3", x"4033f19e76dc656b", x"d460fcb0b4362b77", x"201717a2bd831e6d", x"562c10d6bb8ea2f6", x"bef63dbe21380b49", x"0487541ed543631c", x"89c77125e2bce392");
            when 13529007 => data <= (x"a40204e6a452c7f6", x"4af431d719690a37", x"59a5bfb6a829b1a4", x"18321f5708ccb2b5", x"e3768b51c76a21c6", x"e3dec036336b05cc", x"a3e34a956136b163", x"614e86d483c8ecc8");
            when 23100622 => data <= (x"def58f882aded957", x"1bdaa98284be4008", x"7aa16266257b5f7c", x"840d55e56f71437e", x"5eaafd1e433922d3", x"c603519dbee16d62", x"23706edf4d4b5abd", x"6504e4925af0f84c");
            when 32395759 => data <= (x"c5f607b8bfcc585a", x"b3326e8425c1cb4b", x"fd085146432c80a7", x"a9447c69814fb998", x"9f4cc7b81db87f1d", x"6bbd2817358b0e2e", x"dd37ed6431976072", x"d57d5198d0d4b36a");
            when 2044282 => data <= (x"c79c40a6674ad3c4", x"d541f32db6ffccb9", x"274e18e789e651e9", x"7255c756d4efc88b", x"d30702645cd41f3c", x"48cfbca2c2306501", x"25806450d54d3db5", x"f43056919d329f4e");
            when 20519945 => data <= (x"21de094fc751d8ad", x"e5fe3e6e04986370", x"696e417a2bc240db", x"47c0de3c6afc6a8e", x"7cfbfecedf541f8d", x"07d0dc63a0b1a174", x"af6b4730098864c2", x"db6816f1fb214f94");
            when 14718047 => data <= (x"475f6eeada6d6e60", x"0180a89c6b92a5f2", x"9a9532f77f0cdb88", x"2d4e0247bafa7a0b", x"668e4231faad5144", x"6e3782458e0f5691", x"cc2f5a67ceaedff8", x"d6a8949e9ce40733");
            when 17882178 => data <= (x"2c22ea0579dde62b", x"831416c119098c27", x"932f49b18ed03be9", x"2242bfba3032f9b2", x"a1cda4c853e723ad", x"13e366c0ed80ec30", x"0ad544c5f170d0d1", x"9baf9235b3f71886");
            when 2200577 => data <= (x"d6af1068410a1643", x"92ea122279141d83", x"2c0b0a64f1250bcc", x"b5246f72bb1322c9", x"4b7c436453e567eb", x"de557c0db2ae0381", x"d6822208cf36d0d9", x"1450a112c4693bec");
            when 23742516 => data <= (x"a8fae08cd9c13153", x"630b6768a0eabfab", x"3f34d3f9c0e6558c", x"6d139aa47c375cf1", x"076fe7dc2558fa80", x"d6dd4e8501274471", x"8edae156df751ab6", x"1a76cb7c07b94d05");
            when 26859910 => data <= (x"5e47182ac22875c0", x"0b573f10607c8a55", x"db184370104ba5ce", x"e460ce54cacd3596", x"d30828317adc50d7", x"5d1bf4722e5d3471", x"c4ad458c9868571d", x"75113a42e71a9983");
            when 15864606 => data <= (x"c826e9b0a6554f4e", x"372903129a3cceb1", x"235bc856ddc7c47b", x"839d467d2b95196d", x"d4c03238db2f342e", x"dd3198af9821867f", x"5900ea0681227715", x"906b365db21234d9");
            when 9534380 => data <= (x"7797d997b30892fe", x"11198ba18395ada0", x"41a054bbee2fb974", x"63fbd7174d5c811e", x"d4819731e34b2e7c", x"f9b94d8ee7ef94b5", x"7bfd3178af86cdb4", x"6a84fdce6e042638");
            when 32570851 => data <= (x"4ba033beba236ff1", x"a408c7c1affe0d61", x"e42b996d3ae73c80", x"894db1777a0b07a6", x"b0fa9b74c0114d25", x"e52c02a0423688b8", x"d6785f270a81a46f", x"9d6ef41b04154b8a");
            when 22383937 => data <= (x"58ed5564332b84ef", x"6e04b47aae0c11b7", x"6bbf24e0593b0065", x"460a7bc81df515be", x"cff14fb936322ee5", x"02fb71c3284c7866", x"915d499efb4129c2", x"9d320d8c95c67fd0");
            when 17823460 => data <= (x"58b0d0f36a310c3f", x"bd7aa360cd3f2337", x"b4f7cf57485150bb", x"c387cfefec1001a6", x"55f1f927f73e81d4", x"8f25e6fa3fef4c41", x"adb4c2fa272e1da5", x"3d40d6966f4fb5ae");
            when 5388353 => data <= (x"aa9ee59cd2c2463e", x"311cd0fc7f7ffe7e", x"8ff4ccbc9d146ea9", x"f40c0a2e60c6a327", x"4d6a412482260908", x"4b6247972f31914a", x"2407e511c0918d46", x"8b701d2035f7897e");
            when 10121283 => data <= (x"66cbafc961e8ac75", x"47d3d3e9e5424a65", x"2e41f4fb353c0c8f", x"0ad19e3cb8336208", x"b094aba25a6670cb", x"6e35c53270ca5b96", x"8312315a8412d0a4", x"408c1bd592f1fcf7");
            when 8398778 => data <= (x"2e4bf57ea18a99a2", x"8c6e44d69104b9e8", x"dc6974986074c0d0", x"f7f33c2153d3a25c", x"07ec19c3cc2c0f40", x"a46ae003949201df", x"5468556f7bafd6f3", x"bac53689bd2404cc");
            when 16617594 => data <= (x"4ffdcab40ae59a2c", x"7082fbd32d830615", x"a7148d868935ecdf", x"93babbf60cfc246e", x"c9e0a0fc9902749b", x"e00271de71f1d99d", x"24a2bf2bb413e568", x"b166e8aa761d7c74");
            when 25617698 => data <= (x"26eb5a9b08a01772", x"9c56781e3382ead7", x"a534121007e0c990", x"aab6227844d2d994", x"edd6d4205bbd8d5c", x"fbbc6773190007bf", x"3844efb6e0d2c8b2", x"69774274c9898eb4");
            when 21866512 => data <= (x"58209d60d4e1fc96", x"19ef78fbacfb969f", x"78fc385a4bbd827f", x"728e5d614cb3369f", x"9a1f35dd31cc61fe", x"142815e2d79fefa1", x"7dfb97dba286c687", x"51203ed03bb11afa");
            when 1697049 => data <= (x"73a2c89c396a5fb0", x"bafb0ee6378f011f", x"e29ff88445ab3c61", x"8451b11dcba4ad09", x"3f4b99bc16f51654", x"5f55adffd407305c", x"a871de335a5de3df", x"04fd040725446c15");
            when 1367440 => data <= (x"0228ab3d2d58729d", x"64e3a143ce802bd2", x"e8fbbcf7425ca545", x"217cb6e9c6d2e170", x"a5f42550a6fb5eda", x"d7ded42c40e22f3d", x"8fcdc8d9a55a61d3", x"4629d2a2f111a57c");
            when 24023893 => data <= (x"6b51c602ba70bdbd", x"814e71a30a641f86", x"64366182cd43fa23", x"7ff617660f6302e5", x"49a388bdc635adcc", x"82b47ccb80d4a824", x"97b66025f01fc1e4", x"f304e46204467498");
            when 16041657 => data <= (x"320429c2a19e722e", x"ac458252c39a8118", x"271f6b6cccceac41", x"dfc990f7bf8ba44b", x"afaa21b8d00a4baf", x"b85c721d00f86aa5", x"7409a5bf20bba5d3", x"e61551b6b1fb84ad");
            when 11693158 => data <= (x"fe5ac24781e9bb7f", x"a3ee1419eceac560", x"fb122e36ad787839", x"af37af361261a1f2", x"0b0b069f2897c562", x"ec55ffa1242fc178", x"acf0277bb6c4de9f", x"62475fe51bcfe433");
            when 23237968 => data <= (x"3333b674c268144d", x"345101ba9ed1df91", x"914f193c744b5c83", x"13a9529e8752432c", x"628f92237fac98c0", x"2b6abcc158d2f871", x"1522730ded97559f", x"b32f350081bf63aa");
            when 15142134 => data <= (x"54db51a4c4412923", x"930097bccefa6dc0", x"cc2b3a092fc44382", x"ae5d130b7ba3ac89", x"76d6eee6da3f1810", x"7b7c8d0265175542", x"0f2cac7c29cc562d", x"bb4b8c9cc7f3667e");
            when 12798362 => data <= (x"12d83acbb0081a3b", x"353ea42010961c9a", x"f29ae768defece9f", x"54a7d0f8904a548c", x"409ac1346f46a73c", x"fafe611f45012201", x"2a929fe793010a40", x"adef9c8293a14c5f");
            when 14312403 => data <= (x"ba137a8a1963393d", x"251abbc2bb69b8a5", x"046d9d2ff5f935e2", x"761beaabf04dbf19", x"f17b17517390768c", x"7d4b9833a4c3ae5e", x"d320fe5251b8110d", x"554ede62457a9e65");
            when 28513502 => data <= (x"6647e40be0eca293", x"33a27f8d8655bd5e", x"b7d50ff47730745c", x"6ed74b7f12fbcb09", x"9c64ad7be37d8f6e", x"fde7f9ea3d286fe3", x"59ae4ff5d8198837", x"b373b3296d6a34b7");
            when 3728759 => data <= (x"7fa2f08f9ffc2145", x"d9146e86074a9046", x"c1a20ee76b4fe1ba", x"4acb729a1e5798c0", x"81842e6d8fcd0991", x"0be432bc3a50f678", x"b4b8e74a8ec51020", x"fa82bb2be3b357eb");
            when 28555062 => data <= (x"8acd4e1d330b612a", x"0348b7e4eb280dc3", x"8cf236f66ac17970", x"a6b936bfd477b0e4", x"207e6ead2b55addd", x"134d1296c94c4506", x"ca6259b9bf730362", x"5184bc714a0d59a7");
            when 2169822 => data <= (x"4a8c0dc8b8f40313", x"6c28dab3519cae2c", x"4026818be001730b", x"f7869670b4f9ba3f", x"b2f83c758b657a68", x"9f7023ad71b51b2d", x"c5426f962371d0d8", x"6df70785b4e610f9");
            when 26135215 => data <= (x"5c6d10a59f44f96d", x"9deab230c74fffa5", x"c4d36cbc5d4f7b19", x"a9d16bb1fd2a7027", x"780a4f42a83c3a3f", x"e6f4bbfc7a5b591d", x"22dd37a67a0847f5", x"749e611e424b8ab2");
            when 21173409 => data <= (x"00567ca1dafb925f", x"9fe596ff6196eb3b", x"a2a0f3959d9025c7", x"8dafe56fd961b0c5", x"6b2dc2f23948361c", x"2d5895dfcf5c3201", x"9bdf462bb88d09b2", x"6a2b200de4a52a5a");
            when 15083967 => data <= (x"65cc906dc9bab70b", x"4e40c948eeb3654f", x"db17b717fd46975f", x"8e93171fccc2eee6", x"9c3558d45ae7a8e5", x"d7563205af6b9b79", x"523806f506862b19", x"cf35db6dbea6f3fe");
            when 31614754 => data <= (x"a043deea1b3e1064", x"9fbbc637843bcddd", x"e55603c143b96265", x"d88f3aa24418eb7e", x"8b45576cf08a079f", x"5adfdfb0ca311250", x"1105a3bb34992af2", x"ce1343856d3c1d10");
            when 27714721 => data <= (x"c484ee05306cb188", x"bfca1b2f9f45adaf", x"9df9133530d0ea48", x"cb4c371e56bde86a", x"e7e7eae105d3d2a8", x"3972d117e84bead4", x"08c337f04da0cc0b", x"066aef42723c3e13");
            when 16697683 => data <= (x"700610fa1f93fe72", x"4393f3240048019a", x"cba79bc4d39505c7", x"d824a7b289e57cf0", x"0a9448698096e79b", x"aedadbec59056443", x"d44921cf6cc17367", x"f5e26790c8e958c8");
            when 6394681 => data <= (x"260ac268753d1111", x"db6bcf8a476aae31", x"309206e7ebb7eab3", x"e8f404601dbcbbc4", x"206bea69cd60c71e", x"03cb619bd0f24971", x"ca47f68c102293a6", x"3986072978dfb415");
            when 23510899 => data <= (x"4fe3d20d01cb001e", x"624c38c316bc6b73", x"3d690bd40e3de4bd", x"3852104c403216b1", x"3a4210fe6b8a4274", x"b20c6ed86ed459f5", x"00812b52f7288920", x"2e3742e0252c0d20");
            when 31070548 => data <= (x"c12a132aaf245ea1", x"3d9ac5e214c5f078", x"324d62bb3c4b013b", x"460cc16805e6f8d0", x"68491944847776c0", x"559f0508de433042", x"60120b170a064211", x"f2515af2128d31c0");
            when 13212708 => data <= (x"7893255adcca9db8", x"25fb4b6a141e0946", x"232b85ad72ee3595", x"a6a7e32fd9e74ef0", x"783eed1d71d08ba2", x"ad334e85f2bf7d9c", x"60c180c8a92f26f5", x"b0010d9fe5800c81");
            when 14198694 => data <= (x"64a437e11c4bb8b2", x"863958c7ec7c7ecc", x"14463d762de47235", x"676be9c318f913b7", x"7c5b5963d1bcad26", x"46a653ccd1f432c5", x"9c9c772de68c3bd1", x"08d2ac53f3b0c7a2");
            when 8712136 => data <= (x"35a0011302f1470c", x"a78bf3cf701d5df6", x"0d9cb60f1cf6e464", x"8d19683f7b02be2a", x"7e1ca735c462a73a", x"d75aed6e16432a14", x"fd24e145bd5de2a4", x"17521fce464c9531");
            when 21678046 => data <= (x"24c0413bbb68b3c2", x"b56aca1c358a587f", x"adf377a133ff99fd", x"590efe1b3437d72c", x"d928a02e6d499e3f", x"ac7693c1b0a4dd2d", x"7553a4f57a3858f0", x"164e85294f6fbf84");
            when 19428076 => data <= (x"90c52f8e0f063ea8", x"500cb2644e22d078", x"0354bd27b63cd8a9", x"2c6c63c312728f51", x"dcbaa8eaa7a84e8c", x"f64ce8b12a6a9210", x"2e4c65dc14810901", x"e81915f608fbf038");
            when 11414231 => data <= (x"af96688a1bea8880", x"f6d9115bfaa68139", x"0351f4c1bde39a67", x"04c653edd9b4b786", x"8acffcc124bf9713", x"426328eb43e56ec7", x"038a7b8c9fd7cba6", x"15c2970419c64977");
            when 25304644 => data <= (x"69a857b6f30fec7d", x"94781d982328b29d", x"b5f2a7b0dcd22f65", x"3661cacaeee1cb2a", x"3d53b1c020d80dd4", x"811db06aeab4af63", x"1e37ea3f0d6a2446", x"c7f16bc2f90bda30");
            when 31811673 => data <= (x"bff2c89edc1bd877", x"7dac37de9dc877a3", x"44d3fb1dcdf9b27a", x"13817aaa5e102fcd", x"7de25d70141d5942", x"cb3037fc55dd44af", x"9f5669f2c64b5e55", x"01546494fef4a913");
            when 24154501 => data <= (x"672a86ae81cd92b9", x"43bcb8ba2c3a5274", x"3ac74c3b053538bc", x"b9dcc5c788076b0c", x"314ef792596135dc", x"68c03aad2cf71711", x"3e4c7298e640c503", x"017ac3b9a67fe728");
            when 33081718 => data <= (x"88fb011b7e08e794", x"9dec1c3c105c9f52", x"8a5ba9eac636720e", x"0b439e59bb3a0268", x"554e86cf7cab8f8e", x"9029a3b7a84af133", x"ae4e4be4d6728e33", x"0c7f16e0864a3afd");
            when 15868538 => data <= (x"f82ebbe9ef439026", x"338453c657046994", x"3e08daa382dddeca", x"036b96c330d6eb0e", x"d1375036ba7d25c8", x"369dafba7affb69b", x"46d783b998ba2c48", x"7dd32bc332434c09");
            when 24329763 => data <= (x"d0b6d070da5c5789", x"11109561f971f58e", x"405d101c137d6a59", x"a219c4aef09cd8ff", x"89f79db8037a0459", x"df7424cbf3870de1", x"dc0b141dcbcf0173", x"497a6cf1ea4ff3bb");
            when 5060505 => data <= (x"3fa8c4bb7cf2d311", x"f6d7695cbf07073f", x"2ab9d0316e9813e4", x"eb93f17e80843b07", x"b5343025047a3c12", x"97df0245da008007", x"c603f12eb46d606f", x"d90c5290b3449b25");
            when 31984489 => data <= (x"862c78ba94582654", x"bde7582ac6b20531", x"bbf4c51fb8e1ea84", x"b4c8d419267e97be", x"1452c1696d979199", x"176eefc82cc21d2b", x"66cea67fc4704b47", x"de9b3f100fb8423a");
            when 27777742 => data <= (x"f853ee15e8b37832", x"5e0f2ecb2accf575", x"d0ee0e2c8aebf12b", x"fcde0568ebfcb058", x"4f1d147c29ac2bfb", x"c4e3c2d4603168d3", x"89241557c54d9e5c", x"f364482c61db2ae0");
            when 18155033 => data <= (x"f7dea7608d7b815d", x"d3e3bc5030cba869", x"b0612c03732ea096", x"97e6ad6cff9f0c39", x"f189fe1bc1339515", x"424a17d6748dc3fa", x"236f0539506d746f", x"a09e9403514f5d9a");
            when 1684067 => data <= (x"a34087159e66d0cb", x"f898cf644fbeacf8", x"37b03996a5821c86", x"26e1e18d52fd46da", x"d9a2e4cd1b914f01", x"1bb083eef8de9c6d", x"4f05a2be5a644d25", x"44287963c3d0839d");
            when 16012488 => data <= (x"e4a410169aa8e208", x"76cb996d62903dbc", x"2256d6943955fe97", x"2735146ea3273ac9", x"715f0adaf4b4a873", x"bc05bfb2eb59d186", x"ec5984db520dbfa9", x"ed3989ed69c81fea");
            when 18886896 => data <= (x"055be6106c5086da", x"058b9e73b44b14cd", x"2e1fc27af286b564", x"7a3df55434ab5d93", x"423450e24ad296a6", x"8cf3054b0a75498c", x"285a235efbf6f473", x"6d42f008514d6905");
            when 32977248 => data <= (x"03b7bb54f7cb9c9a", x"349ed7face781289", x"9e5e9b0b442219a4", x"10f386f91fb0c95a", x"06bf1cc851ac4730", x"e2b9882b29863d9c", x"bc860ef24d657c94", x"a8bb4b0eabe06d96");
            when 28108117 => data <= (x"5dd67e14a067765b", x"d48808ae7b9272a4", x"2fa30db0780d618e", x"ed9f88f48a6abd42", x"ac5cc1f6c100fa0e", x"e85de0c34b1e0609", x"036e1d3e61b0dff8", x"db01fb832fee4438");
            when 1270941 => data <= (x"6ee10bfd97b90ec7", x"b3262f9f895ff7e7", x"674dd72afd642ec8", x"bc50e0fbd2df9632", x"3fab8723255f2cfe", x"6cde4533a7dd87d2", x"687838df4602c262", x"1b247fc9421bd083");
            when 29476041 => data <= (x"0bdea64121fd7c01", x"70d401fe09144263", x"620530d6cb691079", x"e4b58be1c8af2f5f", x"0c4947f388e16569", x"1340030151eff724", x"c8c2599fe6c7f09c", x"76b555a9b5190ea6");
            when 30686153 => data <= (x"0fb65c318478415e", x"bb81ff13cb059971", x"2594f2d4584f5a48", x"9ddc21e4054aabb6", x"b715c8e2d15b63b5", x"e4d1dbf5625996c3", x"246dee764b7df958", x"2f647240413ae3b9");
            when 6705052 => data <= (x"3704effae92e91ca", x"bef94b53c7a141a9", x"c2f1cb72039b5a1a", x"d64ba5d30af67122", x"499bc37f9ce6e31c", x"ac4613d425ac2999", x"c932c13ecfd71da2", x"73ce6efbcc449c95");
            when 11075817 => data <= (x"c20890885f185ade", x"5635c214ca0816d0", x"0e95a627dceae18c", x"0521e0db5b017138", x"cb7944f253544386", x"43fb2d5142e08dfc", x"d43365aec67312fc", x"ed04dc20f5b1149b");
            when 23296896 => data <= (x"007282f682d43a75", x"766a0812bfdc8165", x"137addccf6bed526", x"38da4871011b99b3", x"7581d0c7c7f45388", x"3b9746032d6bdf98", x"164cbf1c766978eb", x"074e27e4dd1354ce");
            when 3502639 => data <= (x"1816becb79af7b50", x"38d1611a534d9ec4", x"ec6f6094f12e642b", x"94991ca2247082b7", x"80f103f7277f2a1c", x"c55e3dc8785fe748", x"345f9ba62e4388b9", x"c6f9a2713ce50b20");
            when 3141338 => data <= (x"6ad5ed15a0ae0c15", x"8ca35a6eb73f7944", x"a9cd5a44af904979", x"fa9193af7d0c53d3", x"84c6e8e6451338bc", x"551d3ab41d0212d0", x"264ecde1296317ee", x"71eeedb8893ac53f");
            when 17727290 => data <= (x"8a513a177ba6194c", x"c72351910751d16c", x"1cc13d58a3f4dac4", x"0e11de56f54b8601", x"83f53753a76bbc13", x"b3c3e72201f3df31", x"c40868e697ebe80b", x"c73f3642894e9c13");
            when 4393380 => data <= (x"bb06e50fa3c3f899", x"a7984f5c8737c491", x"8249d0269eceeb8f", x"02960d250bdd803c", x"268a6c23783f8340", x"60eb4e699763c235", x"eb08f7415f0e0056", x"14ff00ad7428bf16");
            when 16274257 => data <= (x"9ceeb5df4bc39b2d", x"4cbfaa0cf7616ee0", x"082594424c0a7641", x"cda049085e2a176b", x"40e5dfe3ee542ecd", x"f01dec6d411ce1e7", x"a5580ba68e4b1b42", x"46ef07f7167fe8c4");
            when 24019485 => data <= (x"cfd3f34f13fba86d", x"f8a213614a3ca6b6", x"931160495b898d5e", x"230855ac41a6976f", x"3dc2204e9b0d9b2e", x"2178625aa015c5c9", x"d8c1b8e84f34fcd5", x"ad94c1589e0faa78");
            when 8329740 => data <= (x"35ca1e0833767ec7", x"0a078510731a1c4c", x"bd244243d8492769", x"fdace28e94430027", x"8385e2617c177e97", x"735496417e4740fc", x"7c43cdaf646b2ffe", x"fde9312c7655d49a");
            when 20200450 => data <= (x"97a6a3b2aaa2dcc8", x"9657a3737fb76539", x"3a3ebe7abea81635", x"743082173fdf5599", x"6ba2615cbaca662e", x"a89aed593b1b21ed", x"21aa2a6e4b802a99", x"e8f65bf3bf52ce86");
            when 4705380 => data <= (x"53e3f6f127b82d86", x"8e0e61db60312353", x"d9dc291a1f846f26", x"68458343cd7c1472", x"dd0e62bab012ecd9", x"1214c22fd986a00c", x"259f45bc43e14e0e", x"ecb88effb92709ea");
            when 15464669 => data <= (x"b03f7c83a6af34d6", x"c70dfeb6a40e6dca", x"b5c7fb1721d6004a", x"1feca65cd36eef7f", x"e9b70ffeceb04779", x"6164f12016a1bd7d", x"12f275f7f4577229", x"8c3485f101e23e33");
            when 26170937 => data <= (x"0385a455f976def9", x"58319d510a32ae7a", x"0a0df90a975d9d84", x"580625f65f42dd16", x"d314b6f24e67284e", x"aeaedab937a12e91", x"400c0273506e43c1", x"836724f1b5f0ee35");
            when 2455192 => data <= (x"7520a25996b5e635", x"78491485955a8aa9", x"fc32f08281672baa", x"e99fcae8da557859", x"16aa17bac257af5c", x"bf8e83397d8eac06", x"4df490f53196b884", x"573a6f96af9deec3");
            when 5845936 => data <= (x"eb141ad87f5ec525", x"7b3e837f1ea66a74", x"1bcc537d1b5a6833", x"8d6a8362171d3eba", x"40eb54dc1222d759", x"db9b10cc80476c75", x"f9ff74dc052c3d54", x"593f2a55793e5aa1");
            when 5079025 => data <= (x"a18beb4450359058", x"52943db23a918b84", x"b98dd293d7b12bcf", x"e0407c110ab8ccb1", x"c99a08a56ffb1f0e", x"5c32c52085e7750f", x"f54e4a00e40b5e74", x"8b07e03bb04d8cac");
            when 22003753 => data <= (x"cba0c10e03d4e70f", x"617d4245481478bb", x"84bf30c5c0caf607", x"171cea94f13d44dc", x"a99f6c388a5c0845", x"064fce0222a88aab", x"5ab2601e5938963f", x"a1faf3f8c270eddf");
            when 567266 => data <= (x"b4d27ffd7904aadc", x"d79c91c5a0b1b390", x"8907c79b61914570", x"9771bcb21b64925f", x"e98ba3e6ac6a744c", x"30c51344b8df642a", x"a5805ac68c919600", x"755cdae74a3441c6");
            when 10242501 => data <= (x"e595b44b999493b9", x"7302209394052623", x"1e7847b255c66515", x"e694f048cddc15a9", x"16239cd8c85c05dd", x"188865fb5e816e51", x"fc18b7ebe9195b55", x"d7a63433907cbcaf");
            when 12090000 => data <= (x"f0196a83cd2929bb", x"92d7577878835a2c", x"f8c00a706387cc54", x"fcfea052bb45140c", x"327a4256e8eead8a", x"eb23c220324eee99", x"73acedc4073cdb52", x"079b06ee8c3a7570");
            when 10515707 => data <= (x"9cdca16c9b4a1006", x"ff4302cdd6dc134a", x"ccdbd3687afa8bec", x"c690ea6aac1729c6", x"d251a11b714b6471", x"056ce6b1f0702fcb", x"d8e37196a920fc56", x"9d05a8ddc71bc5ef");
            when 12894767 => data <= (x"ce7178f0a75434ec", x"dd8a228c71dc5447", x"3f3b3c1af3363903", x"0de9d8ac26536b34", x"96a98b4c3eef29ea", x"dd65e7ad6dc37228", x"06c38bd870fb8a3d", x"86beb7e86b568736");
            when 12997647 => data <= (x"ddb442fc64230709", x"361d695d10800b86", x"1711dc6a7ffcd089", x"3a463a6828e0cc87", x"cb903660b915d092", x"5ea50ad551238050", x"7897e5400221c402", x"030af4053fb34dfd");
            when 11752671 => data <= (x"1c28f9cede7883fe", x"9cd2bbc3f607e8bb", x"3e5f941851e987c3", x"80c0c3225eb4fdf0", x"db68d80f18520971", x"68413a16e8bfc08d", x"3412924546798516", x"0ca3a5c4d1361ab9");
            when 30537810 => data <= (x"51c032c1a930f146", x"f4b232d15bf374a2", x"93a0911638571d4e", x"94e944da8445ffa8", x"a3cba44af587950b", x"838b7efe32a54d28", x"73f46ec1e2f9765c", x"09afe961747f0255");
            when 23516852 => data <= (x"545bb5320191d4db", x"06485caa71837888", x"41048b033947d836", x"d9a127f733992607", x"e0a30587b8531149", x"cde87f3092ad95ae", x"56052756152673b5", x"2d80edb3afb9860a");
            when 31460483 => data <= (x"b39f5a54e61d179a", x"3d0fcb24cf5a9404", x"4683d0bd94568a0e", x"a4aa30edd79422ad", x"42284e81aedbb51b", x"0f61f12f3e554191", x"a86a8595426b1173", x"67833712d91d86ed");
            when 11659399 => data <= (x"ec86e46b958fdc18", x"d0136842f5e09482", x"dd6613ca1b8f4900", x"7aff4c2194199820", x"3fee537bcf586202", x"9450a619eb8b99cb", x"63a11f5777f08d0c", x"ee6e340d9cc4b6cd");
            when 15839924 => data <= (x"32916bfbc2c36973", x"61e31d4444f5be50", x"f70827b15a1ba9ac", x"5a89f000ca01939d", x"3e5f311b4f08e4b2", x"4f785501937c4809", x"557ffc4365087b71", x"5c568c37e6adffbf");
            when 18318889 => data <= (x"614604d2bc19cee4", x"2d372e82906314b9", x"f65403661d38e323", x"ec072b22b6c81058", x"056ec52a3081ed73", x"4a9591c1b0719c3b", x"d00de9eb6042df02", x"f22337bd130f0cae");
            when 15684645 => data <= (x"91f268ad6a34fc0e", x"b054929584a13d3b", x"2c5341e0931a1820", x"168b3d45f5f48b4b", x"5d3e8d008889f54a", x"0c132a7f667174ae", x"63690f2de5d119fb", x"0d9f40bf9d02072f");
            when 8818838 => data <= (x"5a815c7ed92f2ac4", x"7c5a38eb669d5e8f", x"fed5d9ff8a27ec50", x"10e2b0481433df94", x"e7c13fe86bbe8c6d", x"03da7e771510253b", x"dc061a9dba501635", x"43f7cccffd719eb5");
            when 22110581 => data <= (x"894a1ac4cc16246a", x"3dc44d0dd21bdb09", x"798934fcb7248461", x"c707d94a3d7076c9", x"e1d6ded088fc0a80", x"bddce6de879ee63e", x"8a0a3bc550faaa3a", x"7255d290bd80d7ae");
            when 7122327 => data <= (x"b28f7a193ce18b2d", x"797a33517cdec056", x"654e8ff41295e89e", x"f6f1248f17ae9a3b", x"c1eafd75f639b619", x"143e278f58f977d1", x"16fff0d0299424ad", x"ecdb332d155909d0");
            when 24617247 => data <= (x"6f76625f891baa30", x"3ace403f20f4045e", x"9b3acb0d77859a05", x"88c82c05d882a5d1", x"ee8af1c3a098db5a", x"35e1c82ea6d4fa07", x"ec1c7604915ebea8", x"68f9f566094be4c5");
            when 16745802 => data <= (x"b28d4041d3c65bff", x"0aa5a605d069a66a", x"86ba7a5316fa3b4f", x"32da3f313c7db2ce", x"19457036b56e8878", x"02745bcbb12c13a9", x"c84bad98f4533a9b", x"c520ce102462773c");
            when 20599891 => data <= (x"1cbfa2d0bc650084", x"e8a78238d84fc1b6", x"16b9b5827ad3a2ab", x"a09ee0104bfcb5d3", x"521dc201e9ffd659", x"631b12383d65e2db", x"f599fa1afa9ac768", x"981647f306bd82c2");
            when 33153617 => data <= (x"a00c6c96b26b936b", x"cb732833b454cc0e", x"3700c93d4e885751", x"17eac1b0fbcfc306", x"f42ee2e1e766cac2", x"849c469384c804f5", x"1a2d49e2d123f040", x"f15ea2daa6578386");
            when 10751834 => data <= (x"0de1ac872bff6b8d", x"a07b4b16604b9f69", x"685b8b3595d5a084", x"4a016d3f3ccb60b7", x"cba5a5b0694c90da", x"6e39372abf44ac5e", x"bbeaff3dce2fe7b5", x"05111470c705bbc1");
            when 9969274 => data <= (x"95d6c5d24e7dafa6", x"0835431af95e2d1e", x"d69f08b812c0519e", x"e3ee6a946d252819", x"d0526e0d538eeb01", x"9d85388c3d05cdb4", x"08ca1797a061860a", x"8ce52db354fe81f5");
            when 2465343 => data <= (x"d3c7fb24bb2753d0", x"dcbaeee7af3f9150", x"86e9c0930a45735c", x"d7ec289d6d9bd125", x"f1bd137e1a856a26", x"dc9b513f19d2161f", x"298c18a928722473", x"9a928df5c2dc7c2f");
            when 4009002 => data <= (x"e7e7bf600ae3a5ce", x"a2820ed16274b63b", x"7b3a29478a593181", x"c52fcb2f3b6279fa", x"3c1deff1bbefc0af", x"6fba9caf653247e9", x"3a93f89cb9c812a4", x"04482e9a69897c54");
            when 12459878 => data <= (x"71ad67839c96e769", x"9a59e99b4fecfd66", x"eb3da4fbfd09950c", x"e9e33a7c066e2ea5", x"a1f10cc9364e73bc", x"d952753d3783df04", x"253fa4270a609326", x"4baa49d4e1a763d4");
            when 14537081 => data <= (x"689d88bea86be5a4", x"99afb6bb7d6ffed9", x"965ab9a495c7aeeb", x"d02a88058a6be8ad", x"3cdb154478ea5e0a", x"b2f043b99f22198f", x"a883600ee1e8c7c8", x"a8284abfbb92e691");
            when 26652332 => data <= (x"c8b9e59f5017141b", x"a4bce8d413817481", x"7ea23e3934713895", x"05760e8a26d17ea4", x"527f0c26b2156a8a", x"d9e18d9c6423f37c", x"0b925939aae18ae1", x"c601c63ec713530f");
            when 648853 => data <= (x"ae40671846d75cf9", x"128e0b742617650e", x"f67739b2e433f55c", x"8bc44722e919e649", x"899b0f6ea1b5a118", x"81b7865bd3419bad", x"d9c8eeac24a8fbd4", x"255c5ee52dd2d87d");
            when 32128285 => data <= (x"36e5608bf66d1fcb", x"098abce68def23d3", x"c3009e868cd4710a", x"243f426a731b3196", x"0bc0b7cfe5799ffc", x"b9de3d2c0a13e08a", x"079bf4447613ae71", x"0a9af9bae277347e");
            when 14776354 => data <= (x"8eed70bef162e37b", x"86f21d8f7b34d560", x"5e1f4653930425ee", x"c0d0be0b68f9972d", x"f475d3d06ca4b997", x"e61142167a180aea", x"8917266552aefc04", x"8a8e07be2ac99030");
            when 8674249 => data <= (x"14c5eac11499ece3", x"6ee30e8824d59392", x"e204e90a5918582e", x"baadf5b4a3f1f152", x"fbb9a62d01908176", x"8d49143e952315fb", x"62083f91a61f0262", x"837d82a5860ebf67");
            when 10295564 => data <= (x"4dc08f90a4d480dc", x"c2baa043b40174bf", x"b7b7f592ae722d68", x"f7721debf41ea343", x"e0524a2e7790573e", x"37dca503f59c4c5c", x"704974a3980ff870", x"30f3424c995b57ba");
            when 4275421 => data <= (x"f44b92d282da746d", x"098d078483bbef28", x"8ec8a702632cdee1", x"7fd61b48f8dd93b3", x"f3854417ce8afed4", x"a7ce53607a278511", x"84065ef3806173c1", x"f33d291c12552d1c");
            when 13578504 => data <= (x"13b1a1b22256e36a", x"00d37606a8b278b9", x"40ba848afee6927a", x"8f203fe52b50399f", x"4204933aa25e6d40", x"9d4ef675409809eb", x"3e83391907d7b7a7", x"058a8cf3591fb4df");
            when 12363998 => data <= (x"1ae71d0592ccf691", x"d8544c2b632afb25", x"addd80f4fabb4b37", x"f773f52867d4b74b", x"5875d0606a9de3b4", x"472b29799baa81ae", x"e07f2d656806c665", x"ea819c4ea54940a9");
            when 13454152 => data <= (x"1fe25aa34f26ee98", x"e421fac72faa4bae", x"3f5745a4124e5eb8", x"59b373ee72cd8818", x"bd6bc9960e805368", x"eb69016786562401", x"d60fe47f6f7e9a0c", x"8c29fac3d3fcacae");
            when 24464181 => data <= (x"04f8c877372f609b", x"0fdebe37fcca2e3b", x"8dd46cc3f88f4c42", x"1472371aab91e8cf", x"970268484bd2498d", x"25fb720cbed72e09", x"de4dd0b070af09da", x"024e50ca126c9ffa");
            when 7864958 => data <= (x"0733dae123456419", x"abe15daa21f93e04", x"6eb560078c296159", x"333b2aeffe8a0561", x"b884fff17933282d", x"9cebeec82300a409", x"567ca9be1654f562", x"ecabc51908774ffa");
            when 2672730 => data <= (x"727dae525ac94502", x"9471601de3a0b020", x"e0cc99f4e48e04e2", x"e437115b5d1289b8", x"d4fc4074232b7d92", x"7657eb46ddd1d36d", x"b798a31454a8d8f8", x"ba254d271491c373");
            when 25479127 => data <= (x"bb98043d9fd6f6fd", x"c199e77bce5d07e1", x"fbb84f0f29a66d95", x"24ec6d12e4f31442", x"f502ac98c78bf4df", x"d710a1434d47e746", x"aabc64b642cf0a01", x"9f0875c9ea75a83f");
            when 9782752 => data <= (x"6014e5f3ba22bb90", x"31ff3e5df3d10540", x"765ad460ee4a3948", x"2dab1bc3836cac21", x"b1b6c1095b63ca94", x"e6273f58083fda1d", x"848d12a9d2afd325", x"b2d5ede4f2f9308e");
            when 23204086 => data <= (x"b48f49ca4b492d32", x"ffe9dbff6f72ab75", x"4e3a58f9fc09e0be", x"4b63fae0cf4537bd", x"0ce875a16dbc2ab2", x"08e1ab7ce606cafd", x"7ec88c39c6b18e64", x"e6a4be5ce6550ba8");
            when 9613941 => data <= (x"a32d96cc3b5fed92", x"129f1784db4c01d3", x"a2117ae8e6373509", x"08c6e28c682b65aa", x"add03cc21c611256", x"592984152a380cb2", x"d181556955e28c92", x"3f91c57d2d27c2a3");
            when 28747109 => data <= (x"1d999837c546c8c2", x"50b24423332e0a1d", x"af17879037b5928f", x"065e0ce558cb0922", x"861c20b395ff3523", x"e80da6a086c82dea", x"560e2e95c53913b1", x"f1d2a39f8c1d9045");
            when 3993526 => data <= (x"e08c7a857803b218", x"9385793a8eadd269", x"32a8fe8fac7f4e5c", x"66e2f02e2d317ef2", x"e1f9b29cab8d5702", x"aef60f406c0b7f12", x"844f9adabe61b216", x"d05d931df9781a5e");
            when 28885750 => data <= (x"38149f4a0f748f0d", x"0106c683672d83c6", x"91909c3922b40d15", x"538887adf243b057", x"ca43db3d35b1ccc0", x"ae8f4f3188ce9b0e", x"90d90e5c22d14b37", x"1c37e59c41310c47");
            when 33519354 => data <= (x"9d8b8abfd941f803", x"c27b6f6f10f8b0e9", x"02a565edd0adbc9e", x"9bfdd606d0670dc4", x"3d3da4f004ed690f", x"c3bdddb5c587e9c2", x"09691ff2436ec44b", x"9b8a7101736cc97c");
            when 3395899 => data <= (x"ab192006dc6976cd", x"42087932f7327681", x"353ac958bbf7a764", x"5ee0ff53a972e2fb", x"585d14546013db55", x"386db8e160319844", x"c7d28d8f22806859", x"bcd5b3342c8c36f8");
            when 19883554 => data <= (x"0f6baf55c994cb1b", x"69e46201f99a3ecf", x"c62789ac67137a1f", x"04ccc04d2e5f2883", x"c00e0489aec77a3a", x"2ba51a6c24e2b8bc", x"e597a442d28112dd", x"b4d72ec69657aad1");
            when 1222045 => data <= (x"819db6782721cadf", x"6a7d1a8f45e4550b", x"5650f2c123c7a0e3", x"14319275f8349dd5", x"8098bc8e6021334f", x"86bc32bddb06ab8d", x"6ca221172e312580", x"cc5ed5fc1bc830a4");
            when 29537776 => data <= (x"0dc7603f4304f167", x"f9b52da04bf99f26", x"7f69c1c83e4476a9", x"da6dba05307d7dfb", x"41595c6da40425cb", x"9cdbe7f37bdb630c", x"73325557658f0d44", x"fa6053063f6a5d4c");
            when 11966199 => data <= (x"ecacd6c175a35fe9", x"176126fa2a1718b5", x"eca924352d1c7193", x"a08f48bab17f18e3", x"1f04e6d14eee0627", x"cc7b7174e4a0950e", x"613ff57a2f02e19e", x"8fa824cd4f94e69f");
            when 15967919 => data <= (x"d37f74398ec602a9", x"449da109ac3a9d49", x"c2f5355f71d76606", x"4d6c786a1fea22c3", x"de35e62573cedbe1", x"1a12c20b9019636d", x"1eb16b37bec21e04", x"c93ffe8eb0798037");
            when 1633487 => data <= (x"449b580c891bfaf7", x"4c6a3555272f9007", x"c23a47a443a0f680", x"27f6f4c79ac43294", x"18cd2dbee9db3c29", x"9edb5f685b2af990", x"8fbb09b291c832d1", x"6dfd78e49297df39");
            when 32775266 => data <= (x"6245a53b7e0d7631", x"89e5c79bce844e13", x"f6fd84c250a366c6", x"e67ca53e397b17cb", x"a729791dad8c97d6", x"a8081feb1babe516", x"6c427fbe4e5db7b6", x"5fa006abd61b1cff");
            when 23397280 => data <= (x"5c4c589252841047", x"b4688b4fb90a9707", x"3d85edd4291830c7", x"376789db848aa02b", x"4349e5012b49d8ed", x"eae0af5cdd5bd64c", x"1b75e21fce8accac", x"03a7fd67310b1778");
            when 17268562 => data <= (x"715274a23f0dc4ed", x"4b38e4688767d8c8", x"28125a2d5da4a1ac", x"e709653f759c5932", x"3fe4fc2f77766fb0", x"a29fe94dd318c278", x"a7e6f539d30c55eb", x"d264424c3517b120");
            when 7853700 => data <= (x"a39249163e481519", x"7b5fbdfebbbf2fa5", x"67fa1a2889a12c9e", x"0c440fd4b7a04e2c", x"8ce6cb29753a9940", x"4ed7443cd17ff83d", x"728011a0becaa697", x"93558654f17f95cb");
            when 17230286 => data <= (x"a1e4edc48ec0dbcb", x"8d9694de126f727b", x"3ca9c10559925fe2", x"62e188f2b6609154", x"4b1546e8e99a3345", x"8e7dcc72b18117f8", x"aedd1933ce3a4c4f", x"ef212acb46250752");
            when 24691370 => data <= (x"b6f63cc9c5e9ff47", x"086dcbec18414955", x"ff89fccaa49f532a", x"9437fcdd7e9aa8a0", x"6e03d49a4c26621a", x"d28960f8b07eec5e", x"d36cc95936c88a9f", x"4b47438f85c8cd99");
            when 22950414 => data <= (x"f2a10009513a5917", x"030272baaf6f2464", x"0b090aa577c2a14a", x"372138cda8736530", x"a74e2d335b89e6fd", x"a4b0e65038cb2a27", x"00af95f85a1b805c", x"ae1cc4c5b0805605");
            when 8410562 => data <= (x"0c5add4bc9c8f017", x"838fdbe1309a2408", x"9be36e76219849b6", x"62f53f75103eea78", x"89ffac3371e14249", x"86d58bc05ce8ec46", x"79eedcdaf5653ecf", x"6e8a258854176f26");
            when 4529512 => data <= (x"86dc2185f66ce067", x"a21008a5354072cf", x"d876bc2ce6b383d2", x"205ff88af9bef5fc", x"90bed0258c577f69", x"413efc50a9c893a2", x"ef0e8d0d9211ab95", x"12b2c00bad6704f4");
            when 20888058 => data <= (x"43fc24c16f840b68", x"ca245db039a12b59", x"608c35a6e81a5ba6", x"20fec8d7fb67e1b9", x"4861657feba66e20", x"d32462a26a9c2d92", x"6d007de273dbf1f1", x"7f2744818bb5edef");
            when 19379866 => data <= (x"9e9773620c898b31", x"b0094b2f81466a2a", x"6f480208c62d8dee", x"04900f6165978671", x"50792a6e4cefbaf0", x"7c8f4d979c681849", x"9b72135677eb46ec", x"76c10e935e33b1fb");
            when 23655487 => data <= (x"bbeded99e9a3139a", x"294b2a05b12440d5", x"e2aee5b2b7aa36ef", x"8bbcaf16a02c616f", x"64f5f8f115980906", x"9e8c43a309d15ca6", x"54bf284af60c337b", x"7f0dfd4af569d46d");
            when 17252314 => data <= (x"1d0496bc5ff9567a", x"ba2cd5a69a6d8fed", x"06e2e05636f65b3b", x"dff954e03c08709a", x"027e6172900f06b4", x"7acf9339a55291ba", x"609bfbdf4c19d2aa", x"e4d7265e09f99b04");
            when 28059009 => data <= (x"6459e75f4cadf0ec", x"88e34a5ab7f8df05", x"c2b3819154da077f", x"a5ce199ccf9eae04", x"0f5cd8d1e8f1ddc6", x"e01e27650229e163", x"3e68c11a80389c5e", x"455ba523fd2c218d");
            when 13217587 => data <= (x"001e14b128f0e234", x"6cd2acafa249e205", x"ed9dce33cd93c577", x"4b988c5362c821f2", x"8e5c4daa03fcb8cd", x"dc03ff4daa21ac8b", x"7690d79616a1510e", x"0d40b07f44a5ab7f");
            when 30419269 => data <= (x"b80c4c45e5d1ce4f", x"75fc3146c092b916", x"a00bf10da56fc6b9", x"32a667a94294256b", x"660c35e958ea302b", x"480a7c7212f711df", x"aedbfde63368402c", x"834c81031b4ff173");
            when 24842747 => data <= (x"cbc6ec09a2bcb3b3", x"1a103de6c12b7f28", x"e3bf040421bf3aac", x"b5904b69e731c7eb", x"098220e0c8fe8c43", x"4630f45cd128cfe4", x"6b88910dc309e03a", x"de16f80fdc6d17c4");
            when 27523719 => data <= (x"324c2516d9a4cd14", x"eaa0a4ef59262994", x"dd9283f4e82bed38", x"1c659472519d2e08", x"3f2ece8f197037dd", x"a7a3f21497a3cf7a", x"5fc84bf73e71142c", x"64dd24407652b2af");
            when 23280922 => data <= (x"718b7c34dcf3dd8e", x"2925ca6c1f425281", x"afef3c3b037c6017", x"4a62343d6ba2582c", x"a131d2b62e1c55fd", x"d529aed4534727be", x"de74c1d0754006e7", x"4ced18b8aeacb35f");
            when 22820378 => data <= (x"fd9a5a83aa5bc6b1", x"e206b44a3f7c1380", x"b4e5dc2b50d95ebf", x"a09140b6bbf2a664", x"ed89cae17344c38e", x"fb1641ab4576e8ce", x"4a1a108930625b4a", x"bd5114808b21b8e0");
            when 9062287 => data <= (x"9ca17e6577eb0155", x"605a4c45ae52d127", x"88e04ef90d238384", x"f48a33081f9d3156", x"efd5a2ed6a0fd3c4", x"60ba6eb2519634a7", x"a6a0d33e2ba73dc6", x"3ae19262a792bef9");
            when 12430300 => data <= (x"1b6191cdb71c20f2", x"05ba9b79b157eebb", x"18f0854f498cb530", x"e04548fba6ad9117", x"76f1a4355d788cb2", x"20fd93d9d3771ae4", x"1febea918a40d2b3", x"4f39422d37f69a4d");
            when 13142841 => data <= (x"bf761a8d792d63cb", x"cae429f33f5f4345", x"d8bf28edbf350d71", x"9ff69008491b08c6", x"b019740f94cde2b1", x"22a6add732386608", x"c8a6b7573836b6a2", x"dca8af5b6113c0c9");
            when 10640258 => data <= (x"717d44ce45e9dc0f", x"e77fb391153f80b8", x"3c43a38c29d7511d", x"7e2118fb2da4a1ab", x"d5c1986ef0553143", x"083ed813d9da4aa5", x"bfc7b97ef87a2b7d", x"018a7271d5b07078");
            when 5641146 => data <= (x"bdf6d54b31559dcf", x"7c628d5ba1e76d62", x"b888cc7b54f0ffc1", x"d950db499632cdf5", x"4cba25e436c9474d", x"b2535d4fa1af3693", x"b89142e4751d4160", x"ae17640333b8421f");
            when 15642370 => data <= (x"4694735a637dde98", x"48e690944de51897", x"2968b603f4d80317", x"22438b5edf9e6d17", x"ae964da5584c459b", x"d27c2cd4b35a2249", x"cc32225ab424bbfd", x"5b195ea006d0efb8");
            when 13898288 => data <= (x"16b43e3d42bb6059", x"2d1e8ced36ac51e8", x"8888e06beb5616d8", x"f7ae231ae4266b42", x"f6d7e18e4be6784f", x"2b074b43970a2043", x"e4122585175b6387", x"00ada3ec9f7971ff");
            when 9011143 => data <= (x"a4eba9672022d246", x"69a09bba3df66062", x"0e674fbfef6a86d8", x"1884ef2985a7f59b", x"1adcddc7f1e6a611", x"0e94dad8f7942f94", x"615ea9733ff8a416", x"ac729648c65cc2fc");
            when 2981244 => data <= (x"cea31136d72204f3", x"701875bd1f9c5318", x"9dcc4b200ede2a17", x"5b910093e22ac1fd", x"e707120d7a186c36", x"49d37168c6c644ea", x"90e79515e6a123fc", x"3fb8287113f6aa18");
            when 14891878 => data <= (x"72c90ad738e87f5a", x"eda9764de9e7c7db", x"a1e224eb557edd35", x"dc38aa208a84bf77", x"bcdcf9f303174878", x"0be2dec5326ebd0d", x"ca11a2b4459ea9d6", x"65710fbee258f1a9");
            when 29466200 => data <= (x"6ff1a719519a97c0", x"445c33e85e8bce3f", x"ddd8be929d8f639b", x"24973060b10051b9", x"1aad193b3c3667ef", x"b430aba5a010dc3c", x"526704a675c8b2f6", x"afdb0aece9bfd4b2");
            when 27899852 => data <= (x"bf9de56b6425dc4e", x"ef3ff731e93cd1ad", x"c0292e0f1e2b10fb", x"1c9d8cdbe1cba44c", x"15f658df6189cd74", x"4d4a142c09a0c6c2", x"6d2ee80e9d0e6680", x"d4a78a685e287f42");
            when 18895052 => data <= (x"9dac41b7a64716df", x"d71b2049d9195653", x"d5b7d8608cbcddd2", x"a8c4f26c5d80c479", x"14045b37f6bd9018", x"4837a8353783d646", x"cf5d7d6a385f7c12", x"c507162be34d9ec1");
            when 31512428 => data <= (x"02a0c6c6d3aaac6d", x"677e6533e044cc94", x"842666534ef07843", x"e84ed38716031ecd", x"0f8908ec8478c073", x"aacdd6d71af0536b", x"28681e9a67a5b4ee", x"267a4b2a09bbc646");
            when 7854106 => data <= (x"2175d902ee25e5c5", x"67e0628adc17ab32", x"476ebb93d8e22e7d", x"687d93cd48ea2d6e", x"b7faedc6ca4d512b", x"9b0390449dbb5177", x"e0c35f98538a30b7", x"4e4dccb6fa2673f2");
            when 22706244 => data <= (x"61d96349af12f566", x"cec1a5bca23cc346", x"f82259a08dee60c0", x"63f695e37b75bddf", x"d3aa1f7559bb5c7b", x"18a7c186e05fca44", x"e775b3c18cad22d9", x"c5a2a99413d43488");
            when 22197112 => data <= (x"71bf6cda198d7851", x"784a6d852dd91248", x"17da97fe83bbeb31", x"fcd24fa7fbe71451", x"238f3344b317b3de", x"054a0df26904ba69", x"be422b79c96c94cc", x"7eead401b9bd9809");
            when 24794508 => data <= (x"067c11d6d25a8e66", x"6b27577fb038fedc", x"c1abcff361675431", x"adb562768ac00ea1", x"343518ae70dedf78", x"a20d786262bc2edf", x"4960ee77663f9ff1", x"0efa9749f8dd3096");
            when 5534928 => data <= (x"bdc09e32c20009f9", x"f5eebfb5d100544e", x"d80b562a3fd2c9f9", x"dbff20865edbff84", x"590d95129aeaab4d", x"3dbb74ad6ba93329", x"25756d852b8419a1", x"ac3717441da408d7");
            when 374069 => data <= (x"266de6ba52d347e4", x"95b559897cf4ad28", x"4006928b03cbb1c0", x"9466f093ff39483c", x"ea7050246d13d482", x"1859027dcbbec4f6", x"3027285a09a3b158", x"e96a44c0cb7efac6");
            when 638537 => data <= (x"b6d4070349f43518", x"b492a38aa91899ca", x"526a19ac783c5665", x"870193cc98153bbe", x"c8d549aa820a98dd", x"26c8cfae7c789f02", x"138f559014149f84", x"a236aec7fd3f12c7");
            when 22669432 => data <= (x"71faae474f2fcee4", x"ca634a7d167ff21f", x"1b69c7015c835ccd", x"f6ec7502e5984cba", x"5d9efe34dcc680de", x"df276b378e752633", x"8307dbe9a2484b8b", x"d05b11af71391c14");
            when 33377726 => data <= (x"2a0b2ce79089fb13", x"00e21a3d5699c784", x"866ca20dabe3119d", x"91e8c3cee34c55d7", x"70b3b678d86588c8", x"942c68faaa28d19b", x"71222e7e9aaded7b", x"3172a928261f7b7f");
            when 8241448 => data <= (x"776b43673d399413", x"a83d850037642126", x"bd128dbb2bf09aee", x"817602423b6565e3", x"6e0a0796edb9ce19", x"1383f54d7deb0cfd", x"14898503b89f9f2b", x"4de5b42fcb63b2b9");
            when 21307237 => data <= (x"dea85c72d70d48b4", x"56e4ee9e7b097473", x"57fba014faa90b94", x"f5d173693a19b2c3", x"874afd0b252c6f2d", x"0b027c7cf4785594", x"a98b99355d0ca6a6", x"56abd12eb19b561b");
            when 13972645 => data <= (x"6ef3cd1b447933da", x"9a276aee7679fe51", x"37e1c32ac2015da5", x"c33595424b75583a", x"38de150fcb0f7f08", x"624d3cd89fc52878", x"88e91efaefe11a89", x"fb37f26aaf5accea");
            when 5882100 => data <= (x"26f3895216bd97f4", x"df8a9aef089c338c", x"06f6c518e94b1f69", x"19d5a01ca2668c5d", x"684e62b3ec6e038b", x"911e9f86b99904d9", x"e2fd6461af655aae", x"884df2c2b7bd142a");
            when 13883390 => data <= (x"d9436a0bc15101ba", x"061cfa04f5e1f4ee", x"7426fef0a81796b5", x"4a04d69bf4115b52", x"82e102dbef9a1744", x"dad683484fbe7c7b", x"19f630ec8288751a", x"132c2c753673cc00");
            when 11439530 => data <= (x"06b6a7c7c30c4d97", x"6f0f12032a91be2a", x"692fd93238ad84ee", x"f15521b1ea3c1c27", x"61ee450e61b0fec7", x"bfc4dbf6095ef04b", x"2c12312b5937ae27", x"fb24d4ce4b39d877");
            when 29029979 => data <= (x"bcc50f9803d6c7c9", x"a2701c86effb8639", x"d8c09dc9dbb50caa", x"175b912dfaa63fcd", x"2fc00a5ac4a260b1", x"f3cdddd9980382a1", x"cc45db90bb3aa99b", x"60ebb67bd14fa07a");
            when 6133174 => data <= (x"4f274c444b0bc4f2", x"71798311c4bd941e", x"bd12cd3ff6bdfbbf", x"34121746134f0955", x"521d787c896346e7", x"f6efdd7a36334096", x"df906c8539571260", x"6f263b8e7b5e30aa");
            when 21677665 => data <= (x"17104bcdf55b9b7c", x"512890ca7cab2036", x"e3dd1f74cc048adf", x"4a269deb6d956138", x"a1bb5fe47b261a7b", x"43643d1e42b6d766", x"7af6f925ff7914ff", x"755b31bef0ac3992");
            when 27658970 => data <= (x"b16f7ba5adc55695", x"e290858d271c6493", x"7b6a392e89f8264d", x"95f78e67cd71b011", x"29e0c1060d295ceb", x"91a5b87e769719ef", x"ac7933390825244a", x"d2b75b00a69be27a");
            when 33199289 => data <= (x"ea0b9fed83aaa37b", x"31fc588480fb2207", x"bde344ae6fed7e68", x"4eba2ab9a4e2018c", x"2ae53a1d76857354", x"bcd5876e9d554cdd", x"51055345b4e41374", x"8c633fdeee8b6e4e");
            when 18231169 => data <= (x"de24dcbaa7793da9", x"688638925e8af539", x"f6dc3f30cf6c4429", x"a193d5eefb3d1e0d", x"6f58affad973ae27", x"c22a2380fde77436", x"87f0c7e18ad5a41f", x"dc628fe5ad8e4f03");
            when 26878392 => data <= (x"31fa4341a2f520c3", x"ad2c6a30d2e7aa87", x"69d3f6f833d6f4ca", x"0335f94e77dfb0f0", x"de174d3abb2f7dce", x"288957f6d6f96603", x"49bb55b5f74bcd96", x"ac07f58b82b21ebd");
            when 18621136 => data <= (x"c3af9049b46ed54c", x"aed78fff027dee9a", x"c4c7e650a49b025a", x"b876c4b68f639b64", x"8adcc5d9cfa3adfa", x"ff4d003319dedd11", x"a71ba66bbaf5ac13", x"c3e1844c57a1568e");
            when 27771441 => data <= (x"8a9a1ad1d50e0d34", x"1850130bc3d332e9", x"01219418344663fc", x"9df8302ee5082b89", x"d8fe3c3282f985ce", x"25f77066eaeb4ce5", x"9f0dfe57824f6124", x"056860072ae05774");
            when 11709321 => data <= (x"2e01c9de9ac0eb2a", x"5519b816d268f42b", x"56655e0739944015", x"c13ebb63057554ef", x"93508a458972d0e8", x"3b09cb53d2c3fbc0", x"9482b5498e463c87", x"965029f76faf98f1");
            when 9427124 => data <= (x"216756db43352299", x"4b68bd9f838e6c35", x"9c5408558cc79026", x"c93950283e047607", x"9445bfc320179351", x"9fad38ae46d10104", x"79b37b64e2d35e94", x"d5fec90a59081cbe");
            when 16572560 => data <= (x"885a8090a6274b89", x"08fe812909e2edc0", x"7329d81b62982f82", x"416fa1ceb554a8e9", x"731ef7bc44ee8508", x"a7bf442548ec5e00", x"2ab17f0f150c663d", x"e26040e0261ca786");
            when 22898284 => data <= (x"6541b53f67be45aa", x"b8d90384735abfe5", x"5db26f9691a2862d", x"a4de62cd8438b7b0", x"55bcd057b244beaf", x"d05cc4ccce28a93a", x"270b514eca147a33", x"a89b527f2cbbebe3");
            when 13086405 => data <= (x"43cb2a18bca2e81f", x"5c7d887207b06de0", x"1d7274ae74f2ba4c", x"e9227d66f02a4b8f", x"e47fafd4ea932019", x"89be179214584aa1", x"c404f20adf2a1886", x"660d650fdda59bbc");
            when 23128013 => data <= (x"30fa569b33c6ec58", x"8ff6638fe9e90254", x"0cac994d4ede7473", x"5a5449e546772f1e", x"645f527bcb1b49f3", x"1a9e8b2c7f6edaf6", x"61d4e14d000872f9", x"0702c796b7f3dd07");
            when 4891526 => data <= (x"f5645f2a979b681e", x"cc0212789ed0737c", x"42c412ed4332c320", x"eed6ab3df3ae988b", x"ea3471e81b40bff2", x"7d2d8ebbfff7e307", x"bb17c1bc90732602", x"e412efd9a665fc98");
            when 11218678 => data <= (x"3c8ff195e1d83bc8", x"ac19b9cb47f52e58", x"fd882a36203797d9", x"ebec199c66d0072e", x"076c94716f90a73a", x"04b171d6989a5db6", x"01caa3db1d234b83", x"0bc3ffbdb076ad3f");
            when 16924841 => data <= (x"f9d150c307f22b5f", x"fc3bcafec95a229d", x"0999f1bff1c2d4e0", x"c50eac58b5f580c1", x"4aff819398c1d9db", x"ea31e14a4819d4ee", x"a7622b78ff747d3b", x"a065391af35d9c6d");
            when 29550809 => data <= (x"5fcfb5bfce052a38", x"7aa733fec414c034", x"c288653ad7089514", x"4e99a697739ba4d2", x"6a0d2097e83809fe", x"aabed0d7e2ed887c", x"e9f93c2ed9114ba4", x"834e6736da60bb1e");
            when 32953384 => data <= (x"1aad910821f34e78", x"a55a6d34efe976c3", x"b8186ff13f71468d", x"5d312be4f980424c", x"b4017be02b72d964", x"43dc4e93ecffe8a8", x"4c8920083be60aef", x"569645fde0d4eff0");
            when 1333289 => data <= (x"1cdaa8279e1adb00", x"e87c0207d20b159a", x"6ec4a219b9404879", x"953c0ab149e743aa", x"21d584412b1fbce9", x"0e68e3d72e870990", x"f81a203a5d35e2f7", x"6170dea7104789bb");
            when 13916390 => data <= (x"a2e799d3d7b0b22c", x"a885c375084a982a", x"d86e505a63d0fc4d", x"78389513bdec8f42", x"118e68a3e8c00516", x"61e05cfadd3966e5", x"8167c2568c52db3b", x"a83f5efade840812");
            when 2587347 => data <= (x"d27cacd3870f7a5d", x"e406b0ed90891747", x"b03e1e958b1b5d0f", x"cc6fc64213e2eca1", x"3fe8797a03dd1e7b", x"c390655fdecdd712", x"ca784d818285f52d", x"72227387b9d7e9eb");
            when 7617377 => data <= (x"835a35b81a7b7722", x"defbaaf253433ff9", x"6218192a4018eece", x"acf41f90125005c4", x"9321205209a20660", x"19c92867a6f4510d", x"294b4da8ff42e1a0", x"165c45ceb309c823");
            when 18926346 => data <= (x"a194ca738a3123eb", x"c2dd679badb96e76", x"3e5e100c309fe80f", x"e97c8a73880f2870", x"7d3cf9f51d87e817", x"7f05f273510be1c0", x"472679426b4a6764", x"e44af83cd726bb73");
            when 5897730 => data <= (x"99e636b0b3a22baf", x"97c47a26e0a0b298", x"8cb7453167dc10ef", x"9aecc78cb10475fc", x"15ceb4d5ac3bd367", x"0bf372abe9a52f1a", x"39cdd009f50e1f9e", x"77bd95304c9ac1ae");
            when 32595282 => data <= (x"42fc285fc072d802", x"9119af069230f2ff", x"f0de2e78737c821c", x"4ca1d1883b6681e7", x"c176f7235314ce92", x"545406468042e8eb", x"9ccdf624d4642b24", x"375f86c0ddc22e39");
            when 27321686 => data <= (x"bd6736f65127d766", x"e6f477103a048d90", x"3a1228fafe58c7df", x"9b723c90afa5df80", x"8c730ddaacf5c897", x"823428dc0ffe6742", x"ff6fc286f6de8824", x"933f8bebb50f9ac0");
            when 7523777 => data <= (x"3564a4e46c54e224", x"a2c600cebf7a0e61", x"c6fa3ec5b54f81ee", x"ecd9889ad96dca3d", x"5898d85048bc0a79", x"d8243852d8d235ac", x"62d11e39da22533c", x"a8c87c89067bdb64");
            when 5779936 => data <= (x"9f39eb17d45729b2", x"bd4a2fe65e73876d", x"bdbdd4ea25b4ea49", x"56ab488b4f2ed29d", x"4c541243e3b32259", x"f359c46bcd7b336e", x"4d0c9c11a976f961", x"631990277fd8ff65");
            when 17387354 => data <= (x"061a588c40d2c3ce", x"6075001d5f2de6d6", x"3864f47de82af7b5", x"6ffd2919ff5ab966", x"e338b2df054c4f85", x"489e372fed1ccfc2", x"234153de224384b5", x"883093325c5d55e6");
            when 5137710 => data <= (x"85ae17c6fd7704a9", x"0bbbf26bcf9c2694", x"3c9b1bce0350c488", x"844867d556923985", x"d183c4e48146e69f", x"5a785b013c3ed169", x"245f331823b492f1", x"4210901cce6c2f6a");
            when 19452076 => data <= (x"94b017ae896d91ea", x"f505cd0fa9e7df3f", x"9965cb5b8a4c67e0", x"8ec1395ec4996cb6", x"8c2cd88a7d696bdf", x"8be11bb03699c582", x"5cd8f93173918ab5", x"3c38c50758937a77");
            when 1491744 => data <= (x"144f6a8ef4385a40", x"3f64d13a5e465d97", x"bdcb1b30b0fbb65a", x"1f982f6cb7156073", x"7cf6a6c2481934fd", x"9b872fc0e260fda5", x"ee7d50bffbdb68b5", x"0c5654eb8c5b14b2");
            when 10653660 => data <= (x"76bff9ff1028dc6c", x"77fe36810be1bcf7", x"b76fd5527077a74a", x"f130f6ff146c0402", x"716f5908b85ed630", x"1004f898b2581bc8", x"a8b97e8faa9994a5", x"fc6f70ce75c1e3f6");
            when 21884327 => data <= (x"4ab672c2f647cfb1", x"58010a9b6e7437cf", x"7acf0b2e2d249596", x"a2b53b7f6f4988be", x"eeb6d38920d10c69", x"fa3bc0b787cd6452", x"1630876579bcdbad", x"0291852f56264910");
            when 1449892 => data <= (x"9d4a0c8d484f33dc", x"c7d08f87b6a82016", x"1ce93778d9c20452", x"3fa951e07011df57", x"b28eed6ecc6c8b63", x"40c07f4c72054566", x"e26a9a03c078db92", x"ecb650cc69e41d49");
            when 11740182 => data <= (x"3717ca38cf3a10de", x"c4604fbed5c8d4c7", x"68e59bdcfd5991e5", x"3f62b486c1368b0f", x"f32b5e26b48e2edd", x"b9d34d5b3eacbd4b", x"401578381ea4ba5c", x"e5138084d28b6d51");
            when 29902886 => data <= (x"9a62f4a046e3c2f9", x"8bad2dd090b24302", x"420df651703a4479", x"e183f7bb9b147130", x"24568acff7fdfdbb", x"885067d10a9275c5", x"89c46a5fc33c4baf", x"9d099c5199780072");
            when 29724810 => data <= (x"5005f64f47508bfb", x"8b57af62c8198555", x"ae841b873d752829", x"e42754afc2c8b352", x"e02c72be09e5a8f0", x"42f54025b57f8aad", x"35b39c30d8b1e57e", x"fff7af16e3977396");
            when 33384839 => data <= (x"6d69ff3a62d11c53", x"4e56e652219667dd", x"c1fbf49a98c28b8e", x"005a2be70f7114ad", x"b49a9bcbed898fe3", x"1224be8a4fc3d3a7", x"ea89f5f37090cad4", x"fd335bfc92c009a5");
            when 13275633 => data <= (x"a8082e9bf7f04eea", x"4ce0a865d3567e08", x"e835904a6f2c6398", x"59f9dd428b60b832", x"c512c34692a78cdc", x"d5313f08177206d3", x"7797b57b8533074d", x"393b839f86d6b843");
            when 17177779 => data <= (x"76a1e86c5937fb95", x"512d4d0fb78ce0e8", x"ddb698b60fc18ab2", x"8b8be552141fa2bc", x"90712e0b4bb41fa2", x"79adef0913c43e1f", x"6c641bca1384b53b", x"0bfd762633859a7f");
            when 4006418 => data <= (x"67636e53f5d39950", x"b2f6b513fa3e00f7", x"4bd2f3f09fc6c089", x"3a9316d30860956a", x"41f4c4e7159c0e54", x"e5e1fdfcbd5d4814", x"8c8bb4c52d332948", x"a3a04b8d2d546ee5");
            when 33535002 => data <= (x"1a1679137dd8a5f2", x"8b28ce2eb4cf1502", x"5950fc3a5af652bc", x"a6adf1f58293c9ee", x"9568c43ddc2af2b4", x"dd64a0d5e133cffd", x"b21a9a1f7519b3bb", x"595e1f70111d0e39");
            when 14599332 => data <= (x"5334c9640f4aca17", x"a4cb07ca7cc78a1a", x"691bd704cf5839c6", x"e7e83cc66b7825e3", x"9ec30b73b2c5e9c3", x"ffac5307d45489cc", x"d1bb8a8e1d6d4358", x"dbfd081f5b2477e1");
            when 1923146 => data <= (x"a08727885da8882a", x"868d8cbb1df221ce", x"6c257ac5ba0b36b2", x"3b593684fbb808af", x"13a477417500e1b3", x"ef8a3d47acb1b62e", x"9e2bede095168280", x"50044efd4c5093ba");
            when 9165355 => data <= (x"1191dbcb85530315", x"f504c79fa8c4c565", x"e0d4cc384eaff7c6", x"d3acfbcb5d2caaa9", x"c58258d209140dc6", x"e46d098b5a51e755", x"16dabbb8125f8f1f", x"6e11cff51bb6067b");
            when 27753472 => data <= (x"b754d0440a62d759", x"7df32b056cc784fc", x"ee3b632e779e4501", x"77d1e8d9386d922a", x"51e3a5817c3e2c2e", x"5454df34edb43a1e", x"6eed6425379c492e", x"6511e540acef357f");
            when 5393403 => data <= (x"12f0385a66acbc7c", x"ab37545083517140", x"f9e88d427c3a3b7e", x"04cf09d5ce547734", x"b16e6e320b06842c", x"0641de80597c1fea", x"4174d9404fec78e1", x"31a7c13892655a30");
            when 11837957 => data <= (x"467f7f495c479faa", x"0715b5cf28eb045a", x"742639057fece305", x"e49d6389fb396183", x"27d3f159edd076e1", x"6eebfacac4f791ae", x"4371b271cee0f069", x"1cd4fc377f97674b");
            when 5336240 => data <= (x"e1acf49cf2a5bf90", x"60483478be37a748", x"7d464607deb1fa27", x"f3ad3ab289b75b0c", x"afd2cdf18e4c2c1b", x"c3ad1b18aca08720", x"45b3ad49b395edba", x"4aa817b09d14e576");
            when 18935143 => data <= (x"cebad4e3994ad5de", x"d15437b8cd60e509", x"df186621d0cb1494", x"3684ef5da0d83103", x"fad1675bbdc6e7eb", x"d2ef07d87f897812", x"f78963b33b39358e", x"8914abe16bbb1798");
            when 9497964 => data <= (x"bb72dcb37f6dd88b", x"7b3fa5ca01deebd0", x"debbd7b6ef551fd0", x"393f161abdac2f67", x"3669494a68f91475", x"5699fb4408cdc5f1", x"bd4074b2719d4edd", x"b349cf5076b85a6f");
            when 9998109 => data <= (x"816d34e8db2c9e47", x"c19fe6a8dcf5073f", x"c092ac42e9e2ddc0", x"96feb893ea46f57e", x"48ce0617bcd8c881", x"ddcfe244fa17773f", x"e3bc39d660b88e2e", x"cafdd2beeb71eb99");
            when 27554644 => data <= (x"ef70b8cecc21df24", x"b8f3579441f6b447", x"2cbdc7c890182785", x"8c31f4ed89c57ed4", x"3a35bd3e5eab6f19", x"0cf9e0d47b5b367f", x"cd8cc4edf03cc071", x"d8f4d7bd5a3bf665");
            when 904471 => data <= (x"aa0fe02ff21a89c1", x"685e9afdf2e7ed91", x"a22ec129a1160b8b", x"c1044ef1dcbe85fa", x"f004f499aeb5cf0c", x"03f4c728458163ac", x"4cc400e6a8461ae5", x"19b4f2e095c13216");
            when 20269470 => data <= (x"ca462fdab768bc22", x"e9a1537953ae4692", x"ad5e45b4c5a033bd", x"f575b5f50be14b04", x"505619acac7a54c6", x"fabde7d254d08be0", x"a1eb3d273a0c0bcc", x"1b71eca8b05b921b");
            when 23847645 => data <= (x"57d4fdee2d400f0e", x"629c24b01b7615be", x"ff0186cfcc084db5", x"6f242834ed4fb377", x"d711ada0f4b00ed8", x"bd225394f6d234bb", x"2a669bab30963d9e", x"67a9a1ced2af6b4e");
            when 29630608 => data <= (x"625e1a3657cc2059", x"3b3ebf55ca6d645c", x"31cfd51c6e49f2fa", x"b7888ef1d750cbd2", x"c9ade3de5c7fe102", x"3154569bc470c6b4", x"c601423ca35e9b3e", x"e2147507c873a177");
            when 28118630 => data <= (x"cfaf02bff8cbe8d3", x"f1141f3863efb86d", x"b5721baf772d948e", x"746182d4c6068ae3", x"bf9cc646775308c9", x"dc3e2578dfeb0945", x"51e95943600d7360", x"596dcffb513795ba");
            when 8467556 => data <= (x"8307399bef2b9c3a", x"c0daeac66a2eca54", x"b2ed2f84a3ccec91", x"d0845226310d0d58", x"3382d4835aa10022", x"7c20220667c6118f", x"294bcf1e77388779", x"80dfb6b8c495c85a");
            when 1252903 => data <= (x"b93aba6a65bc7eb7", x"2e6fdbc5b22355e5", x"e6d29080123bc182", x"f6fb1fb15f8fbe2f", x"18cae141526d7af2", x"89ace8da3913133d", x"beea75173a0fe4b6", x"65cc8efdc51f81af");
            when 26710593 => data <= (x"1a1ff8ac54a17514", x"e24a81310c543184", x"e8b979fb30addc2a", x"c0a9494b85554295", x"f7f8ea9c8d710cdf", x"fe4085ada15910ca", x"daacd47fcc59bdca", x"d129c9e79f0d2d3f");
            when 9887251 => data <= (x"565b859bb23e1cb1", x"fbfb61184b36e644", x"18ada885759b5807", x"54f3df5d41fbfe43", x"a96393f387f86e6d", x"d99fd33570657a72", x"19a14e555a840a46", x"fa0704966eacb048");
            when 5886842 => data <= (x"758447fa676c7ddc", x"6e26a92aa73f43f5", x"ba123c9963f1f186", x"1697feaa8c18a062", x"8e1ecb5cced43bc6", x"d3148fd4c292b015", x"67aabff96693427a", x"18c124ceb76c230a");
            when 28723939 => data <= (x"78208fe50f696e2f", x"c2e6f11a15d7e3ff", x"923525c28cf652ad", x"31ac7e258597954a", x"e214ac70013199f1", x"b4d5c2998dd1f1be", x"5d12caf4c83a1583", x"aba70035612e9837");
            when 23400802 => data <= (x"77915cb8b1e9a468", x"344703462299db43", x"5533f70c3b4dd594", x"cf93d81dceb99cde", x"226f8b6bcc40dd3f", x"80355319c428b096", x"0b4ce42e66dc0453", x"8aa6e7a02ab6a2a0");
            when 18259052 => data <= (x"b548e99756b870ff", x"adc5526cbdc0d4aa", x"c9fd4b46369a8af1", x"58dc37c18c693c2d", x"4477272962d5057a", x"1d1c64a7f3a0e501", x"1b4804d39fd75f0b", x"7d3aaf86e9f88538");
            when 4101372 => data <= (x"746d0c35cb7470fb", x"36804fa56ba8a28e", x"56954a4dc9fb8f0f", x"c51a79df24ce54bf", x"22ebc38994afb650", x"a5debeaa28a7e327", x"887737bcccb85c78", x"b680584c200c7524");
            when 19223428 => data <= (x"bf865e300d30103b", x"6ca13594ea329cac", x"56e1e3b86b3e8c9a", x"b24af8f143781734", x"81b9e4218fc03907", x"911f81e8ff76a56a", x"d0192728ee14e0de", x"d1c293b8abee488d");
            when 30754438 => data <= (x"bfdad7c0326d6e7d", x"e51eb07f1cb0eb47", x"21afcd63ae0293f9", x"905673eb4a0b4619", x"d7f6ee6f38c9f4fb", x"6fa77a93311ab3e5", x"58227bc8a616041c", x"20a185e7088e1425");
            when 9706564 => data <= (x"7f5003522af08444", x"3fca968fc7709943", x"14a7f01bde85e414", x"624b0dba23b8d71c", x"ba9842450db50b32", x"98cfb400f0e2e5d5", x"511bae9610c1319f", x"1e91f236833865e1");
            when 13519670 => data <= (x"883db398da8c3531", x"0dfff332228e217f", x"779532ccd74fae4c", x"0cc4de0f1fb941f5", x"e63acd1dbcb4adb2", x"ba62691916184bde", x"2e54c6091c05443d", x"796b3f6b7f5a6a9d");
            when 6596955 => data <= (x"54ef370a8f2429d1", x"a29b250d564355c0", x"301fae47f57e4e75", x"26c69bbb51789b9d", x"9ca65a3a882e6880", x"568b5e7289801c37", x"103c2a91f130b904", x"9437803bbc4dae8d");
            when 27116885 => data <= (x"e94c83639ed566f0", x"3a603c8feb07d79c", x"523994703603ff92", x"aee2d6cfa8c40b9c", x"eadc8f64f38aacc5", x"c4a10547e18661ad", x"40992401be5011ee", x"a789c265265e1e66");
            when 5465695 => data <= (x"c592a416c3a20e96", x"13d57c47ee2e97d9", x"15b56e16ce41b477", x"efc72beb2c988040", x"2b2e7875f47d157e", x"484830030f9a346b", x"4863ec97af142e94", x"b2ba95fb21770fd5");
            when 15925268 => data <= (x"e93d147e8aa251d1", x"282224593b43a005", x"5f6fbd8067b48978", x"ae8f2af1badce454", x"c28b165a427ea145", x"ee69b9782b2b5eff", x"343a3ee0b54e2e8e", x"3f316d46562c4302");
            when 32709754 => data <= (x"3eebad177f6f780a", x"281d853fe7b16140", x"ad43bfb5ae81a35d", x"bb4b166bda0ec9c6", x"0639524af993eabf", x"b7c4c2da38a17734", x"196b92fc4b0bda52", x"e6c174f8f4766e5d");
            when 8076262 => data <= (x"16e042235a6e1ab4", x"f1ff90ac786ca637", x"ad2d2234ebc3b30d", x"ba56385becb8fdc5", x"4315f5126ba1619f", x"c85b12372abb34b6", x"1cc6e32614e71efe", x"be9b038786db53fc");
            when 10536817 => data <= (x"c5e8fbf804005790", x"935acc21ca981b90", x"0cb674198acaa006", x"27a3a9538eba5970", x"e00c2f0073a5099c", x"0d7444998e1be47e", x"ad43c97b1c2666a9", x"74097bf17391f468");
            when 727848 => data <= (x"6aaa9c9be5c54dc7", x"0d814bba80ef7ced", x"f09ac58a151eca51", x"96b70ed8eb5b849d", x"31244081a8e7caa6", x"e5498eef43e988dd", x"a4c7c5da867cca36", x"59597b6aeeea4e9c");
            when 31191246 => data <= (x"43f34b22fc44d914", x"73a6796673d69a5d", x"9094eb529f4af753", x"00105e42dc4244f4", x"c47a1b77935bf514", x"4084e2feca64a9bb", x"f4e46ed916954b80", x"3c37c1560fdb68c0");
            when 25438583 => data <= (x"b9500f4c2c8a35df", x"369e65c212f8ee21", x"eaa084623890154f", x"e1dda384d574ba8b", x"738c9f0b3b67f5d8", x"a7578fda6c6c1eed", x"48b62fededdd7e42", x"da34eef8181ea4f0");
            when 20070485 => data <= (x"9939aa018ffa5383", x"94a46901fcb1f8ab", x"33b54a6462ff3f41", x"09ca25913224db24", x"aabe0babe8b84ea7", x"205652c91beb16b2", x"12ad4bda95345982", x"251aaaf5a3bba7d2");
            when 24775782 => data <= (x"76adeedc0c28efc8", x"519c773247623d04", x"1f67c5732a5a346d", x"6bdfcaa7dfac13c8", x"f42896d92d44d55d", x"b5505b6b1863c00e", x"524bd8975b831461", x"74ef3ef3b87cd5ed");
            when 28174262 => data <= (x"342833b23a3fc844", x"5a808d6bac66fc0c", x"6c30ed01b6178849", x"408332876291b782", x"bd1b57393491fe27", x"191bfbe276b450ce", x"e58efbf619fbef5d", x"26646f5b4cee0786");
            when 22990892 => data <= (x"157aaf0142666aa2", x"514f3f42166025fa", x"004feb1d5e735d3e", x"a03849446981a702", x"ed7f5cdf030218c9", x"160c5a8858e1d03a", x"95ac1713e540d6f3", x"3bafe021c7dd93be");
            when 26762392 => data <= (x"c449403df4496865", x"9cec4be149c82692", x"a39ed74de60a29dc", x"7049258fe162cf53", x"bd4b0cbe3182726b", x"1381690de8bf3958", x"23abe1e7400728eb", x"61ab40c368e48a78");
            when 25827350 => data <= (x"4ad13b8c8d204d45", x"5bb19b5051407ed3", x"369c4963a28c112c", x"09f636e1af33515f", x"74337b1d0ebe9508", x"5f2eaa830615c169", x"f41731ff086b7d4c", x"455b74f427acaf5c");
            when 11186893 => data <= (x"71ac3b4df4ce1a9c", x"aee17dae3837f9d3", x"53889a4172de7f47", x"a74695fc3317032e", x"c0a23a85d11161eb", x"c669e2b23a580d33", x"050f8df8ef72beb9", x"8ee69ec097860bb3");
            when 30074938 => data <= (x"1d6c5ae5ddb9aac5", x"2b6bf34b82b7bc99", x"2085c5f415172491", x"04e4c36d5c70861d", x"9bd3dbe296f0b2df", x"472865146e7fcf4a", x"d3ce445835e733fc", x"db4724b508f5ec46");
            when 23754625 => data <= (x"d0b85909a7465c92", x"6e90694e56977c29", x"eb9b00bba7e1f18f", x"c6266ba882ba276f", x"67e3ce977dc22334", x"995572c4d77d3830", x"43dd0c74e45871ff", x"5394e88e54bf6593");
            when 575896 => data <= (x"ac0202f634c3d632", x"70b93ac136aa4127", x"d24150a70afb4600", x"d8973bc252feef8a", x"e34bae3fa477972a", x"1560021a87660116", x"a447456416c6c821", x"25f6d923389769d7");
            when 6944450 => data <= (x"d0302e4069a3dcb0", x"39eb4c234b466683", x"4ffaa9faafd74e3a", x"e698c4239e7fb0e3", x"b450b13aee11e037", x"3d77ec3166f3c501", x"9e7f75edb330a309", x"4e9ee04942d96967");
            when 10449240 => data <= (x"ba4a351728823f93", x"1942fb12a5c8019c", x"2acacd66b087c927", x"eaea6bd957dab983", x"b200332081c53fb1", x"6b70363ccf69ef63", x"bb63a1522e558b59", x"d4fb19d94bf62044");
            when 4691088 => data <= (x"58934d36a74ace97", x"65c4e398d553eecb", x"ea812e61ca6611b8", x"8e0a7ef0c20b583e", x"478582d7ec1d7797", x"52f9d72b60bc8c7d", x"ef1ca1019e7ed619", x"f3630cc5acd63c1a");
            when 14556729 => data <= (x"cedec500105fed82", x"7949c76792c103ef", x"8e93bb44f3cba19d", x"40adc5fe6d597eaf", x"8009b28249e0797f", x"801024bdf2a1b28d", x"febc84bbe4b6f2fd", x"71d070014727a9c4");
            when 22374955 => data <= (x"4e181475fc67896f", x"6e951181edd51c3c", x"d4fab242dd50d7af", x"ab3fce7306f3da92", x"8741a4692d20505e", x"6cef558b0c42007f", x"189fb54b5c35a828", x"1541fe051ec9266e");
            when 33109025 => data <= (x"ddc7b8b932c175ad", x"40ff361054eb381c", x"ef752155bd8771de", x"5d5225c605fa1ebe", x"f1715375e1399c34", x"e8c18e174aa0261f", x"9c0cea41ad982ef6", x"40251540d5bcd23a");
            when 19113631 => data <= (x"2151ef96aae902c9", x"2d9a336d3af2b3d1", x"63f293850868e5e3", x"756509bacea6d818", x"cfd1de817a6c2944", x"b4d418c6b0aed854", x"05a2bd5fd8a2af10", x"3c3ae073494a27c9");
            when 18232392 => data <= (x"964dda0de74f4d71", x"0729bcf2cba7889d", x"e2b1b440a0033678", x"1cb41d054f6dba70", x"4da560b3e2967ff3", x"5fbe53cfebdf8045", x"f0e08b1385d99db2", x"7efe15556dfeecdb");
            when 12016467 => data <= (x"0820e0333c15b2c7", x"b3f0b8270d57bc01", x"d4d63bb88bb79126", x"b464c1a4f0cf1ed2", x"5f8d3b3b4bd4b030", x"60cedab018a4b105", x"581530d7abf841f5", x"b733cfb2ed5ad05e");
            when 19133932 => data <= (x"5f85443233da9f09", x"6cd2a474f2f3c82a", x"4b88849a61cfba45", x"28639543a53292e0", x"3dd95b5f598fbc96", x"26e8f3b2ed424881", x"48130566da176fac", x"56583d6754be864a");
            when 17976074 => data <= (x"5aa83ff2db629201", x"6f963e457c5d1c91", x"0947ccff55999693", x"3e409c6e3697ce17", x"5d5e15103980b8e9", x"89d4a7a1c000e970", x"f6dfde8f96babc03", x"5a3f92b20bb4cdc4");
            when 6188624 => data <= (x"3fd9afb89a38b99a", x"167e4455a1914da7", x"7066ee5b2f9ad897", x"cf74333e57e2ddc7", x"e53f165ffc3a8803", x"f2ec9e2323f2cebd", x"fb24e9ed4d9e89ff", x"944a2859e71afb11");
            when 11376034 => data <= (x"53f7a39ea4827bb1", x"d07ee0fc3dd671e5", x"81b195c78e4aaf94", x"43dd8d676b7a8cd5", x"bad8e9a1422a495a", x"51b4dc90868c0e75", x"d4fd7c352a368342", x"49d2d4ed48447064");
            when 25179593 => data <= (x"aefcd972d7c8f2a7", x"5298ccdfcae42249", x"b16a640bc872be49", x"ff30d5a6cfc9286d", x"25a1eedbf6f0342e", x"26675daad16017d8", x"15331a357402eaf5", x"8fb6f2e093e28805");
            when 31889653 => data <= (x"5ba00448203a52ce", x"12ae825edd1b02dc", x"9a1a720b813654f1", x"08949239f83d823c", x"80e2712d85d50834", x"11a011edcdaf37ad", x"c1853140cc1be173", x"3b8305bb3e0a4feb");
            when 28054043 => data <= (x"9dbb8ad19c2332df", x"6145dc40127ad1a9", x"174fc3dddff1685c", x"83786bbd051eacfd", x"da9edbcb96c976a1", x"56fb28fbc84a6829", x"50aab3d4972b040e", x"df33b14b06b018cd");
            when 1419600 => data <= (x"6e987b2e0bee59af", x"208c74e438c24f8c", x"58f62a967170bfda", x"61b5589d890d6b32", x"4a15b4cabc1b844f", x"6b02a45700f45e3f", x"8bbc70108cb0d7cb", x"23faf91a404d4337");
            when 2582715 => data <= (x"cde26c0782cb5192", x"a0a24a9abd502902", x"41478ec1c802e383", x"1928370c9b24eb19", x"fc02c4fbc528713c", x"08be9c41435dfd6c", x"d54a2b52d5b7cd9a", x"cc37b9536ad27e50");
            when 13445457 => data <= (x"a146bab4dea34b35", x"8a889928fd1fddd1", x"4e793e1f133a620d", x"d036d7e7c2ab0d84", x"8eb0dee98f9da7aa", x"a7b6a88d6e7ec196", x"1e45558165feab4d", x"0d408400f6c2df3d");
            when 4937708 => data <= (x"4d77e734c93682f4", x"fa4fe4b9306c7539", x"c1dd3f97fde61aa6", x"77d837fd51b7841b", x"71161712c172ce6e", x"678f6613c7828830", x"0b83a55ea76b01c4", x"32ac37bc6306969a");
            when 23745205 => data <= (x"0dfa567f2829d1a2", x"e8ba3346b052bd34", x"7908d0626a87e341", x"4115d800631b3d8f", x"6bdcc279f3431c69", x"c44002f8539f472a", x"534c097f1b7960db", x"d1902a9859e41854");
            when 32722580 => data <= (x"b725857b0e5f6875", x"ee9168c12b869cfb", x"76d86f932de1e6c2", x"a023e06bc6c2baec", x"69475233a69d7c64", x"410558feab871685", x"16b74323e234991d", x"1380752945ade7cb");
            when 11583121 => data <= (x"86af10edd8da4160", x"cdc794e8fe68ffba", x"ab33451364eebed8", x"f73654a3f9fb0951", x"f7bfca1168e0a19f", x"a64f0bb3bf9124b6", x"a0aab82ce068c3f3", x"4be61f5ea6fcb9db");
            when 5876614 => data <= (x"feef1d0c99d8292e", x"4c0c2308989faed4", x"e0bcee716e339a30", x"e948c10f9bf33c21", x"72f756a055053229", x"0b2e7f74995db3c2", x"c1169535f6bbc027", x"b086024f059089df");
            when 28798904 => data <= (x"ae2a59b2897531e9", x"c0611390f59b0675", x"6a94a126d6f83632", x"d6add9de7bfc8c30", x"aa0b1beac7e03301", x"13619b8a909d4ce2", x"9fac2876aaa68e43", x"0cd60a6af6b67694");
            when 5939039 => data <= (x"e4a98e25210b38bf", x"506882a9bc119a71", x"2493551898bf44d1", x"b04141df07a7f849", x"ddfcc2185f435067", x"1a72ad3f2b3244c5", x"e4de94cbf3db33e0", x"e764bdc30c3d46e1");
            when 16726191 => data <= (x"5e70363a01307c97", x"03db89c2c414ad21", x"7f44238cd6209639", x"63258d637eb4777e", x"d9975e9a21accf03", x"81f42b045a36ff91", x"51577bea9bc65f53", x"66adf2cf35d26b8b");
            when 18776975 => data <= (x"86d06e85c11072d9", x"34201487848b51fd", x"c3e5aa69aac0eb31", x"9ecc9b8f8f08b52f", x"b5fdc901e2b8a311", x"3935c39505473506", x"ca511f90e3855b21", x"a08140f3ae1d4a90");
            when 3116251 => data <= (x"1062ffd28735ce46", x"c532f36627dc69d2", x"f6b62c3dd20fbd6a", x"266601f55f9785cb", x"c0a561fe6090fc4a", x"933a24e478056c9b", x"172863324d7fea22", x"910e8e494828a5fc");
            when 31200414 => data <= (x"fbbd0c5f331e209a", x"6abe7dd2d23bf10d", x"273eb6d9c89d949b", x"e649a430c233b905", x"3343f6fe0588b1b2", x"0e0070c760f01f2b", x"ec7c1161fe2ea806", x"c7ea1351f2803c29");
            when 5232039 => data <= (x"3ad904561e119f7c", x"cb1100e4b38adbd5", x"6d1798a806a31922", x"eb453867c4aca1d2", x"d2c95e5365187bcc", x"352ffb3c09f854ca", x"96a9ef3b2871c211", x"600ffb056ac9699d");
            when 25030580 => data <= (x"12ade649790bd7ca", x"dc665b4c254160a9", x"4d8149a19ac80a38", x"5543b7e8ff4ed584", x"37a2bc69576a76e6", x"cefd9fd9afe2478e", x"e5165a1b2a849ba5", x"57180759f1227ffe");
            when 17100781 => data <= (x"0d8d94f11513d8f1", x"75ef16ba1214f055", x"0620a2fe00cdf29f", x"affbc2fd831bf17a", x"060825d5893b8947", x"2d510f35bd590f42", x"acfa8d199db2304f", x"679ba2b1e203a15c");
            when 19597843 => data <= (x"c9645c3375263a3c", x"0eb50e843caefe23", x"1ef371d17369b473", x"1361b116a70da5a8", x"f61beb05621b15f4", x"dca23040bb865cac", x"a3c44b22315c6882", x"fb4ff133d0c4eef6");
            when 18430725 => data <= (x"f0f0574141ef272b", x"5ed835f2674311d6", x"b7bd6e96b1dab556", x"54dad214587cc7e9", x"a3efdd8ff72e51d1", x"402d548508cf0bc7", x"3f69c72c3f757bce", x"05fee974f54c44e0");
            when 20701172 => data <= (x"59fe3689462f3773", x"845b8af669f0e2c9", x"de48981629694e80", x"5bf63141dd8e829c", x"2ce6aa8a3a7628b0", x"fda878c39398411a", x"2dff03f8370ffed4", x"3dd3ba18805b4996");
            when 33822286 => data <= (x"b7170e00107f477f", x"af29fb8d932863f3", x"eb7c1678db923e26", x"30c6e86fc47ace27", x"36752fdb4703787e", x"27d01bcc22bf4ee0", x"edeaac5b58d396e6", x"6496a4a2977ea3f9");
            when 27180998 => data <= (x"8d9413db45783b69", x"c2d5c89bfe47995c", x"f30e45d28d603d32", x"c23ab5c215a59376", x"eb702571a8332b23", x"117007b2545a875d", x"c73f89381ef1a911", x"f5628945d393c94c");
            when 812802 => data <= (x"3d962fd060ff028f", x"2231e89cd95b64e4", x"33cd866bccb91165", x"426d9aa795a0508a", x"331beaf985456c63", x"0663bcbcafdd5d92", x"ae2936d39f6d71f4", x"1b379ce54367124f");
            when 13258176 => data <= (x"03b4822b4532f82b", x"fc83ebc03250e9ab", x"2aa8276199514d3c", x"053da731cb785eee", x"3dc51706db2f6237", x"41dcd933f9b3d226", x"9a4ceceb86644677", x"f09feb33c896c79f");
            when 28659776 => data <= (x"3792daedac4f3542", x"7aa102892eafc0cb", x"facba0b54badd234", x"25d9eb4b68dfc78d", x"8d487dd0f9a66acb", x"6b2a5cc64032fcc7", x"27429dcf23276d7d", x"e1b14cbbcaad8da8");
            when 31130302 => data <= (x"0729b4d41ad255a5", x"b5efda299aff3f11", x"ae995af1d24465b3", x"6f3178640091415b", x"5ce432e852e3f49e", x"8de79942d724ab18", x"27a09f5e96f83318", x"787a00e723c991ca");
            when 31808957 => data <= (x"6b96198797458dd6", x"c64b3a82b4abab71", x"ed4b522add2b3e90", x"a9b88bef8df4a91e", x"1e6fb6f498247b3b", x"838d69d25fd577fd", x"0ef540322e625bc9", x"5f807acdd50cdaac");
            when 23045360 => data <= (x"5775eed05e871d18", x"2c1ee791c2d7c45d", x"bc1bac046bf8bdfa", x"65f2cc00beb5bf46", x"19a2a011dea0598c", x"99ecb48ce4ce7c75", x"39b7b3925a5e5749", x"f87dc3e6c2e491e9");
            when 24397590 => data <= (x"2cdf0f28ed902935", x"87bb72cf6cc2353e", x"1d26c17ede7193e8", x"5c38ff2aa25bb368", x"e305e84199ad6729", x"8291c7f4e69fc65f", x"46d506f9f9e2c3e3", x"9dd42ccb89ba620a");
            when 3822849 => data <= (x"8360681d511be8be", x"df8919114af63067", x"17b5d96c25377ff5", x"1e7fcc2fa2c3692e", x"f5ddbb45ad216090", x"93b206b3502fede7", x"85fd9afea7a20c16", x"68dd07547720c9f1");
            when 328381 => data <= (x"bb9e438920bb0ed9", x"87a572b0049d33a5", x"b1668b42c94f3559", x"6b348025397284a5", x"4df39dd55773d7aa", x"405af59554957233", x"fe46e6cba9b2015a", x"794d3b756cbb53cc");
            when 3193409 => data <= (x"9e768f9f9fa5214e", x"90b7fa2cd91d22b1", x"1ec583ed1c182cf2", x"e0bedbcf679aa8eb", x"296abd193ec80eda", x"89e237f470179907", x"ae40b726fca2b066", x"2487e31ada1c714d");
            when 14154969 => data <= (x"c4b402b1ec475ac2", x"b969ecf2c07fe5dd", x"5c43ba297d916bdc", x"dd31d68c7b995a41", x"d5fd2e4aeef7f12e", x"6470eb2b14b037fb", x"6f1d97e42523dcc6", x"606587ce9474d57b");
            when 28314295 => data <= (x"cc0cde13ca6c2d4f", x"cab3165ba4529ac3", x"945c6ade730d43b4", x"8c3da38ad52181b6", x"424fba1971a37a2e", x"c7a020580323cdfb", x"4074178992847401", x"360bfadfcc4162ad");
            when 26301522 => data <= (x"ce6255664bf827ff", x"ea43094548b865f6", x"793ab222c2664694", x"99b6470f5e2922ea", x"852d1faba196247e", x"9e82b3a37473e0c5", x"93f1f011a192f146", x"be2e1ab0c6ebc60e");
            when 29152979 => data <= (x"716369cd31528f7a", x"74b9b68e4306ff07", x"66c5851159228eb6", x"940ecc0bbb37c9a5", x"2dae4fccada996b9", x"065475d1d203f444", x"d10df5f8828a411e", x"466b5abf0101a170");
            when 24213246 => data <= (x"efa81d7c5bcf7028", x"600a2050af40c54f", x"d616d9ab403340ce", x"0ff05c4f30221d6c", x"472ddb95c8ae5fb0", x"2965f1031207b998", x"866705e603618d23", x"247ac11cbad2f153");
            when 13626984 => data <= (x"2019db582d82703b", x"16dc72403023c0d2", x"3c894eda14164c35", x"7f2e162bbcc86518", x"fc835f69630d6bb8", x"66b489642bbbdf00", x"a70c91b6d5b84b9a", x"f9d2a86139ccec9a");
            when 28103032 => data <= (x"77e4c028420cb01f", x"53f69d92bb8444b7", x"92ec3c5882904c8b", x"57b69c673dec3cdb", x"990d6ae5366b60c9", x"b0afaee62cbff16b", x"4c749de5514f5385", x"665a3529f4f5c03c");
            when 22837480 => data <= (x"e679ceeaf8dbce00", x"cdb09f21e9becd57", x"6347b83329f4ea89", x"e26d266e95f34e8e", x"92553a966b024ff5", x"0ae8a172b36ee58c", x"7770509f599bd8e4", x"25ccf39466246937");
            when 15424559 => data <= (x"31de1a83ebb40db2", x"ff29aff3ef41e85a", x"7365b3fa7335f183", x"257637be00da7d16", x"25b70d3d8a67cfee", x"b733af7a88a06a0d", x"cb57c936b76c39ae", x"40890c0dbf5b66dc");
            when 12382579 => data <= (x"0126e9444d9f03fd", x"0ceafbf9f47b3063", x"e70273b76115f869", x"21a5c9dfd0d9765b", x"376d410ed4678adb", x"d27dab149245c356", x"1cf0e4c5f8f5fadd", x"0295cebe7c9aa1f8");
            when 18735929 => data <= (x"aed7501f605c75d6", x"db7e2224c8cff996", x"cdad931305317d1b", x"422b14686e405290", x"a0bc56c26a958c5a", x"7d2db71c6fff2316", x"80b07d15d61acaf4", x"f7a4b2553ba04b09");
            when 27776769 => data <= (x"beaea4ad06e80818", x"f09b4941c65e528c", x"fed186e2e350107e", x"f7336265f5e4ec84", x"0b90f1f9cb96ffef", x"58edef482b0f34d9", x"6ebbb9d68ee75f73", x"39bf5d018469f0f5");
            when 14513612 => data <= (x"d460d479171e2a36", x"06b2bd308a478fc3", x"9e638c28bbec04f3", x"0cdee26f8b973a5f", x"e06b612bb9ca7d0e", x"00c11ea38e008046", x"4b02413889a3697b", x"63c14d3afc6ff73b");
            when 28520686 => data <= (x"d09ff7ad11474590", x"6a12ab7605cd6c69", x"1f86734200563171", x"29b51e795f3bb655", x"8ddd18da784d5970", x"90de68c18b900742", x"c083e5d3596c850a", x"b0cbafe86740de7a");
            when 25390367 => data <= (x"cba0df41661e6c27", x"323543aa01252680", x"bacd2ee8621ec686", x"9295e53847a58dd3", x"b015e0f9a8bdf55e", x"15acdec4e1d3e52b", x"8208ff464727248f", x"d545cd524e8588c9");
            when 33495920 => data <= (x"c524ce493a6e8c67", x"f77f4b67bfe50e76", x"b2481d505e6def7d", x"a53a17ef0042b855", x"e32edac35d9118b2", x"5d420ea179aa0c97", x"569e5f24d982ecfc", x"671a580481876acf");
            when 29091448 => data <= (x"2ae957f4bf4a5d61", x"804f8b397ff107a9", x"02d1203bcfe7d0e6", x"1741cc27ac9d4c0e", x"13db5695a14e28b4", x"72c5d68a356aad8e", x"b64c3fbb5b3c2c3e", x"e733b6864543fd7b");
            when 23952949 => data <= (x"8230250594a13efe", x"4ed0e7f3aff44653", x"5d7a6ca17e47ea9e", x"3edfa93da2f3034f", x"0dceabcc70feaef2", x"ecc3cc007f02e50f", x"2b8c918b4ad47114", x"85434b371f1b5833");
            when 17462478 => data <= (x"e8bc73e088819cd8", x"77e014d646540a8b", x"3f4554d9407321cd", x"4991321bba7ec03c", x"5cb6441fd61c43df", x"066d3c531858831c", x"f9afada40ea8c869", x"d1d4ae3a3827ea5c");
            when 26492949 => data <= (x"33d147fa203f4e6c", x"cee808be21da51ca", x"a4b4d9401600adb6", x"246b9b563724c8cb", x"6505120a50cfdb14", x"0f721c5b9eae5854", x"2460ee73fab0d636", x"e42e559bd5c587e9");
            when 7277478 => data <= (x"27ca5f9e0a0cc2e6", x"b2bf87f3bb07af72", x"d0a0ccf579c2d5f3", x"37c58a7da7ab929a", x"f8936501a5abd248", x"ac1ee5096d575487", x"3c8a7f527fa42a51", x"6a0b8f1b23b04017");
            when 28711652 => data <= (x"a683ff6dbc0da47c", x"da39f66ae6f492ab", x"94418998371d2542", x"5668c4c5da34d2b8", x"2a747758223364d6", x"f5c5fdfcadde1f7a", x"637d3b85bbae7947", x"f82c9300947d1c0d");
            when 32931103 => data <= (x"f9402bc9230652ab", x"de124f2bd9c10638", x"1cd68771a5d2e784", x"ea2291e13671bf38", x"7822e53108a3412b", x"8f85378da401a8d1", x"d97bd4991a381b8b", x"11fe0ef244a12b7e");
            when 14783936 => data <= (x"0a364a244217948c", x"8230aa806f3ce789", x"1f5272a1a5ce0b6e", x"4cdc3d0951bcf3fa", x"9c60569f29423f8f", x"dd84bf7264aa1660", x"347cfa593a0bb900", x"7beab9279c3de34b");
            when 8033091 => data <= (x"fc0a92be7e8778dc", x"d029ac4aab599564", x"6951518f8e7cbd8b", x"ef94629d35accaea", x"f142cbdf52545c37", x"4a5e3dfe08357403", x"ef78161cffec2dd3", x"b9f42b76a8efe884");
            when 29357259 => data <= (x"6e6c762c8aafd346", x"7de2ee4c6a303a0b", x"b26c9b21045f0835", x"311b603d7bb101bb", x"9be2299e27254031", x"8f3c7dc09724fb5e", x"239f9f9472ea896f", x"4d02b922d41bcdff");
            when 27796390 => data <= (x"fa51f5c0b07ec22f", x"4fb53aa372996b9f", x"05dbbf09519f40c0", x"39a91707614aeb80", x"98c386dc7a1f6775", x"63a80577aed4b341", x"3c0214689f7ef22c", x"d41115524632b382");
            when 31712543 => data <= (x"18565649c439db83", x"18591808ce994c42", x"b546b676d06bd737", x"0c6ab2803a391e78", x"e045bd90afc30d39", x"ce3185a9aac6ce90", x"a7f85dd05bdcb333", x"15aaa275f34da8b9");
            when 30625197 => data <= (x"41a480d188a83a33", x"ef30893d0c8ff78b", x"de5e3ce2e8345cfa", x"637518608b27c9df", x"6fbe3529ceaec3d1", x"6b01386a58f01b13", x"05ea63afda637825", x"f452e8cbe8829820");
            when 6409556 => data <= (x"898bfb7e6b875443", x"091cc3bc425ae7ef", x"5048f8be0649e6d7", x"0e25d0fab77be1a5", x"4786e7e1122ac567", x"6d81d6a9dce1cb04", x"1458980fccd4fa84", x"7be9607ef0335181");
            when 18428091 => data <= (x"b54e8b5a4e2b67ec", x"2477e825d1609d9d", x"8db4a0ba84d9481b", x"08f13329dd9bf7bc", x"2c7c1a80f597e952", x"a2c32147a1726cda", x"d559071e3ffc35a4", x"fc9d9d4bb58115ff");
            when 4913912 => data <= (x"5950f38602b453fc", x"1cf3af50dead172d", x"81dabc14805d0e6c", x"8573731b600a3f6b", x"de2866dca884b97d", x"ac3a120f1fa3048c", x"98444b4f4ee61bf6", x"add01b5b08959f0b");
            when 10339969 => data <= (x"de2fbd10790e9fb1", x"a196818e32a13f34", x"bbd44e749640f46a", x"16779bbc7da78dc7", x"364838fca88f0592", x"8223b6e375ecfefe", x"ef8ce0338d78a2ed", x"b6517c13a9f04153");
            when 25346361 => data <= (x"ad20099e089f3e62", x"6b575dda4249e71b", x"a35c8dbd5499a588", x"5da1a360b0551f20", x"bd36db007d4a9765", x"836938c1b31218ad", x"0d16032a96879cfd", x"bfa3640158a502f1");
            when 30427043 => data <= (x"73dfb1cbbc18fa7a", x"b21b8408da9731be", x"5325e63ecb2da2b6", x"0c200eeadc301163", x"4be4cb3af5f3e304", x"a81a6eef1fe48829", x"cef9dcf09e0d0a1d", x"2a2c463f8765fcba");
            when 24488163 => data <= (x"c1df38455d3833cb", x"1afecb5e25f89258", x"6a6ddae1fb860f3c", x"4b00979aec0cc8f5", x"c16ea27fb75f647f", x"16724fd8edee33fc", x"ef79b3bb820e6163", x"f462170e88c2fa01");
            when 13617498 => data <= (x"e07033403b40227d", x"8dca52aa0928b23a", x"bdb6b5067d2e9c33", x"45508a00dbe88c55", x"b2b0bf9ed12ddc32", x"5fa11e5b33af65ee", x"a78ccbaf19bd0484", x"5a442655b9d52914");
            when 15445582 => data <= (x"5920fcd48f5bd5ba", x"706226fd70893aec", x"fb06cc2a6c546653", x"d0e5719bfcbf74bf", x"b71b81b00afffe88", x"64aee8f5f3604c35", x"cacd2557598e67d4", x"f7a12c6a0314f9c0");
            when 15643445 => data <= (x"0c60ec510331d147", x"0a9b48ec5e308975", x"2298dd2088933b73", x"086a29c841688059", x"f71ca337dbafaef8", x"2c38ff2c42d9d446", x"3334d9d6fc0a3245", x"8affd4e2c4864d19");
            when 11890884 => data <= (x"29f128d953242507", x"657fdbf2230878d6", x"1df6d89169498cd4", x"99c3a8cc568ed7a4", x"0b0fdc0ea7392d8e", x"79459e059b8a71ab", x"c8188b0fda3d09dc", x"ea36b8372d3491b8");
            when 858457 => data <= (x"7ffc71a886566e7a", x"97de5a8d3b63c2fa", x"1f3064397ce490c1", x"de044a63509ea5bb", x"9efef7cca2453d04", x"749dea2640a9a457", x"fd77174f239648f5", x"9afe1c7ed5a02986");
            when 10151062 => data <= (x"ce1bb302737cb6d1", x"bd96b2526022d855", x"6772dc6a561fbd06", x"703b68cb81405c61", x"1509f8d1d78a2200", x"4ff9dde39e5cc18c", x"cdbc6ecab97a776f", x"3e2f61f3df1c6fa0");
            when 17007259 => data <= (x"bb1de3d9763a62e9", x"3cd437b3c93f80c4", x"7a4921b9bf70199a", x"5e37b26d940a37dd", x"6ee648bc4e6b00de", x"8073abfd3855952e", x"72051711a73ac1a6", x"9ad26befab150e84");
            when 582338 => data <= (x"93f13e709564512c", x"1c667f104f1e638c", x"d6343ee1c2dbd4c0", x"5ddd94e6a7353a46", x"02f0917e8a74cd40", x"f43a4eb3f6352438", x"687d782ea5b87724", x"de732afeced10a76");
            when 14380366 => data <= (x"e9bd426548526d1f", x"5889e1b79e40508e", x"bf42edb9198a21bd", x"f20652d1c52c88f1", x"45deef3717b4832c", x"af1cd57c3b085a17", x"2ed4a886fcca3b5a", x"be955a6cec7a52cb");
            when 30464383 => data <= (x"2d216792cee92e93", x"d14c7ab16d153657", x"03f8a7690f89130c", x"5713ce4a6a4309af", x"4ec575caee4923ab", x"889d0e53f92c1ed6", x"2f717775e68cb185", x"39d2b82eb112e705");
            when 19309912 => data <= (x"cf48b69c9fbdbe20", x"c2f05b7298625574", x"53c52d290cb0736d", x"91ee30720bb32fad", x"e4cac518275129e2", x"6462a4b11ea3f53b", x"10253201e917f0c5", x"4857cf2c79e0e966");
            when 16940266 => data <= (x"4781184ce7727b75", x"cda6c26029e07f99", x"c73a18839c19d43a", x"707cb5bbc1c87024", x"38e5adc34388587f", x"02dc01892f3bb085", x"2ddc68e91aa471aa", x"1b88febbb3f7dca3");
            when 22801986 => data <= (x"3c6f426e8c4357ce", x"aadb97b1320480f6", x"df2c87754dc2193a", x"314d80c735c4091f", x"9027f848a38d1842", x"c1929a98bb90f56f", x"c0ea515e903b0ec0", x"189e35fb196a4031");
            when 30464655 => data <= (x"d78d9305b4ebd94a", x"1273231fb503a254", x"8541ab31b2b4cf6a", x"f960b00aba634f3b", x"5db741b26cf3c8d3", x"42aa336cc186ac90", x"60bc8138bd82e03d", x"359bd2c839db7ffa");
            when 26205696 => data <= (x"3b10221b48491e78", x"06a9b3a1635fced0", x"6414169721ba78e2", x"0bf623bf0251b9e0", x"3511e5cd0680bda8", x"8f280488bc4a3c60", x"93409437029061ae", x"0bc1cdbc0401435c");
            when 22874279 => data <= (x"8a575661265e1171", x"79d92727b39906ef", x"06a8d4503040cd67", x"9427ab037ccc25c4", x"7d361f3c578ecaa3", x"4ba88ded2aa97efb", x"9fc7ef4a1118d53d", x"0c688e96495cfe6a");
            when 33790991 => data <= (x"791240aafb34e473", x"9b0778c4786d459a", x"92207f20c2702762", x"a4de8a655f76e1b8", x"67119ab697f9b88f", x"84836a4e2842aba5", x"13099182f6d33e4f", x"ba23595203f290bd");
            when 13946010 => data <= (x"58c9417db855a9ce", x"06c6450e1e89e17f", x"3203f1f167f372af", x"e6586ccfbf32c7ec", x"9bf7e5c163b3d353", x"d12b85000465d10a", x"1d6d2b4b47c4f415", x"98040fef35aab05f");
            when 969754 => data <= (x"e4b983f1d32123bc", x"0d6caf8182201144", x"09ba6bd4c1ff57de", x"6bc0a9ba185fb539", x"83b86bec17216ee9", x"f6dc139f3eb1660a", x"dbeeca1b2b9d0f53", x"6e66bb4d00a20e12");
            when 22847366 => data <= (x"5832e2c4720b37fd", x"2054dd225c86b906", x"f207ec059f16a0b3", x"748257e3c41a7b3b", x"37b40d1855058838", x"d62b69824b2d8633", x"74654e871e3ce405", x"b57745c6a0ec9420");
            when 32355579 => data <= (x"f7492efefe9a4dd1", x"9277feacdacb0afd", x"bba7f7fb9c484889", x"9e68fb46654acc5c", x"396b7f0a272e8b84", x"2bccd33e62a4ddb3", x"40627818f9a6bd84", x"ae4ccf8f49379330");
            when 25844111 => data <= (x"7fcc901bb7830926", x"de9b44dacfaef749", x"4e3f028e01c22c7d", x"4ee1b92803424cd8", x"2512cb82fbc0ea80", x"e1d26126a1515caa", x"2a42ea8dfaff7f09", x"949a01aff9df55f9");
            when 21329948 => data <= (x"d351fe9d222832a9", x"f87fa8d420310b1f", x"817042978b569300", x"e401810a9723f8e9", x"379ed61be534ab3e", x"602d80c902e5c4e9", x"e4b05992459628be", x"bd84ed0a71b40ab2");
            when 23359330 => data <= (x"d0c8574db964561e", x"5b19343c221ed005", x"92d2fcef5c274633", x"f1223250e04beec2", x"976a62c3f36395a9", x"804ef7ffd23878a9", x"c6b447ffffc53eda", x"fc0d4b576c0bb8ee");
            when 2202728 => data <= (x"9f2c105b06d8a2d7", x"d64bce5ff948ac83", x"2715afbc883dd98d", x"ce31418351a09f62", x"8bcbade8cf3968c3", x"135f11ef0dc5ff52", x"e02cc92ba367a03f", x"d7945619dc384658");
            when 2041101 => data <= (x"9b1b7df06a73b907", x"96d5f246b0a208c1", x"725d12dd1d2d3f27", x"732c3b20b2d5246e", x"c2c39db3f63ea689", x"41f1887d87ae7da6", x"dfa103285dce5ecd", x"008d79f282bd1de2");
            when 3068058 => data <= (x"320ea2f8fe1d77b4", x"295d93bae1745c99", x"b828d7b51efe9f3a", x"5acd05d1617f035f", x"2c7d83dec4641d3a", x"8e3060238e009250", x"11e9cd91844cd022", x"095e76e82b84b476");
            when 21885214 => data <= (x"3923fefcef07b864", x"1a24a3945489e11e", x"2a2d41dabe1aab0f", x"cc5c0c09bf967ae2", x"022a0e6d37fa726d", x"b54533f6ae58a60a", x"3a6955498c144318", x"4ae1dd7c9021cd08");
            when 29992929 => data <= (x"0eace051e49aafe1", x"eaf05a11d01f34a8", x"978d071e2a4f68b3", x"8c6020ef349ddecb", x"e10af43f693673c7", x"a059483c4380ceae", x"19d763f7baf0ee9a", x"f9fa7bbacf322a97");
            when 11209007 => data <= (x"f234e7e737801703", x"1bad190ba78d3357", x"851bbde02f643a3a", x"288bea258aa6dd40", x"bf0246a8624b299c", x"53ccf8fa7e3e347c", x"c33611d220187c54", x"12ac031c8e004c76");
            when 7809405 => data <= (x"5ae4c1c00bb3c077", x"068c862d08fa90ae", x"4d61d1bd6e7b0e34", x"a4e59d701c3b6922", x"e6553cd644a1f09c", x"f75ba0c809e49f25", x"5ad96f90212c6285", x"ebf4355244bb4900");
            when 16013652 => data <= (x"2b87e748a9e57da7", x"93d29bc77d8b5ef9", x"07a75f778bb7417d", x"2b8225235202f33a", x"93359a2c7dbb13ca", x"ee71fab5b2deb85e", x"a2cea0620cda2fd6", x"860430385bc4d9f2");
            when 11645231 => data <= (x"bc33ebeff5ff2eaf", x"da8d210d144267bd", x"6bbc354502ac1483", x"b444c0dcc0972cf1", x"2d069d47b46d4e28", x"9f8388ecbc671cfc", x"c6a0ed51e144d8f9", x"82db874f2149c617");
            when 32369610 => data <= (x"88312faa083fa422", x"f16809e6dc79a47e", x"54f440f21ab7edcd", x"851ef50efc5f2eb9", x"07fb9d7cb27082e3", x"250d4c444df97fda", x"f315013bb242794f", x"a730910335392374");
            when 16285352 => data <= (x"ac57a296637682f8", x"d72268a82d98869a", x"9cdf8d404e0c7ee9", x"4ec4725b357e1ea3", x"c4d0c09945a7dfca", x"6a42fec42dc199e6", x"b5b42bd38ab90216", x"d04fb868cbf51598");
            when 18704126 => data <= (x"ba4f71c934be0ad6", x"10b634bb8da2dcc9", x"b1e9f2d92be3a73f", x"1c30a2c55800bcff", x"862be0df1334a41b", x"7d3e729aca638ee1", x"fb4be426be67e4e6", x"31ea0c057da96963");
            when 32760912 => data <= (x"cfc4e0e0b8782def", x"2a4728b0fef00764", x"c21624f23bcebb3e", x"44b6f78562941a89", x"58d245213f8657d8", x"1c91b1e001315707", x"e9385fe49395c613", x"b20ace9812c135bb");
            when 16490747 => data <= (x"1eb3432f77caac7d", x"0252ce90a8d9b52e", x"496d9f2740ac3e19", x"7276d230d6bbdb2e", x"6e083edc24a0ad28", x"7fd66ed73c8d1619", x"c369c4c0ef59db5e", x"ac26ed9d93f49c50");
            when 27875490 => data <= (x"3af78156e1e8ffef", x"77fe35237ab4c935", x"cfd197b3525b52e6", x"6be2b40b921b8384", x"d115918aa6ddaf70", x"1136e66bf15eee18", x"a0b1d2ae0d9d41dd", x"396066da4047886e");
            when 19737764 => data <= (x"6a476bcdb3523c46", x"6a1e962c776b140b", x"0a7165eacc0a742c", x"ae41aad412bf4722", x"be7dc926068953ab", x"3bf89a578b613d3e", x"ce72ab180ad8e053", x"bb9984ee2d7d6caa");
            when 26384309 => data <= (x"e03ac45d07c4ecfb", x"e60bea8fd9fc207a", x"b294b73c52cb71d6", x"d213b6bed3dbfd8c", x"ab5958952acb1397", x"a180e9683bf6d9b6", x"e2b9e950f09ebdb7", x"00a9529da5019bfc");
            when 23592725 => data <= (x"9e6d66eac664333f", x"f35009d57fa14bd7", x"29d4aa460c1840a0", x"9c2d136cf2d0da01", x"7a4649910e714314", x"a004defe9b511fb0", x"c4bff92e19d428e0", x"aff4312fd756a42d");
            when 7119189 => data <= (x"f5c1d7a4d9866533", x"f76bb72228cbd6fa", x"5d126ed5a8936b24", x"97fe4767bdcf86f2", x"62577af9115f9607", x"b575e0cf7af4fad7", x"359251cd3eeff78c", x"863baacfefcaf05e");
            when 5861267 => data <= (x"2dbcdf1ecbbc9caf", x"8807b178d06ea1a2", x"02106145fdf9f09f", x"2897a33beb4407d8", x"2f846ad5af3d7a35", x"02549b422f0ecc4f", x"a6bd803cd7116905", x"3310b5abe8778bb4");
            when 33499629 => data <= (x"9c84e339101c95aa", x"1f71b0e1e01aae50", x"ffe622cceded65c8", x"1f89e6785ad02ec8", x"24515ca5ca1df4a6", x"f1d1733e3cfb9fc3", x"0821e40f5e9bbd56", x"167d0983568020a2");
            when 17373831 => data <= (x"ae8c249a84470b4c", x"69f35739b6f04ca7", x"272d693e489cd690", x"4ae2b9db55ff3fd0", x"c8d73a8748b3f0af", x"59fc4c1b3bc3886b", x"5b2e3ae466540dc5", x"67a2f9a28c6d85e3");
            when 9132421 => data <= (x"27606fa10fe63f8e", x"e2467640fad86849", x"cf5f9a7ff6d8fe0f", x"264137670fe0489f", x"f09b29d7dac2f566", x"637fa75b8f3f9a1e", x"6937578698735a88", x"ea1ddd81af617c64");
            when 21655415 => data <= (x"09820febb7296c87", x"f3ff288da0dceaef", x"a77c48bc10f2da32", x"be897651bb136d5d", x"7fece4b0218cbe4e", x"2567dd72cc43118b", x"2d418a33b4b48de4", x"386b65e8e76dc3a9");
            when 16998149 => data <= (x"04f38cfa3257bb9c", x"fc0a763eb3042227", x"162767b409e6b1f0", x"b1266707571eca3e", x"07fd878689410d81", x"87fb33f92e675346", x"b2ec82d94f7e5084", x"50dbfcec95ab02bc");
            when 2554205 => data <= (x"9416b7510309fafe", x"2ec065bee91e0cad", x"17ea8b620bf4074a", x"1dfeac7b721aaaac", x"8fe2411c89cdfd6b", x"8cbb971d174bf601", x"82b168315fc2d968", x"a30cbaeb246cf920");
            when 7322848 => data <= (x"b341caeb4689964f", x"d2a2a11595ec0c01", x"c0406e3c820f81fa", x"ef46e8fd29ab7d82", x"cf5b4d6f27aa9f6e", x"75052008e719850f", x"af3a32317b44a02d", x"33b1a24fa288bbbc");
            when 9768291 => data <= (x"1b0cd1ae507b1369", x"e964da60a986e4dd", x"cbad2c4cc697fbd5", x"d63f3fd170be0037", x"c7da09359709fd9a", x"35bc2608fec883fc", x"9a45e709eb704d9a", x"dd1d926f35e11538");
            when 8249027 => data <= (x"a24d93a94fba9346", x"1a42bcd2017b0d76", x"cc3f771bda0b0373", x"a394ebce769df97d", x"9969a8a87692da9a", x"af8159b4ffce7d1c", x"2e8a78f3f0477e7b", x"7d7b276bbccdb9b8");
            when 7402006 => data <= (x"b060e07bc8933de1", x"184605c14368e5fe", x"bb723e1bdaa6d9ba", x"2a7569bbebf978fe", x"3359b3976e212104", x"bdee5da61a72abcf", x"d5b589c65f222c02", x"e3eaa7a5bac04fc7");
            when 10928313 => data <= (x"201f949b95f25e39", x"cbc797377c3ecc5c", x"b05760adc7beb3ae", x"03e820e6b8c75804", x"cccd4c9b5075d5c1", x"fcb346e39d4a1a7e", x"96d3eb7eaa756b27", x"d2051467ba54ccb0");
            when 29603995 => data <= (x"817c5186acbccf60", x"ef2c8cf926598f11", x"e221ea06389c7dfe", x"da7f384d37f62084", x"676412dd4024d02e", x"f0b6936f51043def", x"a14e600ffd7697e3", x"f1d7fb3c07b3cfa7");
            when 16734775 => data <= (x"36e00f5d81f398ff", x"e357944a9053e832", x"74a73e1a0da5b652", x"47701624e96ed3a5", x"551d7350f72fcbf9", x"5631a050e50c3b7c", x"2df9e3a089192176", x"6e50b972b41b0847");
            when 4072276 => data <= (x"a07a30b71d143af2", x"7b47a450944289a9", x"54ddd6d7228ae980", x"f5aecc00ed83cea4", x"3012f10b05cd6a51", x"ebba56ed5e1371fb", x"9275203494053cca", x"dd94d9fd17f55213");
            when 29050322 => data <= (x"61ed793a2c7b09f4", x"b8ffaba7eb6565cb", x"6ae4c7390d1e079a", x"a46c59925cc5f809", x"033016ed7f590352", x"09763988317ddafa", x"0cf0d5f84ee9dd97", x"e8f2e7ed677c8074");
            when 11954939 => data <= (x"9fc909fcdd2994c4", x"1cb080da0840c8fe", x"a3d496c7343cb91d", x"ea8f053fcb976fd6", x"226759740fa49f1e", x"10a7e35aa809cdae", x"5184168cf2fdd3dd", x"1965e91d9a33120e");
            when 788058 => data <= (x"b5f9cdd3e980d96c", x"8800f2fd6efd21ac", x"07fb03c8cb0e9f31", x"98ee060b20268cda", x"509512afe86192ff", x"0f26a35b87cb1ab0", x"04817c037b929983", x"8abde5ecd57ae758");
            when 19383688 => data <= (x"d90024daa94174b2", x"76ce5988b288d96f", x"8541a171c660ad7d", x"dba4f69e730fbbc8", x"9485d7fe1ac7c0db", x"e5a048dcda67c8a2", x"d7a9e57c19d0d4af", x"ca7f2e96641ad59f");
            when 28587638 => data <= (x"ec45a3fbbe597544", x"013f1e8e72e8732b", x"e24db13c9d1c2743", x"8a8841b3e76981fb", x"3f029973883c10de", x"ef5199d9787c6f79", x"adc6dca44726a666", x"b865ac8232de1b86");
            when 24491468 => data <= (x"7e26ad6e06fe5c94", x"6202ab00891df249", x"e10bf18e71538deb", x"57451fee7222ff16", x"f480f71a70cc7ec2", x"6ce2b01db9c3b54b", x"82194e6e0b013713", x"950599aeb1efadb1");
            when 8606690 => data <= (x"f8fa4c26e4fe0848", x"e6b147deae964dc4", x"2da5c5bcb65b843a", x"d18f2723a9995785", x"bd0a35b86f344c5f", x"2f32baa256551904", x"d3e26156aa6993a8", x"038569c5fe0f13ac");
            when 13848555 => data <= (x"f732623daac05432", x"20fca23e203119b6", x"a678367bcb905305", x"60f3bea36860e7a4", x"a95738222540ab6a", x"d130258a2d37d1eb", x"0b47c0257ff3b952", x"417d2f2b0adf8582");
            when 23448775 => data <= (x"cb15b52b8240f9c3", x"198f86f6181a58c7", x"c3958388ca2ddf50", x"6b4b1b61b9a71e12", x"d5a0d3b4865517eb", x"4401e0e457c97155", x"6c95568694071b71", x"2dd8a7458e03f16b");
            when 12525873 => data <= (x"61dbbcf42c30c2d4", x"9152153f00cfc356", x"c1e14b8e663abca3", x"0ff8fed731fe1a2e", x"23d2c96f1cf6311b", x"a4c405b932b1ea76", x"ec0208f4fc05293b", x"0fc24f1618cb47d9");
            when 19143704 => data <= (x"87d536f71046101e", x"e5b2310b704e500a", x"a8dd9f659d49fcad", x"da83f854bf15e197", x"a33475ccdd0d22d5", x"f589b885b6c3c096", x"5d8f17f8727ec32c", x"7ba3d8bc46ccb438");
            when 6436368 => data <= (x"7ea1c08daee5c25a", x"8add033a764fdaac", x"071c451c9caea973", x"53f9301f663c69f3", x"7c92c9e19c093318", x"867b1f8fdecf0a4a", x"d1a3532696cb7a8a", x"a095d22353345128");
            when 31388974 => data <= (x"e1c035683642fb19", x"c45651a25b12c120", x"8c910250d0a30570", x"aa670d96342d400a", x"22f216baf21fb958", x"cde27fe3db640f37", x"6ec4570aaa769196", x"33bd37b521448a5a");
            when 5861966 => data <= (x"ecdec9cfae1cfad4", x"9d744e21706c5a93", x"c952c18a030b4537", x"90c52daa58acd740", x"0ba09ffd66a61c5a", x"5e79018790984104", x"ee4b8e0aa4c4d9bc", x"9265d72fafacde17");
            when 9573098 => data <= (x"4af58c0dc11b12f0", x"f1d1ef7113677be1", x"ef9c464cc2c02a58", x"f511d6f4d9de4627", x"7179456716a4600f", x"9a0c6c1ec2eeb627", x"f28fb0e9e851394f", x"360ee5f7bff231df");
            when 1868231 => data <= (x"a4ab56831fd2869a", x"e7250388764f5c18", x"6c9b2b525aa4aca4", x"38b9249510ce98f5", x"7af09a8e667af21a", x"b4d4973ad9cc8c19", x"a6ddc1a7e98ccc8a", x"3cb096c2247862b9");
            when 12711546 => data <= (x"d51e0029f2493eb0", x"8e4158fc6ef1de2e", x"48f48324c9674691", x"f7e68fe7f35fd82b", x"b1a29fcf79f061f3", x"116951a46757eff2", x"2c7f591559e5b81a", x"12d7bca67a87dda7");
            when 8431010 => data <= (x"1095e9121d5dd1da", x"aa1f3ccb3909b901", x"02ce76f497e6afc2", x"a8f1db009a285629", x"af25cc3dfb3998f7", x"52e6cf5a4372640f", x"5012e39a7d374e6b", x"503546d4b503190b");
            when 22632473 => data <= (x"ed57331f31e55422", x"8fd0f8fc81e41c18", x"06a6f9f99b36ac7b", x"7f44dcec7348aa5a", x"0c58d85a5dd9651c", x"854d6c9e4e3d3f1e", x"52aceb8b4ef71c30", x"ec3c9bc89519574d");
            when 6381900 => data <= (x"95711f13485ad583", x"109e71ed504ce77d", x"f253c1b74daf84af", x"32b837e20a5fa5ee", x"7e4a7dc1b17533db", x"bb82eadc504f2714", x"b650c840cada8770", x"170ca5bc233dea53");
            when 17243096 => data <= (x"a825cbb45b5d18e0", x"46c74197e45e7780", x"daa194d9af8ca245", x"74dc45b74dc38076", x"67f2a2c553876476", x"8ddbe2483cdf2d3e", x"9df43b9657a57050", x"7c4d0bce47e3e445");
            when 9499576 => data <= (x"7042bdd22f5c87bf", x"ec57061deab69852", x"84fc4a65ea0cf1b0", x"eaa0375c5a215ca7", x"3857199f7dd21bdd", x"a22bb1eac63b5ec4", x"77139a29a2af03ff", x"6b11d2d0ce10fa70");
            when 5524344 => data <= (x"bfac8ef0b9580b20", x"dbe372c7439f5ccc", x"1b2dd0f30c7b20ed", x"2551ae6071ccec0f", x"5ace4db7f5ad9cd6", x"3d51ad3d2a553959", x"20f39e05362cc2ff", x"1aceca4e15fbc3d8");
            when 15821101 => data <= (x"ddd49ca65fa8964a", x"e6eea9cb23eee566", x"700a8030faace38a", x"c0399edaf85f0823", x"75da7df50257cc40", x"b2ea5a513f946f05", x"06e4991ebc3a7231", x"a250bbb00ad310d3");
            when 5867123 => data <= (x"facaad57b9036acc", x"110340db8b6d252a", x"9d4fd55fc6f98785", x"444cd1e388eca46b", x"7724db3826dcfe19", x"d47308a57cdeb830", x"465983cfdeef7c7f", x"ebfbaa9b32ce8d57");
            when 31521605 => data <= (x"70fbed6ec070a9c1", x"e2a08ca568ea956a", x"9081aa6dd12c153e", x"b2a60765407f536a", x"988f43e3587af04c", x"d8f0ef024f1ccba7", x"1b2bb6808fedf09e", x"7f85dca1daf1970e");
            when 7364645 => data <= (x"54fbd0bcaa8a58f9", x"18bd9ecd73d78a16", x"da7825236d420fe0", x"a0a39f4fcc2f325b", x"162ca9e8a0527d69", x"df2b00ec2849e701", x"5ccd8ddd5f2a06c6", x"b242dc04cea5398e");
            when 3266962 => data <= (x"11ddc7b678694c42", x"9e41d23793fcf4a2", x"2915a76a40eadabe", x"69b4853deaa1cdf5", x"b634d0d3e18850aa", x"00991fca92735b0c", x"1e1d7744bd60ef36", x"4d7f8b223c83577f");
            when 17423575 => data <= (x"825a262da2260d91", x"f69bd2d6efe89b94", x"b39d184b942761cf", x"6107df779c3d3550", x"7decec2e768ace9c", x"a2d9358bb93bcc97", x"fae0c02d3c92ef24", x"018165d6b309dc88");
            when 29201298 => data <= (x"fa693656b3207ae8", x"77aa3fcfdcd27ee2", x"78da5da804f926a6", x"b27a729bcb1ed10a", x"c2c609e41ae37198", x"7901bcf64313807a", x"1aa53be820c8d814", x"3813bf5642c349a3");
            when 1333448 => data <= (x"f4eeba0b476c2878", x"68e590bbb0f4bafb", x"535dcd8bd1ef834e", x"b535d07ab5df6a2b", x"bb760a75c1041490", x"7030b495b514bb82", x"2382560c0e08abd2", x"0f4d730ccd68e002");
            when 10281945 => data <= (x"f8b9fb3c3fa192be", x"f3ad4307833a4456", x"4904a13fe387c7ef", x"7d65fb7ac3155b0a", x"8eaa892b843b28b4", x"31a6bec62c523b6f", x"b14fa780f8f9574a", x"80624e140c947e6f");
            when 16337766 => data <= (x"890234e872cfa0a1", x"20ff25cc5753d202", x"5e021c06d57ba8a8", x"2afcbceea5298f0b", x"fbd5c84790d0da01", x"b287d082c2477df8", x"057f2c2ff8e59996", x"61900603060e369f");
            when 26197173 => data <= (x"448609afe6e735dc", x"fa728b05a6ce565b", x"598a44f717601acc", x"ab0912599d283f5b", x"a9c380b9775d97a7", x"810dce72d0d95c87", x"389a7c95dc53cdb5", x"f211d7c046e221e7");
            when 13353730 => data <= (x"8c684b9c07d434fb", x"ca931923eba98f38", x"4a2af18857f8451e", x"8aa8091ce3ea0c81", x"5ab5991528e1bc48", x"b2d6536edcbac147", x"01123898d531a88f", x"dd7b0b04ef4aee84");
            when 33183201 => data <= (x"0206377c6f82a49f", x"5dfa0962608454f8", x"ff79fa7ff0ed5e55", x"b08145ca05be386d", x"c6d8b7b5bf528d52", x"d16f3eedac6c39a7", x"b07f29a007882843", x"b8494b12cb1209fd");
            when 31269317 => data <= (x"3153dce4601ee0ee", x"4111fc234e2928b4", x"3a3e47c2d46925ce", x"7e2675057bb967e3", x"d18a5b3f8ed06967", x"ce3a3de0b0b537ca", x"e5c9fd2590fc279d", x"c2980d8008237cf3");
            when 622993 => data <= (x"5d6f8b6839f9ded5", x"6c61073d247f1506", x"8251c2bcd9580564", x"6cbc9e4502391062", x"5b0279251c28e348", x"12166df090218881", x"75a09271092d9587", x"7c5ce15972d43285");
            when 28350710 => data <= (x"7be96a903efcb7a2", x"df7da46cfd67e087", x"f2353235114baee6", x"e618bc0f8e907afb", x"6cff6c9faddce282", x"b045548f6fea7ed9", x"88f0aec086421bc0", x"cb2bfadfad37f4aa");
            when 20037990 => data <= (x"9e1ebf0719fb20bf", x"7c4a0656aa91e6cc", x"651ebe0bc6d88aee", x"68bd8387a3a502f9", x"d56673ec22b34143", x"a8459833f4829450", x"9d738d5359846d6e", x"897821af3bd32df2");
            when 15492987 => data <= (x"12231a4b98b17a03", x"c6af48a6c3a5caf5", x"21c25490cbef3104", x"931fb244965c844c", x"54c2ac62af6143fb", x"e8b22013f99f3828", x"4b7c01588a23694e", x"a275f5b7b79ebb6a");
            when 27137579 => data <= (x"a23b87b0d9fc3884", x"5982400ff615bf2d", x"aa2c07cf6af5a134", x"c3f7f72cd91d2ea1", x"0db97f0cdf98f0d3", x"058946a45b5ab5b6", x"18bc002ad37d7968", x"b25f8b1dc3f157f9");
            when 789283 => data <= (x"7908a11aea9b1f30", x"094ca3ba52d734ca", x"f8967313e92be28e", x"565655e2b30b77cf", x"04f47c9f4d07534e", x"c82fe16f1cc796a0", x"2952b926f87bd5fe", x"052453022b34a6cc");
            when 17095138 => data <= (x"91f6d99931dd51a7", x"01e7ae756ae1db3c", x"633b2ce636ae326d", x"db222fcccfe129d0", x"5b6d1a4e44224dfb", x"240df739339ae993", x"2c68d1777c84321a", x"e120c7590eca0b94");
            when 10936306 => data <= (x"4680196ccf0d28df", x"88a1e699f449d9a5", x"a912fe3b275f6944", x"5313b1eb8e9e5eb5", x"a4d423939eba2a59", x"944fd9cd0144e0d4", x"e5e0d4eec090523e", x"5a8f33727b06cebe");
            when 25772366 => data <= (x"b182f14b45208f1c", x"5d20688e82dce0df", x"a2699cd4d39dad8d", x"d6a2026106f09043", x"983abfb48b1f529c", x"7a948fae145d1575", x"92db3ea64e68b94e", x"8af3ce834430d2ca");
            when 27386171 => data <= (x"6cc6a8fc090a3599", x"73bdc79055f8088e", x"f7df677db116b37f", x"1dc556d7a8ef1cca", x"773c1e56f99bed16", x"7142e53c90fa5fe0", x"4206ab10dade3339", x"91dc77a262171e9b");
            when 25524278 => data <= (x"ce839c38a88b152c", x"49313e3a857ec8e4", x"75152eace736a047", x"d8b1b40203a646dd", x"c4ac143cb0f936ca", x"68cf34f8382840d8", x"15c2d5336931f187", x"1a06290616b51c79");
            when 7709258 => data <= (x"792b90a516c5da89", x"e5f9322daab4f868", x"d409853a97c7ecba", x"98cedd73728ddff7", x"854249e3af555e3d", x"425acdd579d8b631", x"b8a094c81a5ce802", x"2c06ae0865f8ca36");
            when 33412122 => data <= (x"3aa8cd32b1034731", x"d01029969564e5f7", x"da06025125c6a8d1", x"23d3f966c0118582", x"01de051ff1af9714", x"c9273bb792a07411", x"5845fe573a7613b5", x"547aa72ae56d1a87");
            when 653857 => data <= (x"74f602448354ad30", x"d2d5f5cbb3650230", x"019b5feb63c4fd0c", x"fc3cbbfea5b18be7", x"7958d1725e2ba544", x"769d81de33dd5d8e", x"6164ace82fbe3693", x"0c2d4e72d3c13199");
            when 22507917 => data <= (x"6b7234aa4a4d4c8b", x"e34cb2aae09f0952", x"1ba97bba68f93c18", x"197e146b51661c55", x"d6c5d6579744cc7a", x"76d48ab133667825", x"cd5f5c58aa9cc947", x"b44612cf294488db");
            when 18464383 => data <= (x"45be40450bfe2c38", x"c24091a1e10a5d81", x"a7eb81d7673b14d0", x"f263ecce296c7fad", x"51ab1f36036442f2", x"9f19733918445d77", x"73567248df90559e", x"fef36ff7453596fd");
            when 7109507 => data <= (x"f99eff1d30408b3e", x"492030487d9360ac", x"ca676de788643cfb", x"1a8a9c123edbed2c", x"1d9932a731399849", x"8cffe6592ce17f71", x"c8947316fc730ed7", x"0016afd0505cdbb2");
            when 25201197 => data <= (x"6e8b540ca55d180c", x"07cf2713c0a8606c", x"b8e8614ea4e4c3bb", x"4e882f9d52348108", x"36386d96257f212f", x"8cb993cfa1a8aa2e", x"38d32d91e5d1ca4a", x"29ffd227c8b8d1d6");
            when 1576372 => data <= (x"4d5ce2c93069ca14", x"eddb2138fccf7116", x"769ef74701c26b9b", x"63ad3337e90bec2e", x"0a187e1868184e57", x"f6a46c6cce7a4fc1", x"9755604cb8a3abc1", x"d1307698cbc300aa");
            when 30974187 => data <= (x"28d7ad078fd55d55", x"c314ab95bfd4e4fa", x"d0f7a0a8ce3f6a9f", x"557cfc60045ea59b", x"8a42dfca4b478d51", x"0cf60459acffbc4a", x"08a717113f687551", x"a8622c94d50566a3");
            when 20089517 => data <= (x"ea0ac4da1175b253", x"fa32de0162d4ff7a", x"56fc7699822d7b92", x"a345cb39ce6cc58f", x"3e28adc64923c854", x"48428ea067881c87", x"96003231df27f56b", x"25c641253f6e6008");
            when 16904162 => data <= (x"82c13bf21b90eae2", x"bebc663edc00529e", x"4fcbcf15c68911fc", x"91b6168d976ad228", x"dd1bb3fcc572424e", x"d9b568a00af77404", x"3fbe1e3e2eedddf8", x"eb93be9392df8128");
            when 17769077 => data <= (x"4e5529aadd6cb241", x"d7d396f52a84bba4", x"ab6793895b1eac85", x"e3bd90d693862f9a", x"d1f7477f2640b38b", x"d9bfdf2583a2c32e", x"88bf8d0b5f4a9ed4", x"21df71942b224f99");
            when 23732147 => data <= (x"1ff7f267b94551ec", x"a82a17597b4e6513", x"545e86caf3bc36a6", x"2ae526de599d6fba", x"4490eee3be7a6d40", x"7e7144893dbeda73", x"fa7ef8de4e4290da", x"8e9b00cca6031042");
            when 26109723 => data <= (x"efaa440bfee767e0", x"3e09d8e3f2f8c698", x"16f2b012cc3dfb82", x"f3aeb69dbfabdfa3", x"578ee8730e80848a", x"7c1bf8e81f41371e", x"087f7aae8dbc2f45", x"1f32fd23ca92c7b1");
            when 19010398 => data <= (x"22477418dfda93cb", x"46503db814479e18", x"59e4ebc6034e18b8", x"c7242749ec31a8d4", x"80d16e36dc6127dd", x"7b2b5977b61e0440", x"cdb73b693774365c", x"9e6c56cfe8c516dc");
            when 18089175 => data <= (x"69ed614591b97546", x"d4e6154b4a878228", x"5745176a12ad78e5", x"e869292a07a3ab53", x"e097fade73af4656", x"561245e4d692c528", x"8e7532e5091e747a", x"6657d52fed1105a5");
            when 31090970 => data <= (x"d0e3b7ded0336289", x"532f9a6a24729fee", x"af151d516051362d", x"20e6f8b041f01314", x"18782f3a8dbca99d", x"d7fc77e11ece9647", x"60ae19f05c3aa569", x"897ca9c99ae0e4b3");
            when 3333028 => data <= (x"9955ecd17d6d2452", x"1f5c8a7646e9fcf4", x"d9852afb3b54dac8", x"a8e76a25e556f412", x"4f6b5928f01fcd46", x"69deb102d78dce3b", x"74630957a82a6ec7", x"cdc0506a6e00d4ec");
            when 21423030 => data <= (x"b21b2a11391fe6b7", x"367d541138402d91", x"5b151bdb30948fad", x"453c36fe4e266401", x"c1771a1191adf796", x"7c6191e480694ff8", x"0e03fbce9e7cbf33", x"66c8e0b242f02f97");
            when 7658230 => data <= (x"6fed85dc1f49fed3", x"095377f6ea860d36", x"354090648a58a5d1", x"f6788c0b9d56e010", x"eaea5fd42a05cc5b", x"0d71cdafa8ea6c0a", x"765caa17b011e5a2", x"00612e518881d2f9");
            when 4493132 => data <= (x"179ed702d1ce538d", x"14bd5f945d32ac0b", x"a27ae579a561f64c", x"5cbfc4dbb6885e9f", x"0b57b8b38ab951a7", x"b117af3545f00cc3", x"02abd74119513180", x"cea6970eb1c33b55");
            when 21638192 => data <= (x"cc5c996f1a2df16e", x"dbf1face2c920a75", x"e070b0dff2f5631e", x"2080cdd3bd157a79", x"5483079b6548c37d", x"9b0b8bf1f5222b67", x"f37cee02d0489b55", x"6f11ebda039984eb");
            when 13698145 => data <= (x"766ec46fe62c11c1", x"0c0dc359e208352e", x"581eeeb05a9b351b", x"c9aee72b4c05e578", x"a9fa5972625da778", x"2cf7d1124ce070da", x"605011b647497566", x"77f6a34e4baa154e");
            when 33043648 => data <= (x"67871f418f295739", x"c3eeee8999c8332f", x"8a464d60db39fb17", x"5fbade2e593a94be", x"445b4a71bf6c231c", x"ea4607af64f292fb", x"1c9719fd8f2088b6", x"ce25d5cb46c7a5be");
            when 19499550 => data <= (x"6e52b7af1f69b209", x"d4156ebfd8f1219e", x"f58a927d7c9efba6", x"18358fc8667fea6c", x"f8d954ae67da45d8", x"e1c93ab8b5eed654", x"b6a2d83ae18b7938", x"aa506c67459babe3");
            when 24499588 => data <= (x"68082af42d8e64ff", x"5177c8a2e5c643e8", x"ec678ab1ed70e3a2", x"861bf905e66e4c57", x"77be89a51912b90a", x"871d3e325414f4e6", x"5cd0da93a33a56b8", x"a35dede3d8807660");
            when 24697413 => data <= (x"67c31d5ea1900bf9", x"d7d1ad09c81e59ee", x"388dbf71e006c98e", x"db202a0931cadef3", x"b571c2f0549e0580", x"6f3fd6b7b70948fd", x"aa9a8a7fcf098184", x"55b9dbfffa546538");
            when 24543603 => data <= (x"0232ba4a7fb9f667", x"40a002ef018abe6f", x"e5014a01db0fd311", x"918d3455972416b2", x"d2b2c54b16f996ca", x"395e6988fe88f746", x"d2ac8f2ee28abc6c", x"3b93b0765ac3b1e0");
            when 15387896 => data <= (x"82006184ba2027a6", x"ec190242fec69cbe", x"a387b664459097a9", x"e0e17e4caac1a2e8", x"5847cd8cd993c169", x"81726c6b339041ea", x"6185f19b2929fd0e", x"c6843ee63a00429a");
            when 6879332 => data <= (x"ce254ef68d451944", x"da722695d2f7a2ec", x"33e324d1dc253b70", x"508be99273ea460d", x"5dfe5dc5230b3128", x"4fb8f3c4fdeefc9d", x"e18714924f32fd15", x"51b41ca4d899dcea");
            when 10495921 => data <= (x"b1c1b6a98b98b432", x"12f9f5e5b5e5f1f7", x"adac2cdda85fe753", x"765cda79ed76e290", x"8c803e5f971023d1", x"f56c09dd7993de7a", x"4dbe6d469157b5a4", x"6aefcdad60cb3b71");
            when 28176710 => data <= (x"6319b115bf6f757f", x"fe694923afc0f846", x"b415a05d7e26749e", x"59dc699dae46abfc", x"f54b7be16f8708f5", x"5cc392d3b03a2c36", x"c410b4f66617a15a", x"2a6d132882183ac3");
            when 2796519 => data <= (x"a7867b4bb9c437e6", x"9f8fd950681b57c0", x"824c755fb0994e81", x"44d63a86677ab506", x"5b3635cb1baade6b", x"db7dc2a72e3c16b4", x"2f7e84bdbe4f2593", x"95d55a6f249962c3");
            when 7485442 => data <= (x"f6453c093f78759d", x"d80d7db7b2c55ff6", x"b16b7d14f4d7ed18", x"cab5970cfa95ba00", x"02d8f0d4a0ace622", x"066bf5895515038f", x"bd9d8f47258a4429", x"779d060f9a94fc7b");
            when 26789150 => data <= (x"bf907ee17de2d8ec", x"e3c5162b8e65ce11", x"82dbf06c94e7c7c5", x"584e59e4b15e7663", x"744f287dc0dafe5b", x"7ccd4d64f0829bd2", x"f9d9d98be62db86f", x"899bd070656434b7");
            when 14060677 => data <= (x"7a4aea2702e3fa11", x"36d458cf1b44eb94", x"eeb85c6e07f288f9", x"40662070d0871e44", x"10f82e3fe6afbf2d", x"fdc631c0e069181d", x"4f303f269e0d6341", x"8ffb4db2cb843308");
            when 16360696 => data <= (x"db350537fc09a898", x"825a0af01dc83cc2", x"b64d9b9faae6f747", x"ccf61db23a9a6e1f", x"2013b9a4366341dd", x"739a445722c0e070", x"713a5cec06ec00f2", x"77a37b641365ee54");
            when 10732384 => data <= (x"162fd46e6d3ed691", x"b2b2393f96ce4580", x"a032be579b938a66", x"9b4372e63d137f1d", x"594753670d9a18ea", x"2e88c79afd4b4880", x"5d9cc7756ea4e908", x"4016dfa7bd82215a");
            when 25343312 => data <= (x"893b42d74646a15c", x"573bc8a5ca20cdec", x"6921dbf350a17271", x"3dc35a00eb0ad85b", x"d90192187054bb8d", x"9a1caa04d680ea47", x"8d633528135e586e", x"8d545819bbfb1fe7");
            when 28275762 => data <= (x"33e872181006aec4", x"0ae1fcd24ba8e694", x"04b79d449ca7531e", x"ef1e87c0b327c270", x"fdfcf2fffd3e3039", x"b8c5eb2c55078575", x"84a76007e0c1663d", x"8189121f22c2c266");
            when 10556360 => data <= (x"81071a0fcf1a2392", x"f2c37bcb7de147c3", x"54adde05783bd1e0", x"cb888f4d8547e484", x"d066086d9987be6e", x"0d301809dafa360b", x"4f4fbfc4a89390a4", x"b8ed1e3a488e6a24");
            when 16963431 => data <= (x"935050bfca829ea3", x"7b1a9fdb060a849f", x"e5a25f68beea4d3f", x"1c8f394b9907a239", x"c4568dc4e6c3afa3", x"17e6810ba00a164e", x"666ef709f22f7f1c", x"daa26cec4a5c1f97");
            when 26919456 => data <= (x"fd686f4095596657", x"ab780be5bb6e89aa", x"ff7f279117e404f1", x"0b6626f9d792d241", x"a180dc8cb852481a", x"a612f3077c1df716", x"f4f29b6333cd6bd2", x"82d27787fd37d6e4");
            when 9655700 => data <= (x"50c38377eec6b5af", x"92a1d616b3cf0e74", x"f118610bd078ac3f", x"74ee9e3151b28264", x"9bf5870fac6c3545", x"cb94c1f0e299b7b3", x"16a9dbef29ef579d", x"233714e196c08849");
            when 19686551 => data <= (x"08fe6591f6ccd931", x"be6867f59670b0cd", x"40f63a4ca6e7ad74", x"a014cf0187a53984", x"a5b6f7ebef4b63a1", x"5a875c2b012713a2", x"832fc218bc487e0f", x"3b732f5f5f3144f0");
            when 4317184 => data <= (x"7304157352c66433", x"a082289148677246", x"150548da2d1efba9", x"50d55e50f1aea574", x"9225d91a140259f7", x"4cacc1f2d2fb6337", x"89164685498a47d5", x"5485b47060a09ff2");
            when 832878 => data <= (x"8a2f7232d8f3430a", x"d685ab57e8576dac", x"90da261fb58abd36", x"d965434c804e747a", x"21f259bae9f56560", x"115875d14c881b41", x"3bd206d43365b306", x"cbd84805b0fe93da");
            when 18706769 => data <= (x"2af65159e6933903", x"fcb85b665978c47b", x"b84ea0e59c7ec6e2", x"541c83e97445528d", x"09c7de82e5829ace", x"bd36c0bf6beab973", x"35e4c130b31347cd", x"9f5a1a5639d83a26");
            when 16156637 => data <= (x"986d18ce5f195e0c", x"f8808ffaa0e83826", x"0495894fad611536", x"94b8f3474e9bb646", x"13454494491c3098", x"381691c2fcc2e8d6", x"d5a50c6444308a66", x"3d00ab6e5b65edb8");
            when 1567820 => data <= (x"e5d4277546e9b4f6", x"dd86cdb7a328d893", x"b0478dfd86759d34", x"b4b4f45a5b044a10", x"06ad2efa411dc583", x"1a0b04f20fb8ce9a", x"51327541073211e1", x"6bf22aabc47e38d1");
            when 11265709 => data <= (x"70c7b4b34c4eb0f3", x"1b8469fafbfe25d5", x"96aac55d7c092c5a", x"752fe10fa0ac929e", x"7f78fe8585859522", x"efbaef0dc4b81ec3", x"16e47bbafa49b551", x"4fe28f0d1febd598");
            when 12961871 => data <= (x"a8dd8e65e82a764a", x"94e2ddb5b2af0162", x"96543ccd073d528e", x"c473eb8ecd895537", x"3bd799d46b1d9471", x"a235f3c7f439e221", x"bb956d958ae3d315", x"673701a27f9e35b5");
            when 300368 => data <= (x"f6f93c5a913a44e3", x"d4977d58cd18c63f", x"09bb4da345a27472", x"bc887593b259c7ba", x"8002fe19bb1b235b", x"39bb5ddf11e3e518", x"72860118a2a8d360", x"e21c14b8632b3ad5");
            when 11499734 => data <= (x"48781ce6f73ccfb6", x"d2bae8355c9fcb83", x"d96d9738a5ce16d6", x"ecd2f64a4251d752", x"074ebd4f42dcd701", x"653cdb7f465bd2b4", x"9182b23ec2074ee3", x"08b98a9625eae27d");
            when 25662110 => data <= (x"35b185ed44de16ad", x"296e1cec8591acd4", x"1685bacd190d4f37", x"79f58bd932516f56", x"c4aceab50851e6c7", x"4a831411c76978be", x"f1d85d34294748d1", x"5472859edd536465");
            when 9312282 => data <= (x"33184a89378f16bc", x"0242d4a7f99a8c43", x"aa2c87adad4d7409", x"1f7bf80c3ddde2aa", x"716506e8d775872a", x"f9227e47c262d09f", x"253099f4e14892a7", x"007ef9a2a13814d3");
            when 10943588 => data <= (x"2cb48dd84a729c74", x"33519b0370a5c273", x"5f273c4c39a633fa", x"2e82a0ee11b9a5db", x"5b24f6aa5de5335f", x"32918f5237d3a4e1", x"cf0c35d58034f8b1", x"da2f3d62b71dccd5");
            when 17156427 => data <= (x"8d49b319197cc292", x"51bbeec05f814c6b", x"b385514b492c4fd5", x"eeb378dc099197e3", x"6c550f59dfd4654a", x"da1970e4a7041eda", x"63cbfaba7a27f47a", x"884c8dafbaa8edd5");
            when 2299349 => data <= (x"71f017417c4a2910", x"5f0d6913ec0ab0c0", x"89a4d51a8ae5e4a1", x"2a2f4252b4455d43", x"865b42e9c8da3643", x"f871f24f71f93583", x"2b307f5b1b1b5950", x"301f59dc8897ccdf");
            when 15942910 => data <= (x"8ba0eed4c448ddff", x"774e17280b634a72", x"214e8d8d673d38c5", x"2821978aea46367a", x"ee2d0b6abbd5b152", x"a79fe43b6f3e27a1", x"48e0662d0d1ecb42", x"397c83bddb1b55ae");
            when 5342402 => data <= (x"062a4e60714429f2", x"5cfac224ecbb7b71", x"ae47c39be9aac8a5", x"0eb9000e80412afb", x"33fee17be4a78985", x"dbc0ef58ecc5e02b", x"5498a82e2f6c9c09", x"31b55f50c7cc8fdc");
            when 8732558 => data <= (x"e805e3d4785d7a5e", x"b3b0614bfe662a1e", x"3cbdd725a948aa30", x"d339ea8ded0432a5", x"783a2898674ac284", x"4d83b18b58a7efec", x"1ac9e448fb447c23", x"7f3f9924f7fe5472");
            when 1964889 => data <= (x"beb8c46058028465", x"4a9328f66a57e31a", x"6d65457c35030fd4", x"53c641fe4d84f4db", x"9e68aca82c4b78ff", x"a52ac6c9a4229bc9", x"9571ec1012316c88", x"52f0c2fbe929d599");
            when 7551777 => data <= (x"6ee6ccfc4dd65ea8", x"8c57039f7641e8f6", x"792c41527a9c8a28", x"24b6e564ae768ccc", x"9653acd59a1d3213", x"243cb27ea56dbfba", x"155ceab5d3a34b7d", x"b964608937d988a8");
            when 9875430 => data <= (x"ef744da9897b3461", x"b82ddedcfa4deba3", x"6dfa1c51307f9242", x"2a14135525f8cad7", x"e4a1388400866f4b", x"10eb4b62b9459be3", x"17736d745d5da84c", x"0881cae607e29df0");
            when 19858383 => data <= (x"146d6284cab9e406", x"5356d46d48283430", x"676073b427a4ae83", x"7c67aeb567f4e4ad", x"797a6cac265925aa", x"25b45b6b5f48d81e", x"38cc041f0ff4f6f1", x"912bcc6238b04738");
            when 17999346 => data <= (x"0d010b15f5fb5442", x"398430e6e04eeff2", x"4c26df91a7418cf2", x"12ccbde718e85aa3", x"aa9745728e7a9849", x"5dd1f0cb98e87090", x"36cfd0887850a826", x"4695694dcec8324a");
            when 23585717 => data <= (x"4577ab7a07141222", x"528971c566bf0675", x"9784dac50471c04f", x"7fa5ae11a5361696", x"a60db619e6b67cc7", x"1a91b048a5f2de96", x"5618f54732053c99", x"7a4f6dc9187fff14");
            when 23131438 => data <= (x"2ab4e62ddf59cafc", x"178d1947a567ec46", x"18bfedf7d724308b", x"f8437987512833d0", x"4f44618ddcc4891f", x"4fb39c7448d3ec40", x"e69ca8d4fb235272", x"62bfef403ccfc415");
            when 25201764 => data <= (x"ecce01ce5d57cf42", x"d5d837e12ea6bd93", x"605d60ab055fdcfe", x"e7c1bb3fbf66cbbf", x"4c2ac0effdf09de3", x"8c41e69cb104d5dd", x"16f74252362dadaa", x"1852c849ff2168a0");
            when 11840861 => data <= (x"a06494dc93bad35a", x"1199981bf998311d", x"5e2a861f2bfb5e2c", x"dbb3f3300563aded", x"6d5c6784d48f835b", x"7b4cd01983ab27fd", x"c997ef5405deea9f", x"ce49acfb6800c58a");
            when 24199792 => data <= (x"d8625e8637abf9d2", x"f53c8b5c05ad7f41", x"c84e3057613e8716", x"cec904348507e2c0", x"4598b01b59be9d90", x"628a6e97a8127afd", x"44fde51a1916231f", x"cb6d3484659323bf");
            when 2434573 => data <= (x"c27604d14e758364", x"7e2bb8f07415af48", x"93f723b09060bc55", x"1255f5ab1bad92d0", x"65f56ad5cdb6a399", x"af6eaf07980c9a23", x"3714ef7a7a5243a9", x"0d37f4e8e38ba0cb");
            when 13403855 => data <= (x"ea22bd3bcf620d17", x"e7d6678cdacdf5b2", x"7e32b1e54289dcc5", x"25c39b367892226f", x"f60783824857e781", x"bb9b7fcb03e1b175", x"cd7005826bf11e4f", x"d2f423fcab575375");
            when 31821408 => data <= (x"42c90654f2ff7f11", x"ab1b7beed1810a98", x"cedefdf548e2a87c", x"8c852e61b0f16962", x"af2c8a24f0a5f53e", x"6e9a7f077a0ac2eb", x"1e92f75d076bd098", x"ad9c807a0501d879");
            when 30818874 => data <= (x"e8e6e8445c49df51", x"6770e0af83350204", x"dd3cd87b5947e4b5", x"a5684615fd88cb3f", x"9fb95b1621a5a845", x"fb7c73a4d9d96eea", x"21770094ca6038d5", x"e578c0e5f7df9935");
            when 6889244 => data <= (x"e453fc553650b35e", x"c2ee3abe37684d8f", x"a8738df333544e9c", x"fe55c28470ade100", x"c7bf8f39fa37b097", x"d7317c9d52150151", x"3503bbcd5a7c4024", x"4343235f9a95d3a0");
            when 16282379 => data <= (x"9182721342f147ff", x"90cdfafa87fb071a", x"d283bdb6fd420f1e", x"ee3fc6f020c6ac64", x"d5ef35a4e8ed3f5b", x"ad833350a5c094c4", x"cb1c26559570d391", x"203ed506e4743b03");
            when 24498884 => data <= (x"e82b5c393be521cb", x"cd61a00b8abead28", x"656a116dd3d94821", x"8f637b0caa74e480", x"a83b9fc5d78f1949", x"92019a7dc3131ba6", x"5e11c17cd5c2e291", x"d2c9e4c6456cb4dc");
            when 14863574 => data <= (x"444433e47efec6f9", x"bc12796cf5676667", x"7e8f6e891c9672a6", x"4790d7705902fcfb", x"93bd0edc592d0d1b", x"e75f58760501fd99", x"5a5c8f90a137f22c", x"ef4f9527ec4d605b");
            when 21355402 => data <= (x"d872d10f92c56698", x"bb92f9009968bcdb", x"482fa75f96f92510", x"4cd0c16d67217e50", x"197d9567e6e0fa2c", x"0a7822b7cae17709", x"d741679dcd6a6f6c", x"80ce00ebeef1beb1");
            when 11697625 => data <= (x"eae983635a28e346", x"ceaf740c8624bddd", x"e1cbadde3df79653", x"e4bb5e5aa7353093", x"6fc80be263cc3d9f", x"0dbc71f26ba44ff4", x"286f98de31a47b5e", x"8fb694cce98f931f");
            when 20367888 => data <= (x"608bda8ca1b4afac", x"258fed35516e5338", x"c1cd6d17e7f4ce19", x"7d66f5921cd2c2e7", x"578ec6879bddd51c", x"cb17fd30cb8054ee", x"150ce25573f6efe0", x"1e67860e769533ba");
            when 26197884 => data <= (x"9f61b9959802282a", x"40f1c9566d35b1e4", x"c9d7b82509582564", x"1f0ed67ab45b8370", x"6ad5e29bbafcf588", x"624c920d69ed21c3", x"aa2048a39e778ebc", x"a38b0f19ee560134");
            when 3525876 => data <= (x"12881cb1b5306b72", x"d9b2a6404931fdf9", x"5c9e923c93ae3975", x"351da5ad90366a73", x"8dc921ffa8ee17f9", x"77268c7545391600", x"ba2d7a616b2ebd11", x"11f3c6a9653fde02");
            when 30221126 => data <= (x"fc1cb844d1525ae9", x"9c2b018bb9a65463", x"21d1443dcd25546f", x"211c0fc0dac9641b", x"c39f728dae9cf4e8", x"44230436f3778dd3", x"44ecd79e094aba68", x"b955e6c24860936d");
            when 9015448 => data <= (x"7a6d18bd2d73546c", x"af54f9d18c4fc8be", x"2c50d4a19ca862d9", x"484fedb5035b2150", x"71da03648701e6a8", x"bb692661ddaf307e", x"a68f4229483fdd3a", x"0f71c11b303a6980");
            when 4521881 => data <= (x"11377f079bc515ee", x"c29bfaca3349db15", x"402bdd462e67bbd6", x"9c42beded5915a58", x"71f6bef531ea3437", x"b2cf2bd866144e94", x"b356f1e0462fba06", x"6d835cd6bb0bf28e");
            when 20159410 => data <= (x"cb0d2a01747e1ef3", x"8f58285c87c5ae16", x"02ceef327dc03a7c", x"dbc9afa70e5901ba", x"73b7574907ee1d81", x"a8ac68ae0d8113f9", x"ae1d39d52dc00ae1", x"78eacd35a69018c3");
            when 30316000 => data <= (x"5080c73176aa12b3", x"8e07b640d8a849a0", x"b591447b7f6be098", x"84c42684b56206b7", x"456462cfe798fe72", x"66faf3d451892a77", x"f199dbc63699cb38", x"71f6ff9b8340bea9");
            when 16317987 => data <= (x"af277274d2ddc161", x"0f48e6a762991f84", x"9ad4e796f66de395", x"ee6aa7212d870ae6", x"f8a07c91850736ea", x"4bbeeefd80524640", x"f6156fb77a9ddf25", x"0cf217b99a68c884");
            when 19525723 => data <= (x"e34be7cdc1ff0235", x"9005774f1fe2efe7", x"8578065488d33250", x"f0ef0dd900ab1207", x"9c447b504df6f4e2", x"ef188d799e52da85", x"4c5b9f1b48571aa3", x"c78d41b93add1821");
            when 31741408 => data <= (x"61d2038ba320fccd", x"49b4fad68a57f92b", x"175aa1b3715ccea0", x"c6bd9a1b83b974bd", x"66f3722dc0018384", x"53840d0cf4158d80", x"f0354e48486541c8", x"2c318649554e0ec3");
            when 29024172 => data <= (x"4717a1637599364d", x"859144d31d8eff2e", x"ecc5c7fc77fb9d50", x"8812026cf7919a03", x"6b441d18bed40310", x"337a61bb053b5314", x"979c1cc6cb94eef3", x"b016c98d5295bd79");
            when 24700859 => data <= (x"6b058cd5a347c558", x"ecdfcd7856e8f9cf", x"b5ffda925cd5683b", x"7d779b3ca902ce91", x"fa62bd59b6c8bd46", x"66ea1a88bc99fcc9", x"5d9546949be9d5fc", x"d659d895a4ced948");
            when 20340607 => data <= (x"f024a4fba2d2c2b8", x"4c360947201ed40a", x"21a681fb63c4ebf7", x"ca2cd188b261ff7c", x"b22d932792d08c8d", x"f86f76d8d5cd5a72", x"ad49224409457158", x"0810ce6ac32a8088");
            when 2869684 => data <= (x"33e284577bd0f3d1", x"ee8031171da41fe5", x"cb7d4fd8c0ba1cbd", x"837d6e0a6f529263", x"494f39c1cc909f5d", x"03e2c4b1cda2e180", x"34d138352ea125f7", x"de52af426a2b457b");
            when 1947580 => data <= (x"67155819f608d85a", x"20242afb9d26f547", x"d2118f6e1304ccd5", x"36e1747876a9f020", x"9495bc4c26f2965a", x"78671e59036c2ba1", x"c00c7a349aa2497f", x"1f097927f3c4463c");
            when 27574813 => data <= (x"db791bf61f3a5b85", x"169a9e075b930fde", x"e21fcba39e727f2a", x"d49af65b6f007eb8", x"27076ce7225a4cda", x"eca87c70be688de2", x"36c53509d0dbb1de", x"0fe26c45f32925a8");
            when 8791045 => data <= (x"2a73515283bbe955", x"4961938085c3145f", x"fa98b0002dcfff0e", x"bf0f4b0e45030f73", x"fe05ce9a66e6a9f8", x"074bb1b63c4ae61d", x"d0e09bdeb323c0e9", x"14016c6c82c4e8a5");
            when 3898330 => data <= (x"fb6f7fb14761fc6c", x"ba9b66e81fb4f683", x"b0d6845f172cc0d1", x"481d3a946ac7873c", x"9f46bdfe0353dae4", x"ccbda4f1fae9479e", x"9fb2cf9f0a7df635", x"170407c245ff84a0");
            when 25273987 => data <= (x"e69c215685c8aec8", x"3a31d5ca35e6ca97", x"f8013b8026c48ae9", x"eb2ffa9455abeacc", x"4e6bbb821118ec0d", x"863dcc5c89405281", x"7041efffec6ff3ce", x"9740ea818732ea0c");
            when 32264895 => data <= (x"102604362d128454", x"1ff48a1ca5314f7d", x"fc419cbdfaf739c3", x"92b756abf71702c9", x"e17ffb1836f55c6f", x"2d896d8a41a1835c", x"0d3268b04191abf9", x"73ee12357325feed");
            when 26572524 => data <= (x"235ca8165884c0c1", x"e3f14960b3e42eff", x"9d67f4b4c7eff307", x"b8a2039853322cb2", x"17d3ddadbb6fc206", x"bb1d3a4c9fb23926", x"9ef61a1f37579a1e", x"d6b62cc1bd1c4e08");
            when 15549458 => data <= (x"ec1e756a7a025212", x"bcc0ef4ba8a5e624", x"cf55fa2928c09186", x"1ce8720afa5b87df", x"0c6d00a06604493d", x"d8a4750b6e31c2ff", x"f332d91059d77e01", x"e1f49b397c5eb21c");
            when 9193309 => data <= (x"15a314c82727d83f", x"05ee129193773417", x"f84a2548106dc3b4", x"e25fb24a29b76114", x"2cde980467dc4337", x"92c65c93642c950e", x"7b850759efd5ddf4", x"8d7f1beffa5eb2f5");
            when 17539723 => data <= (x"2caae287344deaf5", x"48aa09c38105f0f9", x"62f32a05d563467d", x"7a57cb842830ff08", x"685e9beeeafad37f", x"610c35732da3f01b", x"7f94287520c65b11", x"1c7a39786b244e78");
            when 7617732 => data <= (x"479d40b780fa0915", x"16e8fa5d4c1d65d7", x"96e61e1fad612f1e", x"821aefd95c716537", x"592eebe8a3aa717e", x"84984e87e82d230a", x"12266bbf93994c35", x"d68cfebff8be8486");
            when 7796925 => data <= (x"b3214ad3792880df", x"427f7b2ef73beb7f", x"52f7c24f0ebcda81", x"60032cccf1bdca29", x"7266ab7555748a96", x"75e3fa5a2cd4414a", x"9abb275e4d61abb2", x"bba393dce48312ea");
            when 5222868 => data <= (x"99ad609cb8b88d8f", x"687e7f779811011a", x"529410a28f864d51", x"db4f0dace766fe79", x"d672b33bd0ab58e2", x"9f8e5d15bcc8c8d2", x"7d130b7c701dfd80", x"a41bbf4a9f681185");
            when 16773616 => data <= (x"1040440b162bbc89", x"20d9a290373dd65f", x"dae945b3e7e58590", x"93ce6b5bdc4a52d5", x"e76ad8ffe52d8af3", x"18bd0d19dfa4c6ad", x"241b9f56ebaa841f", x"91b2b6454ede15eb");
            when 27254832 => data <= (x"b0352d9f9587fa74", x"4d7799cb3cf7f522", x"58f1eb2f692428b0", x"8ea0ca44dbead8bb", x"fddd0de5b102b3b2", x"50ecdaa999fd3115", x"0c4019939e74a152", x"9be62a0ad63e420c");
            when 29201861 => data <= (x"602b4bd1cf13dea2", x"306594059d7a0345", x"251f23a470a27e18", x"b0db3ac4436a3235", x"1c5969c708871f06", x"ee660bbcbab2e3c5", x"cbb3beceb0b639c7", x"b7352dbb54b1f1dd");
            when 12401227 => data <= (x"2c736886c16702b3", x"6c609fdf5fd2ce40", x"5d43f9487affc381", x"5ad81a8b14e6f1b6", x"b70b7bf17d9e5a27", x"0178ba5d54848d33", x"1f6c5f9fad17d885", x"bfe59cdca0d275fc");
            when 23022185 => data <= (x"27f493f85934309f", x"735c2493bdacdafb", x"c22db282f8e60b0b", x"07227997d0e80b99", x"ca0aa692c222f8f4", x"b4cd09ca91758f6d", x"f17c4f1af35482be", x"ed63c79f2b52c5d6");
            when 2867593 => data <= (x"5c0a2f2056b683f5", x"b14a391f370aab2c", x"8e83be9306cfc9be", x"dd47eb0e961dde8e", x"4a48906bb59270ff", x"e259c278ff0e8e5c", x"6f6f58c3ceb1248d", x"86cf83b89df5d372");
            when 33018167 => data <= (x"615e04e73c8915a8", x"64dc8c2e14427393", x"023a334aa0e5422a", x"e26defdc28770f90", x"d487746f424e3156", x"50aca06f5bf214b3", x"3df133e5033e044e", x"d6f1cb7aca439d8e");
            when 26027140 => data <= (x"46a9e9632807dc88", x"e466a4b00429c088", x"4ef71a5dffbbeb37", x"e28338c00e2044c8", x"b9dc6d9aae575089", x"f84074b59f722bf6", x"43648806d594dbdc", x"2dc6e61e383233f9");
            when 19083799 => data <= (x"390366fac417db84", x"5293024a9213a88d", x"06b4ca69c451aa4f", x"48f6983adbafaa78", x"b84e74bc920e1769", x"b9c17cd6c1f2c9b2", x"62f245260c3be2fc", x"6b139d3e0f7ec0ed");
            when 33650233 => data <= (x"1f5dfaf472a98064", x"ae716ae7037071d3", x"6f32b91fff5f9336", x"e3186ed2af8bdff9", x"888939ecf3e26839", x"b5d87d0b1ab807c6", x"7a64906ab1f252b6", x"7fbfba99fb4d1f23");
            when 8334200 => data <= (x"62927710eb044161", x"f82c6007499aaff3", x"cabae942812b7ec2", x"0fbd285e9393d8ce", x"abea8eccff38b7a3", x"ac91aba2273f16cd", x"1d672bec72246f48", x"18c878c90f1e8095");
            when 14786682 => data <= (x"59414545b7c6d9bd", x"c3cd7a25d07fc888", x"82720722f63d025c", x"4fbb76c077000c23", x"b5900d273015dcec", x"389752f02855a8e2", x"420b767363082d6c", x"e61c49bb3955c178");
            when 31927944 => data <= (x"e64e43a78b1ec1cf", x"1a18eedbbcdbd9a9", x"53e62eb81c77d525", x"5a58badfc89abd20", x"e4a985f7a4fc5dbb", x"e31c33392c115980", x"f995ac7b0a08af6f", x"6e2e0d7b4021453e");
            when 13561325 => data <= (x"a514ec2687131226", x"d1fe6f3385e70db0", x"7514b9e5ec02d352", x"f5a8500ef3a91415", x"3253bf9895222a3c", x"7c5d08177ff5600d", x"0ba1210dff01d797", x"ea1f04100aeed32f");
            when 4384753 => data <= (x"c764ca6ae3defc59", x"3a6bb58bd0aaf7da", x"e6d54f0e2f763382", x"326a25e2c0c85a46", x"a710ff13840ac085", x"5114a03fec23afbb", x"1caeab94b93c11fa", x"def5478159e64895");
            when 8958634 => data <= (x"cf744fea1cab995e", x"3d090b2368f49fc2", x"88d9c29edce67ef6", x"100462bf7f1d8a4f", x"de82ccf85a305534", x"7bd52457e2448320", x"e0d65d1afc64ddec", x"b32607c459bb2650");
            when 3391043 => data <= (x"2f4bf672a05eb128", x"b53ccef0c7dd9d1e", x"514312b21a674eac", x"746c07ec3688988d", x"13408cafb127da80", x"712ba229f741c918", x"7985fc16e07b15f1", x"5b23f3b84a32d9f3");
            when 21623770 => data <= (x"2e82bc2007ca57ed", x"0d16b38f6d8cd2b6", x"c3153dcefd19af21", x"91b16e7a51f9d303", x"2df1fa1ec746b199", x"a9f822570a67a214", x"045be536d15d66bc", x"05bcebd399f3adb8");
            when 7010876 => data <= (x"1e93d571dffc850d", x"a744065b2c8b16e1", x"f9d39a4997d52538", x"18fd0ad0e991243e", x"7ae3de37f2dbcac1", x"bd3e799a0b8ccfd0", x"1e564886aca65b7a", x"b569bab63f72076d");
            when 15771455 => data <= (x"9fdc74684400b024", x"4d84bbe9cf5c2cd5", x"56763314513418a2", x"f31c88038d900184", x"4446bd99a69b9efa", x"6a8876148dcc2c58", x"4185885b286b21ac", x"3fcffd7da13d9568");
            when 12292420 => data <= (x"cb036129c0a1f289", x"2352ec599ef72ef2", x"19e1e09a2e671562", x"a976a879a13c6772", x"71564daf1f72b7bc", x"ad1793ee554544d9", x"d6c1b95b13b77ab3", x"6c29c121610d8be0");
            when 23065440 => data <= (x"3dd817abc4e73f67", x"c613b0bb75c4e9e8", x"76f1a9f24cab6fcf", x"a18e94d5a2e9d50f", x"1562665629eecf8b", x"8e79bdccae47005f", x"e06f04f15974fbae", x"cce623dd1ad87d79");
            when 28305664 => data <= (x"b0e900642d98e71f", x"2ed292704b512713", x"5e7d34a66a8a7640", x"119369f93db7dc1e", x"52fbf378e0ec5158", x"42b5071ca91b90db", x"602bcbee08e90c5a", x"37a19a20561f06e3");
            when 21697012 => data <= (x"09dd184767207ce9", x"c231b21592e5e409", x"74cb60eae4e9bfe6", x"2a093e658740af68", x"bfa84e595b28035b", x"cf1620a0225711a8", x"34e5abded8318d5f", x"674216c394ee6b90");
            when 25910977 => data <= (x"a5d35f0c65999206", x"7c701e91498ed53d", x"b00157a101d01bc9", x"816de06f01b73c42", x"3cfb90512c246ae0", x"5e53b4eed2319bb8", x"2ba2dc8647a9e347", x"54ac154c1308f71c");
            when 13862192 => data <= (x"180bfe760c272431", x"2b43982ac3109a74", x"8fe05b9d467afc27", x"b3c28e1f1eea3cad", x"4eccf2efe4f54142", x"c7e02aecd05830f2", x"bcf844d838f8ace4", x"3a84fe0b8b98c28a");
            when 15393417 => data <= (x"e21ff427346a3d8c", x"bf5bc3a63d96d718", x"ff51f9182cd4e15e", x"6297f8958ac81eb5", x"30a7c970b60a721d", x"705497d8736619d8", x"b973ee33f10c18f7", x"b0fd3d21d5e42469");
            when 11761523 => data <= (x"820ea5d1d7bb51d0", x"2432180f39df9d0a", x"f98f37cbc2f6e717", x"8f9ce3483915133c", x"2503d9238acde5bd", x"bbcc826a30116792", x"bf250c013a2ba87f", x"1c81b424256ade27");
            when 19694341 => data <= (x"8513907d0f654435", x"bf2b4237d1e0f3ee", x"6a4ccc0fc63b62e2", x"cf0fd2ca8e375e27", x"685f16b95416fba0", x"a7ee22912f78079e", x"42f0c3279c65f803", x"d68e503039de105b");
            when 28120888 => data <= (x"d3e34912bf84e2f9", x"3e00e37fd529c965", x"554f54384e754840", x"ad0e039d5f73033b", x"5f322d5f769bcb8f", x"aee95df688799dff", x"b5963211630c7774", x"d2ae30fa7f660b31");
            when 4354234 => data <= (x"b666197b9fde637c", x"b62e3ebb378f2e2f", x"9cf5744e9d4efa6f", x"d75c9e1c29ef9ad2", x"b3ccf06fa4ddf8fc", x"1a1004a24eba1ad5", x"c880395f29a88a8f", x"b7a3bf58c872b6d3");
            when 5235316 => data <= (x"2e89869109be58b0", x"0acaee3022827db7", x"b60fb7aa5edbbb2c", x"feb3b72baf9b41a4", x"0c9918cb7878c5e8", x"d5aff700d04fc47b", x"6035c53e59c3fc09", x"d2582a9da92bc803");
            when 3093004 => data <= (x"351efc5ca938552b", x"f59c21f2ad034468", x"f66573d53e4d35d1", x"624c5792ce2a9e05", x"55cbdad24e27a569", x"ef1b174711d3aecc", x"8ffa79c3ba046ccb", x"8500ef57064aa7b6");
            when 2856856 => data <= (x"995f294302dbfe5d", x"de3067b17a2f9b1e", x"c7747b2c18d22337", x"bcd9e833c1621dbe", x"fbe3d9695a96bf64", x"d3558885dbb58796", x"fb0815e1014ed4d1", x"253a018dde120412");
            when 2748945 => data <= (x"522390143c886c38", x"4ab75b58b722913f", x"0586f53ad854b939", x"df69a57c3c0a21b2", x"615de5fbf6c04368", x"4901603399cbc979", x"1d851c9bf474bb6d", x"3f102bbc3f3af51c");
            when 20023672 => data <= (x"89263ede9f45bf19", x"c495efce81394bf0", x"3857a49aacfaabec", x"16c9cd8515b2bb6f", x"526ddc8ea430df45", x"704fd6f508ea4a30", x"64d5004ee280dcfb", x"f65e7e58af765914");
            when 1656836 => data <= (x"60c734e197272bf7", x"ebd80255dc2b4ddf", x"50ed69af65bf7b0f", x"d83a99e8af7c8fec", x"5138e95eddab992c", x"b9aa25d0f4e66705", x"189727ffe1fde4f6", x"324a4e0eb9f26b9c");
            when 3247583 => data <= (x"e11235e42034a032", x"8c24e9fbcb13b814", x"bf8e58ecb286f30a", x"cacabbe97db19682", x"b37022d639c76c8e", x"8bf7cc83debe4bde", x"5e44243d2af2abe4", x"91f3d748e3d27863");
            when 12403074 => data <= (x"c2debea21fae15ef", x"cf5e81f7b750107c", x"aa2a86c9a0757f67", x"80c0b35462a4f259", x"891faa6926088874", x"58dcd4c4044cdff5", x"62edf3d992bf6dc5", x"16f6ab40d4d189ae");
            when 31886189 => data <= (x"f81258bd5c0445a6", x"53f0a2efc08bc244", x"495ea0ef73b918a2", x"5ce56b5cc6044ac5", x"744a0b6ece9de469", x"22027006ae45f7ee", x"1ce872edea65648e", x"9edee802adab71b9");
            when 7274851 => data <= (x"cf57e0c015a112c4", x"ddff6634e37c1e61", x"a1d5a029da15ef03", x"4fd7476d0efd4a19", x"66245391a1640965", x"d917d6ae312563a9", x"314c4770309445be", x"d92e5d1e6d8bde76");
            when 16081620 => data <= (x"b1a7d3fcf111a114", x"24bedf0fadc8579a", x"1c7d54c3a4d7edcf", x"266bfc9cd52591ee", x"5073277ce2579fdf", x"97457b9e0b91918b", x"5f6f476c214f49dd", x"a5e2b37cf36aced8");
            when 15107463 => data <= (x"5ba59f91f8a8824c", x"b30903b949a12e7f", x"ddc2c9c6e0544f24", x"2851560c1ccbb6ed", x"de15499d9967c06b", x"c2204f24c59bcbfe", x"75ecd9af335f56e8", x"cad34a554861618f");
            when 20675149 => data <= (x"66d7b89d688a6e46", x"e3719d9ddb55de94", x"b66ff08728f3ce97", x"3a59a42f39567995", x"80a32dc9cd4696f0", x"2a4e3b5283bd24a9", x"7bd5098148cd56a1", x"06beba774bd72b52");
            when 32416495 => data <= (x"21f78274a008d4bd", x"3f94f229e6e8b037", x"f8c905007cddc3ba", x"445c6f4cb8825b0b", x"5db8d75cee2e9cde", x"02fbb8fe91c063c4", x"36ad7827c1f2fa0e", x"32772a1c85bc46ea");
            when 18237038 => data <= (x"b02d98a5c63f16da", x"5818f87458597f3c", x"a2e63c1d8433b97f", x"accecc6b0138a38e", x"5be8f1fe4c3124d7", x"e3c0959b5ce2a999", x"9155c42addd5ede4", x"14a30cb1fc35e9ac");
            when 14974371 => data <= (x"93fde122d1cc19c6", x"362b9eec3e449773", x"7cca2ed801e9ec9a", x"f8456564f4b0fe32", x"b5a1ef1f0aa4f746", x"5b8d650c9a2494a6", x"1ce13ea2aac639ba", x"7241a7d04d29c059");
            when 4839843 => data <= (x"128f8eacecd04137", x"65a3e61a83112907", x"2693cde2c8a6c01d", x"077309875a367405", x"dfb8e4f318c71911", x"2073d90d60a1ee81", x"5f97216b9008fe76", x"8b754e31e0a57369");
            when 8333901 => data <= (x"1486bd3ec11a0581", x"0484dd68bee093b4", x"826123ae5f181ec1", x"1d809272156c0add", x"6b03494c30a7c5cf", x"f24208803a773bc3", x"7e828dec245cbff3", x"daeebb570dc2138e");
            when 15333266 => data <= (x"15c3fc02328dbfb3", x"93100e7434d3fe9a", x"515c3781b4ce9ecc", x"90150048beb73dbc", x"b5568986193975e4", x"0f8027c028610927", x"efd2f1e0f83d133f", x"646e3c2b17459265");
            when 22769976 => data <= (x"ed707c2fd9146d9a", x"ea5b0cf865069593", x"eb22b87019def9b6", x"804b8cc59a491952", x"ac3c2c88adc430eb", x"7520514c18612811", x"778620ed30418da6", x"0a17b770eed82ef9");
            when 25633074 => data <= (x"4762e03e73d60831", x"ca3d8b1d1cc233e0", x"b9aa1ee6f1266d1d", x"d6e842dc582f2528", x"9054d9fe14f076c5", x"f434135cb1cbd956", x"88757f3a85d197d1", x"7c075cc50f7b8c32");
            when 26894808 => data <= (x"2c7b63f28d3fb48c", x"bb1c5efa4565bb78", x"26a67f7903959fc6", x"ddcbdabf54205877", x"c24cf9062800891d", x"b6a52cde9467930b", x"c152f062e1400015", x"df54ae670ccaa463");
            when 15355945 => data <= (x"a6e5bd7bd2d1882f", x"663b4e56a8586639", x"308db56ca34556d8", x"c25a6d0eb51e4075", x"86ba642f73c94a34", x"f644e74fc5bd408d", x"cee8d41e0e917e05", x"e5396bd28207266b");
            when 32600187 => data <= (x"f740b79db509823a", x"bce496428397c95b", x"9d5d3ba486e887e4", x"3187dfdc11741ea1", x"df87b50ab851b0b8", x"ad38e65b865aee38", x"8ba93ac1d0147421", x"1569bdf6f8ad6acb");
            when 31207856 => data <= (x"9a878cd46041a711", x"daf258371fa6a1ca", x"ab1c3aeb8cc2b70d", x"2b83ccf33c750ab6", x"4ee2fbf3764f7c4b", x"59f33816945f39c2", x"704f88abacc687e7", x"98e0078e768e7116");
            when 32679162 => data <= (x"150f86b284465308", x"1d5fdfe4075b2afd", x"de937f95f2065d6c", x"5f3c68f15ca9f6b8", x"7136bd94c664926d", x"a4b94df7f9562b8b", x"7fcb0cbb42d1a6c3", x"ba0954d7dd315c4f");
            when 1179530 => data <= (x"2a3de406f39c4ec8", x"c60e41d51b14a81d", x"3d6fce270b0480cc", x"4e7a0f63af47ef09", x"9c1be96a9c887d40", x"6149f26dff79dd6a", x"aaeb66f0141ddd99", x"22129fcd8d755e4e");
            when 30343341 => data <= (x"ed2fb92c661a11a1", x"f617e73f8aa12e64", x"bdfbdac276a05496", x"2cdea0cf28d3218c", x"d6bae416002ea46d", x"b9704dc9e2913cdf", x"d25c8d066cce635c", x"c5683e0a8005beee");
            when 24694703 => data <= (x"409ee91c142b01dc", x"2bed308efd60207d", x"647bda751632b766", x"486285c71dc30d10", x"0eac828e9ca4131f", x"0cdfa5f117bb0866", x"e398f95a51d54d3e", x"54cdf2457be320d7");
            when 1080339 => data <= (x"0b3cf3b32f05110d", x"a92cc51551883f5b", x"0f976c19ac3a1bca", x"f22418bf56a52abe", x"7b366746a2e0c411", x"bd0561dbe0e7dfe7", x"0ea7808711a45d91", x"225ba9769650cf08");
            when 5776823 => data <= (x"bb1fab95e4212a48", x"0684d4eb410a3a6f", x"953b055e33f49a3f", x"7bcf0bdcc19aa65b", x"10740ba5d7df7d27", x"e6bc766c5a337b56", x"6fb0ead2cb121d7e", x"5b6da36f6d8ee5a8");
            when 15273475 => data <= (x"d52f702e6eb4e45c", x"21a0b443576c9693", x"cc370ff3d48e1944", x"3a0c8c81cfe449ce", x"c001e46a277a651c", x"d2a18538bd50715e", x"ac6d5807a335b4f0", x"6ebccc0c94d3cd4c");
            when 9400934 => data <= (x"1efac77cbc7e2931", x"03357357fee4b330", x"c08ba9685e99adae", x"0ddf21d4e0876efc", x"7f9b0e9129bf6ad9", x"c554e86f21e6666b", x"e8776ab73e846134", x"38b389369e9d3ca1");
            when 26350262 => data <= (x"755e3f5bd0a6bd52", x"9c52f5c67390a58b", x"f6c3990bc58030ea", x"26d8d8f7e7a93c86", x"d3ca3818b996e7db", x"3233169fa70d6667", x"41a3c9759bc0c79f", x"f2338dbfd6201921");
            when 6599454 => data <= (x"bb3677f56bbd19bd", x"fabff6ef9cac2513", x"5537e73cdfa5e632", x"1b1d3a4ee36dbd06", x"6ece5bef5dd0b561", x"6135e7e6d184323d", x"11d60a8e0d6cb99c", x"d74c5a3ff40faa41");
            when 5165905 => data <= (x"6df20d586c227d9c", x"b3c223ae2a9050a5", x"011f11cc42e84df6", x"bd25ae687073c353", x"5e7b9f321c3c118b", x"ddf514774d310c81", x"500364452c58d31a", x"fdac9a97bf1f478f");
            when 12407203 => data <= (x"9df09d046f04e307", x"c55fcb426c33fedc", x"1cadd3cfc08a9489", x"3676101ab1f4cbfa", x"322644b6ab671997", x"28f5e7a87668c068", x"9d1828757054bd35", x"c886a4e6c5f33015");
            when 32499957 => data <= (x"647b7b82ccaff6af", x"f1f1d2a9d66efe1e", x"377b2282acf53eab", x"d9e0dec9776e72be", x"37233240877ef51c", x"cac1107e48fc1661", x"ba21b1b24ab56042", x"6b74185c86fc6f44");
            when 33307114 => data <= (x"d022178cb5f78f0b", x"11ffa09fc268f171", x"3ce71fead20cabaa", x"fa14c075fb722d5b", x"05bd9046d3798bc7", x"ded93d8f1521bf13", x"06547d33860df34d", x"84add85c5e99c886");
            when 21009907 => data <= (x"fd765103595afc07", x"1525d3f218849c2a", x"5685d67ab4fc4b37", x"8aa1971aa726dc2b", x"5278eec90dcccd16", x"61c222a2a2dc40db", x"208764980c350643", x"e41b99425ae635ef");
            when 31444014 => data <= (x"a42c7361dbdd8657", x"4dc25e47195ca5ab", x"3feeaf46f745bd42", x"d3b546c570975f9a", x"5495125795ff6d82", x"ecb7654dc2d9b055", x"9fd08b099f5fe519", x"27b0ac4c68a35e71");
            when 17599553 => data <= (x"67428d1ddd524828", x"2b3917289fe363e4", x"0c7d347a51f55ed2", x"824441c0cf4c8a51", x"c3f01ac25e259143", x"7ce5daf23157e8e5", x"5e2ee8f840b30a60", x"8382fcd0d60769fa");
            when 3442509 => data <= (x"750c7004cf09ca24", x"080224578645870f", x"817a3a49942fad38", x"b88a2b4bba82e95e", x"f2f6918f72c80238", x"5e5cea5f1bb230f3", x"c5aed5e00b317ff1", x"280cd27bb4464b03");
            when 16788159 => data <= (x"d1704d2c011ecb3b", x"c3fe785a27ea79be", x"616e2684cf06da3d", x"6727c19aa8d34e48", x"1a49657c0d067a54", x"9a7b9838a6ab2ef9", x"5179d46fac533f07", x"5def79fa2ddaacea");
            when 33061819 => data <= (x"8ef6dc2e45219478", x"68136b3d2be6d599", x"6f3074ae78a909c4", x"05bb4e39d7f03cd5", x"cd9183ebc80a503f", x"e3f51348cee6f738", x"be7f33d6da6affbc", x"a1458e51323015ea");
            when 26706417 => data <= (x"9e4eb08d62519609", x"bf3afa05c8a2fd02", x"33918536b7297477", x"f33518a9f2a5ce5c", x"2fd06e8f7c31fcd0", x"819286562f6001c0", x"877b33e314d4d8c1", x"6b34919248e75222");
            when 986337 => data <= (x"c15a45bcb0d3177b", x"79c09a5efd5b1950", x"a725a84850a3c4ec", x"34a307755034bd24", x"4e263a141f734b93", x"c9e138b013ebddcd", x"cecb162d7f1b689f", x"cbba704aa9db1655");
            when 5810739 => data <= (x"511fd828648ff400", x"cd7c5507f63a4883", x"683db81f28a97925", x"3c5764c56979fabd", x"a4e02a62a97e04a6", x"832a20593e7e15fe", x"fb7b7b4d488f7914", x"c6e915dc8cdab2a9");
            when 9853993 => data <= (x"ce36dbdb5638a030", x"3205119d358be9b9", x"686c883c79187576", x"7b254c5793a4cbd3", x"44db2550b1a7a690", x"b82a80b02691f911", x"15cee4fac197915a", x"d4fd9dbc520f6673");
            when 28113625 => data <= (x"6a70fd2ccb21cc29", x"c94677e8b26f2fc1", x"802eaccad7350f65", x"e9f280bfe698c335", x"9b451e411b51a62d", x"3a93e2ed08413ded", x"be771bf14493c961", x"a3872589f3d10159");
            when 8161206 => data <= (x"0487536557fe7ea3", x"eed740fd7729ddb9", x"0beffe5734cd42d4", x"e6cc83556722edb5", x"8dc453023732d218", x"818a9b6c88075a93", x"4dfd1e38b4de4c79", x"2d16b95b4e53895b");
            when 15304481 => data <= (x"96a70449005ec91c", x"cbe9781958c6dd69", x"a59ea496c10f24fb", x"281ebbdc9008141a", x"94cbd93e2de06096", x"6d4301d641f7539a", x"6f9581603434e290", x"ebd823913e6f8b51");
            when 10080880 => data <= (x"c509427a993db7ed", x"f7daad435a0338b2", x"fc3c1260dc4aaf25", x"eb5d650bbe43c8f5", x"5e8540ecad67dccd", x"d61c35aac00d2a44", x"e139483cf2ba7396", x"e7ef278087d875c7");
            when 3104734 => data <= (x"6af857aaf7f7e940", x"76f6895d252214e7", x"266050185eb1b8fd", x"2b61eff11a12a309", x"e94970b19986fe04", x"deda1cbf9c2862f4", x"8df8207af87f9262", x"0c0fd538f79c36ea");
            when 21782456 => data <= (x"82c345ad160adfa3", x"028305733db9c405", x"fc8f55af96914d47", x"c94f12b595bcfe0c", x"13490aa6f53b36a8", x"1cec479686974968", x"dd25b693122f0d29", x"7df689206bdb5e15");
            when 5564091 => data <= (x"295a84e63493f085", x"984562ce2ff6dfdf", x"f95b32e6ee001bbd", x"50971cc33634eb59", x"6d7443f360954ae1", x"d5ba272f37c20799", x"734727f543944a9d", x"78427dfdd70b3ccb");
            when 21055497 => data <= (x"c76bd3ed395c4b51", x"c9a86c49599efc77", x"7292c7a56f5b065f", x"832f8167a48b15de", x"bc44edc8d2e3aeb6", x"c757b2001260054f", x"fca23c4e7496708f", x"596e4c13cc260056");
            when 19652113 => data <= (x"6dc50470f84d494d", x"42d843ed89a453c4", x"840cd520f46da4a4", x"8956076d030a6c59", x"74019afa25dc0a23", x"2ebbd945ff7396b4", x"2f41be18a32d54fa", x"3f3e425ec7376c87");
            when 10229857 => data <= (x"c47c2a4aa743b9ee", x"d474dc6d1128eed4", x"7cbb648c4941e0ac", x"18a1db4d64f12eaa", x"d6ff8d45c8782106", x"18950e75a4db741e", x"c9413f22ad0a8e6f", x"878729cbf9f44c50");
            when 20501018 => data <= (x"d6671f8e36089f7a", x"565b438ec70cd29f", x"8bc387db6dcf8288", x"8ee8413944c15bc0", x"81078f22720d7986", x"00e1e3c7dc1b059a", x"4cf7779ff9e4a241", x"96842c722272e59f");
            when 1506004 => data <= (x"ab5e417f3828b1b1", x"8f83e1ac179cf1af", x"ed19e7c141632fb3", x"bb9073dfe6cb08dc", x"56e66908c83c2b54", x"21220ee7c2cd5ece", x"0aa546dee32648cf", x"33591a410cf089f0");
            when 14139331 => data <= (x"8acf5e45a2c349e8", x"cbeee45b5dfbcaf1", x"0e6a92156a448dec", x"ed6edf3af7928966", x"a9142595e560fed4", x"db1dc6cdf11626af", x"52ccd9957c5f3e07", x"08f2dcc6f4f86dd9");
            when 26751651 => data <= (x"910e7b94918ec2bd", x"05baa00cd721e9cd", x"c89a4e14471c7cbe", x"0baa5592077aff23", x"aa5d1803226ab50f", x"f78ae36d381d1abc", x"9233dde7e4f3a48b", x"367cd7967b3dd9a3");
            when 343437 => data <= (x"557b05fd0015d1ae", x"cd74356927d76a7c", x"f93007bfd229a0a2", x"794ecb603ccbf27e", x"f8b69afec7cad83a", x"248664656a2b80d4", x"32dc7db4cda49559", x"77ac8df4c35af91a");
            when 17569353 => data <= (x"abf627e7ff9d8d86", x"a6dd1fb1625ceeec", x"4827f50eca7ccb43", x"8ab8ab80c053f4cf", x"002172dd0ce7bf1f", x"fdcf334f9c25cdd5", x"ed7dbb72af15845a", x"1fbf52946ae2bff0");
            when 26721718 => data <= (x"162086df7b4024b3", x"e08b28a259f7bf81", x"78d5500ca172040b", x"555b794ced95368b", x"49d01acb9f1120ab", x"fa71b753c952b484", x"fe3bf87f8d5f98a3", x"1530150d7905dfc3");
            when 6923260 => data <= (x"f9014b3f2c93f613", x"d279507d388b50ac", x"8d242237a015d991", x"49f59e4f81e66ac5", x"4716c8e2ca50928a", x"217e464d0e394c14", x"250e2bf36cf45517", x"9e77aa2eea5ab5a8");
            when 10406034 => data <= (x"75d397e6ac1d8d0b", x"21059a8228cf70b5", x"cb0892dba149dff1", x"02cfccdcf20fc195", x"c475144eb9a0a7cb", x"cf7e9f0ac485a584", x"f26c99845a5848ef", x"723422fadbf5d5e9");
            when 28358148 => data <= (x"4e2bd055dd231c25", x"15f621529cc22f39", x"96a94bee4d9f3801", x"b59eeed4b2b7d3a4", x"c3d455166d9dba55", x"28e25e6b1b5c7522", x"511fc41b7f8f92b8", x"eee697c1b66ce852");
            when 5442007 => data <= (x"afd84a5ab7ed650f", x"5396183483c3775f", x"ada413dba7baaed7", x"109a506f4a0a6f12", x"2ee2956b1cdf5642", x"ac64b59a4916f969", x"b9cc88681c459d42", x"7eb9aa42bc217231");
            when 7724488 => data <= (x"a22ada08901ce97b", x"a659e164aae14370", x"1b60c058df2a9adb", x"a2c81a7a04aa7a9a", x"65a335185be3593b", x"e5229aaedc2172d5", x"322e0c6788311b76", x"ce39fdd40dbeb56a");
            when 18423261 => data <= (x"60dff0935c8842e4", x"090f0d73c6962df7", x"43092de43f4adb05", x"2f9a7dc3230e04cb", x"0d8b0c0a02db1675", x"cd21de403a0f2c1b", x"afdf18732b137622", x"1812a3fde0e4884a");
            when 22188898 => data <= (x"31c8787b18f8b06f", x"cc85e86f49739241", x"3abde1d4b5e5a830", x"7a5a34f04b08766b", x"2104561cde0ddc67", x"5feb59fcb32c9adf", x"69bfd4d462203de8", x"abd6d869ffb3e1f9");
            when 7063583 => data <= (x"6e29c27517789050", x"0bc2c66aceb3fbc1", x"be580732375d4baa", x"4b0f95127c6119cc", x"1f5a41b2c56d923b", x"498c4d20e299a1cc", x"25945bf2249dde56", x"80e6be28718f5b2f");
            when 2022859 => data <= (x"0913f5c800675f7f", x"b8103b0c769d55de", x"f4d8ea570f583b31", x"eed2858e822723a2", x"d079311f76601f95", x"b14c1f8369e3b8ec", x"1fd3610a8ddeff09", x"26fb7e0d95a8c492");
            when 25094561 => data <= (x"cbda5f6f05cf4445", x"d9007a66f6c97fd7", x"14361703ee3632ea", x"4325035efc0f3b7e", x"5a2f41ad00dfef64", x"c924a899b6b7688a", x"91b521b172c5a5b6", x"fa8776716c21d0bc");
            when 25827381 => data <= (x"8d27ad58ac01c938", x"873a121eb157ebdd", x"fdfedd0e1179381c", x"2fbe2955aa385dc2", x"dbde83b9c50ef0bd", x"83535630edb82dcd", x"ad3479fafea271b3", x"29121aa5931e86fd");
            when 7623047 => data <= (x"877982f2bebdfbc4", x"06fcc36241b69a4f", x"86f58ee6ad43005b", x"e46e8fdf78f45261", x"aafc3ba4c5facd4a", x"d5fc63721e828da4", x"5b6f8bf273cedbac", x"2e8279665df609a0");
            when 2713374 => data <= (x"68323a7bd4c774bb", x"ed053c32a75a223d", x"9c1ecca9a22095a0", x"a27f6d5c5c5bbec3", x"1f726b24650dc47f", x"2942e58305f0edae", x"36db3e2af0829796", x"774dc101c124f487");
            when 21571308 => data <= (x"3c865a106d08ea74", x"6ec581530739db57", x"f4b7147598ecd1a9", x"e47f53d0cde5de7b", x"62682137def0169a", x"11f21ba664568aa9", x"cbc450c67ab14071", x"7a0c84091b2db211");
            when 14343069 => data <= (x"e1f6f81c779c7f85", x"36c7895cda56f3e2", x"d0cd61c2acf6394b", x"53c4e77e1245c8e7", x"d1526a7d4b89112b", x"490ee35aea713a32", x"9aa3d55bed9b7a6c", x"c0d47e63307b2b56");
            when 25419342 => data <= (x"ad0801d992e7cf1f", x"a552832dc239d4b5", x"a410c71b1325888e", x"f17e126e41c73144", x"0dcafe60b86d11d1", x"380f82ade8a471a8", x"85adf56246be03ad", x"4b3abe65b1271568");
            when 16487877 => data <= (x"dde9f5b3157064ef", x"a815bfb516f3c0fd", x"1920675da45f95fc", x"15584688c23e3112", x"40bf48707bc39464", x"9e2b026b7f7cd204", x"a75df697654101bd", x"efa2b9bf1e73ae22");
            when 1366643 => data <= (x"8c3c74e22eace380", x"72a2dedabaccf5ae", x"39db2e2fc5d4c545", x"3d61d8ca7cace96f", x"554f8f9f9a324c95", x"409c00ad8e3d3a5e", x"97cee7a9e11063ee", x"21358add939403f4");
            when 8129482 => data <= (x"d943f1a93d9bc0ee", x"63c8846747b96296", x"b394ebe69de6e506", x"2cdaafb8c27bd33f", x"cfb31442ccf5534b", x"d0331e37c9cb1e22", x"c9b3c25da86380dc", x"22d9c634503c60c9");
            when 19505302 => data <= (x"bb7ce0363f9c52f9", x"47c942564285edd3", x"7664ec35f8e6375a", x"d896b2bdce3bb781", x"756204e83bb7a349", x"6241dc42fd27543d", x"05709eeb775ead7e", x"11772aba6c355cea");
            when 17600520 => data <= (x"b2c2a9d5122508c5", x"330e58eb2b16a211", x"001a45fb2ee66d28", x"8c150abafd4cfd8a", x"c6d99c0bc70535ad", x"f97012819d539a6d", x"037394b9d58d4215", x"54d3b37e8c49fd25");
            when 18076439 => data <= (x"ae5efd1a004b604e", x"d6311fa2c32018e3", x"c2c69b4cbad22a30", x"03169d1da5c45186", x"4fd17bb32e2f81d0", x"cc12f1afbe32e0df", x"ff0e3881968af151", x"c0b137e0b0a5f747");
            when 20050755 => data <= (x"e4c801bb84ce978d", x"991e4b00d3e5c9cb", x"867f731acc8648d0", x"04acbb99989641b7", x"f9c4a295722ae1ab", x"5229055a30b6cb6c", x"6e4a0cc75634c105", x"ed6e20742ef1404e");
            when 28300136 => data <= (x"e2f16a1926a9da3e", x"9e4cbb98f0f33487", x"6eb8710c6249e588", x"354894bb822a97ac", x"0c46994b753b97d7", x"a7e1359cde4b548d", x"db051872d6256649", x"7039d7f4102c971b");
            when 20163070 => data <= (x"40bec7b5bd58bded", x"0604489b3523e4c4", x"82eb3e10e7c71f19", x"4dafd96a0ea711aa", x"c8dd49d8bdcdb3f4", x"e9f8382b4a3df2eb", x"c2512ea8d1f3dcf2", x"6a10069a8cd4792d");
            when 10916466 => data <= (x"061c73a6ff0af74b", x"fb5aaa0cf6b195e7", x"d1c9a366b473d270", x"566884846d9d2674", x"ed14aa88c4031798", x"9a473da643dd9eda", x"5d507684e0d20485", x"580d71ffd978ff43");
            when 21245529 => data <= (x"6fd25f14ed4b50f7", x"e15ae2f647696017", x"641b123c60a4d226", x"190c6c5be381cdea", x"43757f5eaa212920", x"8b89d00b6d27c3c2", x"fa5e46aada1e83c4", x"3fea2886f2623ce3");
            when 7898999 => data <= (x"aa7dc39c2acf80c9", x"7e596f0ce8ddf7e6", x"16559789bd94d2d1", x"68af3b6d399834d6", x"102ccbd9b5c1381e", x"8f0c99c38d210eef", x"3c1a222a47476940", x"0bd9637cb32bd8c8");
            when 22056439 => data <= (x"b25e3dd62ebf0d82", x"725d0fa6358816f6", x"b67ef429440b0539", x"196b011b04103c38", x"a405394d51b8aa96", x"59231999a32977a6", x"d7d5925ad751ebae", x"71a50d3228fe1c74");
            when 8644947 => data <= (x"d3418832d4c7c02f", x"57b75d14012500c7", x"7a9af67cb9422d4b", x"b3769744d2b805b3", x"d3cc9bb7c6ed2a61", x"134632dbe42b644e", x"760bc348e33d2ab1", x"540c0028e372da25");
            when 25528903 => data <= (x"6aba83af0d0d9da2", x"6a2a232dfc150ec2", x"b7d39009d959bdc2", x"0a46a302f459dd15", x"01c986211714b2e6", x"0f12656e8aefefa2", x"833736d202b5e7b5", x"282325f3c0e143e2");
            when 1124096 => data <= (x"167459dbbef861fd", x"49afbd2c74a032fc", x"a2402d0ce9b4f5a0", x"2a36ea3d79746375", x"9e096928bee7d4b4", x"2846a49c400cdb8f", x"2e06ecfea2bc8c13", x"87f3542cf9258d0b");
            when 29088922 => data <= (x"972e27104b0b503e", x"9f905df5280e0dc3", x"6a28ed24c50bd250", x"9271b69ffcf805dd", x"deb1ef321904fa37", x"04e14249f62b07d7", x"63905af6162cdd38", x"6714b5f2b1ad7517");
            when 903064 => data <= (x"f331c3769daa5fdd", x"68f08ef964d515ed", x"0522ea84fa360837", x"500ab1ba156387d9", x"528091b14cb553b2", x"adef43af482d2e50", x"074e67f59469f318", x"36bee07c75893018");
            when 20469463 => data <= (x"59d6b6e451827f59", x"c83b61984542d83b", x"aa3518594fcd132d", x"4e4347b8f8a55c7a", x"2b1dd01a6f7a862d", x"f252272591e9c9e1", x"ae3b45026d74be09", x"d026d6313a62d854");
            when 15655464 => data <= (x"69df8349df753ce4", x"366fedfdcd96d990", x"a4570313c5f6cf55", x"9ae4bfe2be56d2fc", x"d4ea3b8ab3c6ed04", x"0f1e8bb49b76b28d", x"333e7d2ef01be0ae", x"bf399de827a5b999");
            when 8317472 => data <= (x"6b0cd313d065d5fc", x"ba4455818f642910", x"e8782dbcdf57218f", x"7a061481452b1aaf", x"a7af54cb8504b6ad", x"96aa03cdb17a9f21", x"4e36a89a622c7d8d", x"41cc5bfe0be47907");
            when 12343525 => data <= (x"d709689b51b73391", x"42b577badce67875", x"25d0bc762e524267", x"8cf39f25a5744376", x"0935ad83dbe7b67a", x"f9ecc66b076c5355", x"f3caf1eb006dd077", x"737f03a89e6b3cb9");
            when 1762825 => data <= (x"e45a0627bbbe2dd3", x"b2d6ceed526e5f37", x"44613301f051e63b", x"3142ce475cad3986", x"8457ba65d42b7877", x"f328d6ff17ad87ad", x"064041544c5b487e", x"39bcec3bf6ad2d32");
            when 31577695 => data <= (x"2fa245a9ba1567a6", x"dc698bb92938b8c9", x"ce0018516ecb5404", x"6932d9e0e438410b", x"f2ed348531a2c0c8", x"03e00cc4d513877d", x"4250599572c3642c", x"54c196447b1a567a");
            when 11216570 => data <= (x"7f1c72e66bbf0d1b", x"01e3aa618e99fb72", x"e6cbff44914bb385", x"589acab7b414d778", x"98613805dc1f5e1b", x"c6b4b5d93669adea", x"bac45081e73fa614", x"6db569d38d86083b");
            when 19392038 => data <= (x"661b21f8ca94a5d3", x"0adf00add1f0067d", x"c6cdc2a2361d527d", x"3a5009cf6cbf01bf", x"d5d114e62b2004bd", x"9acce2219559c7ff", x"dbb919f1e23d3304", x"85d9db89defcffad");
            when 23775941 => data <= (x"97f9191c906fa5cb", x"ea4f2ccce41f0a3b", x"086342c0462d761b", x"5701292593dd6e64", x"52d6ca16624b1cd9", x"8db2a4b7af80ddf8", x"ab5df8b3230d95ab", x"2cba324431fa853d");
            when 870239 => data <= (x"0430951b706aba77", x"84479d481ebf8ffe", x"600144cf358124cb", x"1829c441dbdb9228", x"64ae0b77ec8bae8d", x"af9c75d8e151b729", x"71bc19b4a95f6a1f", x"e4e5a01dc7776b99");
            when 33468284 => data <= (x"b25322afe10966e5", x"491ba924af19df04", x"24379b699e386fc1", x"79ed43b5fb577738", x"9bf02ea9fec03004", x"87719d2031ea051b", x"6a4dd13a9c69cd31", x"1e283014a9fa4112");
            when 24308574 => data <= (x"ec247fc74bb91a0c", x"8f66dd7300b08576", x"e54ba1d6536f156b", x"3a14bed74ccdabb0", x"47cf2799a6ec745d", x"4502357f645f3397", x"32788b52b434df89", x"de21079b55105909");
            when 3425723 => data <= (x"b515680312b463b2", x"9c62b15cd860cb66", x"20dc96e660e5a2a0", x"1cc9ed259018956a", x"6a55b196d0b09429", x"253d43a3a8c39dfd", x"591ac834f971be0b", x"787c600a280bad42");
            when 15209554 => data <= (x"3401f7f0ea3f0e7b", x"c2f0f5808bf5c6f4", x"7491f1ddf0258a5a", x"01d80c88d95e3f78", x"8e5e68f7d4b1fcbe", x"7e21ffa72b0746dd", x"f592f54a65530583", x"c7b39b9c9d2eca3c");
            when 8606070 => data <= (x"21a0794b47c986ee", x"9f1a2095a15d05ff", x"2b0de257d3b43132", x"7f8c7d6a440e50fe", x"d4e5a379f547bcdc", x"f98de1603dde480e", x"e1ec257022ee322e", x"cc607674d30ad413");
            when 15170486 => data <= (x"a7bc71dafffa8860", x"555cc89b89d14424", x"1618af1ccd583b9e", x"dc78dd16412b2608", x"f4e7fa8b3386ad06", x"7a7bf8f2b4833fcb", x"4234a86ba3f08daa", x"314bc919a31d9eb1");
            when 33265540 => data <= (x"fd17d15d07875847", x"daeb5a166fde6cff", x"f24f7540651b76c3", x"6a43fe6f282d1259", x"3624832074ce86df", x"01091a6c78d44edc", x"b6188a930879d243", x"e67c3a1e974b2a03");
            when 2942930 => data <= (x"c2a98fd57f616bc1", x"af6e53fb8bf4c86b", x"03f3118d521f7bdf", x"3ab4a81a781c2cb6", x"0973d68d25b21efe", x"63d34be9a021c2b5", x"dfe9d672a7a982cf", x"a510a284cbeb8476");
            when 31627743 => data <= (x"a342f5b5bc5a0a06", x"13ef161c5bb246d9", x"520e5adfc423a7c2", x"815f53884575900a", x"06c8b8fab0f8ba01", x"73bb150810143e1e", x"2db0e2a82d4211f8", x"9669405770ae8b5c");
            when 16486997 => data <= (x"59b027fbd1a4a89b", x"790b1567cf8bc027", x"cad9a0b26721ee4a", x"9be0820bca9444d0", x"e43deccd86b980c7", x"aea1abfba77d1d5b", x"62ae75ce825fa6c0", x"7b6be56ae93cfa21");
            when 30641991 => data <= (x"59e3d1f1dcdfc306", x"b37df7144c7061f2", x"b435268eda337737", x"bd1224a4430f82a5", x"31a7904079c93db7", x"543159030e842ba7", x"5eb588d42d12a330", x"4329e4ef72f1c6f8");
            when 6391867 => data <= (x"4ef4c542ef984b75", x"9de36120639d587e", x"87d4b13e23757611", x"7ccbf652c730d8ae", x"b8e985870285d7c7", x"df38c9f71757551f", x"8aee641f5553a7fa", x"451aa89972fd258c");
            when 12785599 => data <= (x"c693ed813e8c1bde", x"0c4ba6d540a7a2c9", x"d9b59ed4ea89f1c4", x"68940b74c793d322", x"7a349bd4fa71f70a", x"c20a07c000927cea", x"71b7e8481b35387c", x"378e5a61888fac1a");
            when 16705492 => data <= (x"b3293b86f92d319c", x"9399b40bb623b68e", x"38916dd49a30fac0", x"aca3e1e77b7b5691", x"63fbc14fbe46a3f0", x"f8fc35f8d6f9cb43", x"7dada7dc1426a7f7", x"17e447efe5175734");
            when 27029030 => data <= (x"42a0aac6630c1400", x"b4955f877393af5e", x"7922b1d0cd781fc1", x"0b0b187a850add29", x"f3557b75c793a0e9", x"daebc0fa134b2090", x"9d01c1958e2dc1a8", x"2d3b000f571581ff");
            when 2299688 => data <= (x"72071bc5a6fa2f22", x"afbf0923f6d3d038", x"ab00e5147cd7d6c7", x"ebbb7c5912e1739c", x"5837e17c42830411", x"60581c3948d7516f", x"aeca7c2e3e0267de", x"85608ec8ccc16801");
            when 1707305 => data <= (x"00f807a61e74bcef", x"16495e264d9c7a57", x"e2f21d2dad20d172", x"3caae2cbd807b2fe", x"4ba9c502ed0416c8", x"41fb929d3018213e", x"e1e061906523c4e9", x"3b04d3b118e47d8e");
            when 674861 => data <= (x"2eedd9f3534c3976", x"bcabe6ca3f193751", x"38839e8707d6ee94", x"62ded2168e0f465c", x"fdd512a67e4f5bca", x"29269c6c84ef1a7e", x"f8ce10537dc10c80", x"7975243e8fca9510");
            when 5898615 => data <= (x"122b8aa819effe82", x"6106cb4b0b9357cd", x"a804b9f12fe144d2", x"2fc493db4a72efb8", x"882f9fd3d9e0d9ae", x"25faecb7ccda5e8f", x"284de4c1eb0d8a42", x"55e8ed651830dd59");
            when 11175724 => data <= (x"48ed85f986bde304", x"1750ffcda2c8161c", x"47ecf2e133232ab6", x"57d875e99cdf4143", x"1d1a8f817aebc7a7", x"e80c986f17c81fa3", x"f3e3ca39fdf5fa3b", x"172a9ddac1ed006b");
            when 20917972 => data <= (x"bb9039616457829e", x"8cd80133618d81dc", x"cbb7eea07bfaabe0", x"7f1c90b6882ccc10", x"ad40a7c4144179f8", x"29c2802f57230ad5", x"81805d7bf2e95b9f", x"77ba70a0e6d0f714");
            when 12241068 => data <= (x"b51dcbb75c7eefdd", x"89e76a51277fe1ef", x"dfd6b63bd2f168d9", x"f7d57ca8bf56c190", x"8bc8cafae1f406b3", x"e744560faf91be7c", x"9708e8a2998afcdf", x"6c94418575a83629");
            when 20016482 => data <= (x"d445f18d1137e92f", x"f177fd3aede8951e", x"291a13d1e1dd8e27", x"1c4726dde3752cb1", x"5f3c0c67603e42d3", x"5a5dd7c12d570e59", x"897b8d15b7e45f33", x"58728fa747b9ad94");
            when 29549419 => data <= (x"f588cc60537ff906", x"a2133c4ea452281e", x"69fb4a49ac09f255", x"d7d926ba180ee10c", x"132e7bda8711d6e6", x"6f7fed1eeef45782", x"71e64c301e744232", x"f7c787c7f1226cba");
            when 11569642 => data <= (x"fe54d10adc7ad045", x"e734cf2fbc53f6b0", x"944225db92c06aba", x"1241432e747e6a47", x"87cbb8c756a16041", x"20128b076f306ef8", x"f53d910957f2da5a", x"00d08c12ccdc061b");
            when 26501313 => data <= (x"ddb420a2cb133d5b", x"f4d5c662bcd6813b", x"20578f8743428732", x"e399b144b5763efb", x"856d0550980e47fa", x"67ac5f1b726f357f", x"ed1554251dec36a8", x"c5f6004b6e02967b");
            when 11971185 => data <= (x"a9257fedfe9d4111", x"3947e3b3a81b0b58", x"4b5b7e74ac091d89", x"6e7b7adff8fa62ba", x"3f193f56a5765217", x"372604f9fea22f57", x"a171751d8d3feafb", x"aa98c7ac1aca9c7b");
            when 18707686 => data <= (x"3ac9c63b85e31344", x"736401f3ea1a88d3", x"92b0b5668bd9e12f", x"544573896de3ee36", x"001b9505cb624b65", x"ed358e60027d4c0d", x"4b57bb873da58bd3", x"5dbf3f6e54d50a66");
            when 19749136 => data <= (x"bede6ff1080a1a30", x"70666d9531008845", x"2be941c0cfc2ebc8", x"64079561b77beb3a", x"f26af923bea20948", x"a5d4e4aac4be02a8", x"e46c1c63dec33e36", x"ff00832b801b5eea");
            when 5322402 => data <= (x"b57e64632afc1649", x"cb027f21ec7b7fad", x"8fdcddd8e2cc1951", x"43c96fcdf63df666", x"849ce1327c49207a", x"95926d553771bafc", x"2553604b616de1db", x"76021a83e3336dba");
            when 29584862 => data <= (x"afe23d4bfcce8c13", x"b4928bdaa8c9e499", x"c2d8ac8375e6f8d3", x"047a8a6ed3a09f7c", x"d9ab55baa3d41dd8", x"8a496d3cf0f0e2d5", x"8e0d4853efec9d71", x"a751d060bbf4ad24");
            when 23838894 => data <= (x"82a97b00ee2b7d0e", x"7b3254629a58c6ee", x"95bcbb83d7b3aa2a", x"f69f96e9925e5a23", x"78e330024eeb244a", x"d116e849fcceb08f", x"ea5335937c475468", x"c563341bc54622d0");
            when 31315619 => data <= (x"5bd37c585743f6bc", x"58972af957c0ee5c", x"cba128ce8d92d7b0", x"54f4237fa9f230b4", x"6092394a7d386d60", x"1ef341b330f0956d", x"08693eace09a40c8", x"2ef6986d2304952e");
            when 12087565 => data <= (x"da0694b62c688721", x"2cda9860aed4f697", x"8fda4606278ddd20", x"9fe1ad60ecb4a548", x"315e53e4238243b0", x"2acef15b05d2ec3a", x"4c1696fc9d3bb90a", x"d5099bbea8d2b46f");
            when 4777750 => data <= (x"ddec1ea3ad16ed55", x"44c8ad6db0fccd5f", x"0ab54c7895a5aa0a", x"ec84c770610759a8", x"dc6f207652788b18", x"70fcaa654aba848b", x"9565e0b8c5bf73bc", x"fb910ca0dccfe6b9");
            when 1778977 => data <= (x"4b9bb3ff507e03d9", x"f44851045f67cf78", x"b6a495af90a67985", x"504337f5cdd79d87", x"31ea8492c4f34110", x"e9c6f4e6bdfc88fb", x"ce2015167f95d880", x"cedef2b19f4d53ae");
            when 28471732 => data <= (x"27b575949e91ba60", x"6d118bff6f9e79b2", x"08accb5b6e6866c6", x"0490059b18b4f463", x"242dd5b3a33ced16", x"da66fadaa42a450f", x"eb9e952fb673848e", x"732ca5f721b8ec57");
            when 29462224 => data <= (x"f0fe31b4921863d3", x"b3b2c8f6071480bf", x"66377378904b1eb0", x"db605e649e9d9a2e", x"f4436ac6bb7ebf7d", x"792c3da01b6a9f99", x"5299bd24769d0f01", x"5274f10a3059ec07");
            when 9511150 => data <= (x"88b37e555eedf2d1", x"f25ca5d689ba804d", x"e0efd31ee75593f8", x"91850bf5d46b83f6", x"2fdf0e15493488c3", x"3ab84b8f18561f1f", x"99a8ae8a839d17fb", x"58d45fc98e70795e");
            when 9943372 => data <= (x"73d60b4c9e4b2514", x"e7667c3b67832725", x"b874dbfddbfdfe8e", x"5bdaadfe7bb625f3", x"8106d95b5cf0c32a", x"79fb518e3a0af44f", x"cd12f842283d13ad", x"e2f272f7c9b12b32");
            when 24119559 => data <= (x"5c068ece6cf6cfec", x"40b11124a9ab9fbc", x"6f2278e5a5958956", x"78cc51eed55ec106", x"c1529a2615774d96", x"bd9fd86f98c91ad4", x"6b153ec49304b02e", x"df1db7bdd1397c7e");
            when 20960565 => data <= (x"720031979e2b9c7a", x"91125e12e079736d", x"2e1428ba05fa79e5", x"12187497643dc815", x"b75b47092ef672b6", x"959294e25e550b3d", x"97d30655d477dd54", x"8055e48668036eb7");
            when 13243299 => data <= (x"6ba21ca6a8fa13a6", x"638d2d4ad7b0bfa8", x"193b267a2a060264", x"1ab0bfc942d5fadb", x"5a28c1d72b40e31b", x"61f9fe7130f0059e", x"1181cb41b356bdb4", x"4c31fa436c81a3c3");
            when 20312224 => data <= (x"e99ce3db48e9fb54", x"2674881631cb9f22", x"7fdfcf40c9d25215", x"7dc9aebcc55508c3", x"3437be37ae2edc42", x"40d98c39df1e50d8", x"ae624a1ceb52d710", x"b9b1cb9e723fef35");
            when 27090501 => data <= (x"1e546a1e5c172a68", x"2ac45622eb9e92f1", x"56543e79f103b9b3", x"157bad3a83649c79", x"3f24af325aca060f", x"92a301ed45977541", x"2118f2e51b75950d", x"3796ad6435022429");
            when 33287959 => data <= (x"a324e77e0c065cd3", x"90f6a7ef8386ec1c", x"b772a8791e0766b1", x"f0e023eda09827ac", x"b81cfe860b43a1c6", x"8082411de2795c47", x"0fe9f181adcecb97", x"ecafeac46667218a");
            when 23140319 => data <= (x"6bb7dcdfd9141a39", x"b13aa8d1748b3f35", x"05d7ce57c99e34b3", x"5dfd5c009c8959e0", x"bae7ac2071c22ac2", x"26f45e92a96ea94a", x"331b5a8d4e630463", x"0136e1ddb448f77d");
            when 9384539 => data <= (x"8d8906c696669932", x"6dfe95630452ae6c", x"565960873ee0e1c9", x"d5972641c1ff443b", x"f5dfe45ff7e33bc3", x"21d1628613fa4002", x"1f6b9cb12339eaf9", x"6d2b13386c106642");
            when 32053144 => data <= (x"81c7dc587e88c754", x"d7266e5047ce41fa", x"4cc26c28314c2465", x"226a1485cd56a6d5", x"feaa35aa2b0b31fb", x"2372e7ded1083def", x"2e7d330fe694464c", x"0367c9ba567ca118");
            when 33341103 => data <= (x"bfc6a2cafcca2905", x"576b630ebb980c0c", x"93fe44dd40aecaad", x"6d3a8d1dd553b18b", x"37c3948f99c91c06", x"c9b2160c98dd2fab", x"d305c0b507898b02", x"52fa40c0984ce334");
            when 5290192 => data <= (x"e1b2c17c2598c13f", x"f9f21e8630434467", x"e7be4c60843f1b49", x"dae678fc24ea0fb4", x"f07d71d533ebb60e", x"6dc474af78c75098", x"5761ffa613c7081b", x"451c27a49ecb0a17");
            when 3961446 => data <= (x"7749d249c9498a72", x"1e46f2491f369484", x"e0f2649b82b4fbdf", x"b85240cb9ff3c3ec", x"dee9de1efe2c039a", x"e2c79b9ab415d2e8", x"27c1ef0ce8d9a007", x"fc72d4d4b40b0bd4");
            when 13572486 => data <= (x"ebba97c75b50cbf8", x"a5791a0a2f3005ec", x"468b046f982a3ba7", x"11a3cb40bfdc4c24", x"74ebda1378482571", x"19346be7bfbba6fd", x"f04d2b25f4471318", x"10636f3383124e16");
            when 29503509 => data <= (x"da32f2adfcf160df", x"5583a4ecdb04ac18", x"a5cfd2d243988332", x"eafdc38f54f428fc", x"5c746b35b2383990", x"ab89eeefc918e175", x"4f61abaf9b6c2db2", x"594721030b36f433");
            when 19746771 => data <= (x"a48094566d9b7a75", x"fd8e5272b58ae8ae", x"d86a1698f1d3d699", x"117a59e53273dd30", x"81780e537622641d", x"f37276eb68dd4aca", x"6498d924aa656571", x"38c7b26010bfbdcb");
            when 2924768 => data <= (x"49830bbb045b2ba0", x"59821aaa56e14523", x"f4a287ca614b857e", x"babd7e3aa8d7e231", x"8f1e486a2dce407a", x"667a067118fe1ba0", x"9d16e294917d81a7", x"f9abe9796c6032a9");
            when 2172746 => data <= (x"8725ee4e7e5472d8", x"00adecda35e87b3d", x"d01d4c2980e38b5f", x"95f92a0cdf8f437f", x"4721969eb02df022", x"345c07727907a869", x"af3840ccf6b7cbfa", x"827912181921e318");
            when 33649304 => data <= (x"d4c45043d91ca6b0", x"2211e670acf8eb08", x"597e8b643bb26728", x"bd42e300a05cfafe", x"2a01edaa4f63e90b", x"20688951fad35c6a", x"c3a191a271fdcf82", x"7b918451280b93b8");
            when 9546195 => data <= (x"4b1fb22272e6ac7f", x"da2db7c15c0f9b64", x"b5dc21bb3d0c5e09", x"6be40b0f31b36e56", x"7568edd6ed1899c0", x"cc485c72e6034354", x"4efd83c3416a24bb", x"e951e754a8083471");
            when 21110232 => data <= (x"6029f2ad2a2e67a3", x"cad155bee197f16c", x"a76b5cf1fbb3b4ed", x"e4aa0fab0590ab86", x"ec084d0cc6288954", x"13c1b3ff18cc0d1f", x"fb0d7189e819e9cd", x"16ca191c8b3a3b0e");
            when 7754272 => data <= (x"82cc4c4ebb1ab9a2", x"f1e8ec690052fe04", x"e0b9817f17b2e2c6", x"8013c9b8085e2cba", x"1b9fe259d216bbcb", x"8c863aecb977ac7c", x"52a954abd88cdf30", x"2636d92fd8e0fc3f");
            when 31972974 => data <= (x"6dbb48895104b52c", x"af5f580dee2c2789", x"45484ccc3c947e7f", x"21ae7998c9709e0c", x"0b6ed2bd27ae1f80", x"7f102310b4ed78f0", x"e26dee0d86ec47c5", x"7a2d891a091dec44");
            when 30543481 => data <= (x"59f14c2305b67deb", x"d688645ec52bb4e3", x"bfbcdd89f15584fb", x"78c514e41235241b", x"1f6582480f3de1d6", x"38ca042a71258c3a", x"e338960e9fbd7d7d", x"46864ef263e3072d");
            when 25175116 => data <= (x"587529a556afc197", x"1c51c75a675b032b", x"77677173d67d1b2a", x"9fcaa8966f045715", x"045ea5f2288b474f", x"d2facb12ebc239a5", x"1e1fd8e991de199e", x"9f645fe5840ff8a4");
            when 25512769 => data <= (x"d929bc952150597f", x"22c2d82df946103b", x"80533522f9ee45b9", x"3b51980eda23d657", x"8dda0d8f213a59ae", x"37a82818d21b19f7", x"7aba68456da75ea9", x"2183214969d7c692");
            when 12176196 => data <= (x"cb94979e439ee11f", x"5e64d96bbaa2f18e", x"eed7d7c8d4ecaae2", x"e7a073db05312486", x"8ba9b5579938bce3", x"d58b8d50f37aa1fd", x"3f15f4dcecdef9db", x"1db21d681ecec12a");
            when 11231356 => data <= (x"a31f25b37523fc88", x"5f5a91c70d737d82", x"058c12b7e955c312", x"b008ba220b27d333", x"560e4dae07cd2932", x"aa26a334f23b8c4d", x"355ed8931776a836", x"a3571fe6f5a40125");
            when 25235617 => data <= (x"d9eceec48c028cb7", x"76ac0c9c29bd5191", x"4bf0c970f22c31f0", x"5afd1f909a9f6e0c", x"765d7c3fa896f601", x"358b6f423986d5f0", x"d46a26befc0592dd", x"97e4bef582d60f8d");
            when 13826665 => data <= (x"47d7762bc7b48634", x"e25ac1634b9ab62e", x"dcf4585cb8805937", x"4b12fe8bf6c9bc77", x"1a5daaca73560981", x"ac7d3c5efd0898a6", x"a431722c713a3998", x"456ab8cc0cbf63c6");
            when 14779505 => data <= (x"d19fe78348d6d954", x"b49c2dfe89c2c405", x"526a04722e449a91", x"66a75ad1de1ff5f7", x"24ed428e38aac8b4", x"aa8c05719ea77e0d", x"ea5d8d9b78279a45", x"1ebe5d84588395f1");
            when 8774241 => data <= (x"fa3663e65830b6e4", x"1f2e44936c37e324", x"7c82a8bef9563c91", x"93edcb7fd7ad10e2", x"a0d8bbcf1de8ecd2", x"2254e74bc6731bb9", x"2abf02582ac97b6b", x"5cbd1b1e6329a91b");
            when 20781823 => data <= (x"32df034e048fc482", x"dcdd0a110ba3f5ed", x"91153e73c5ce1a2b", x"a8c095af5e560f5f", x"25f8a7db42636306", x"9cb9c00203cd0c3a", x"cc7f2d1b903850eb", x"5ff091f9c2314c3b");
            when 28654244 => data <= (x"05775da8bc695a3c", x"936fafbc6400e1ad", x"a641d9fb19386d9d", x"258a955b7c76f14a", x"68971a3b9b88e00b", x"69b2412ea6b2cfea", x"252ef24e61352e38", x"ad120ae6eda9d592");
            when 9213842 => data <= (x"6e36a0addd235911", x"052f779d9eb07907", x"6d1b2a82f50ba00d", x"24be9570b9ad004c", x"843ab2a3340733d4", x"ea0f100713a67e13", x"493cfb0169053e09", x"f5afeb8ef26405e3");
            when 1556472 => data <= (x"f091393c0785e851", x"1b3973517b835503", x"cdae7c1daf919921", x"345121a5aff067fc", x"deadc4006c3003de", x"624409736e82947c", x"f33822f79cbedff7", x"ce50771908bc2d83");
            when 1266904 => data <= (x"6f3a99f91ad900ee", x"166b891503d9255b", x"d2aea9084acaf294", x"9205a81f55076f57", x"35d2d11df31bde01", x"06d9b12a1d407344", x"48ca017ba2bd08e4", x"e1ec172d335cf8f8");
            when 4968577 => data <= (x"de1afce3cb26de5e", x"9b38d95b160e8935", x"d01a1e28f1c57ff7", x"f2e35794495381c5", x"10bf7ae7883dd30c", x"000b99bcbf103f4a", x"8a592661867e3db5", x"4937dda7f0188c68");
            when 29060666 => data <= (x"4e1614a70cecd540", x"7cf8a1e4773ec87d", x"1fbd025787c51378", x"b9d02f878189a6e3", x"98e62ca04e8581f0", x"bf019f9dd02ec269", x"064a3dacb6782ca9", x"82f1560fb9dc216b");
            when 9829463 => data <= (x"3dcf8703ef8ad1dd", x"ad06b5382a3c2d9e", x"3b3a6a273116da95", x"0b0f9367cb370feb", x"35837ffd477dacba", x"48f53d2c0e040ce7", x"76ae6fda9eba1f47", x"08a830901eb8d239");
            when 17838459 => data <= (x"6ea25148a7e96939", x"65e892e8dad7b09c", x"0fd028f0d2681371", x"291b232cd5fddc0b", x"c5f4b868a41c13a2", x"f2ce6a48705fb670", x"8583de944e44c032", x"000fc147862be3b4");
            when 7962624 => data <= (x"d948c12819672a8f", x"f59c43c556ab0955", x"4b4fac1d1949e47a", x"acb789c2da51ca96", x"b4aa26cd663f46cd", x"d6be7a3ce74489de", x"80232e6217c6f806", x"a5262bc2dab0d2eb");
            when 11125905 => data <= (x"491e957feb6d1e27", x"228de29f5b5862a1", x"b23e33f4bf3e67f3", x"4a2db86bbbfe557c", x"ad4e3b5694cb33e9", x"ba7f82102417248d", x"a5f55ed5ed548d50", x"829d6dbca2aab919");
            when 4280129 => data <= (x"4972421b3f4f8893", x"879adb8762a63a6f", x"eb09b81ed896e2de", x"96a5e29ee631ac94", x"10d985a2b1c89fb3", x"fb0990d8b479708c", x"50bf52896e5e762c", x"b68d48aeb1b50ffb");
            when 13704456 => data <= (x"a911cc480e731d40", x"655b8cdfe308ced0", x"a130307a71088d3e", x"9b891618a79519b5", x"4309ec9ce5bdbcf5", x"785cfbbd60cba677", x"4522c3fbc5323af5", x"d5608c62674fedea");
            when 12868372 => data <= (x"015f1be57c56dcf9", x"c95c34e534343cca", x"0c3120744ea62945", x"cd6ee18e07852d9f", x"20ca696517de75c1", x"ef40f06797c94001", x"8869cfa73c8ffb14", x"d98b1e15b7143397");
            when 22704654 => data <= (x"b49243402bdedd55", x"31bb1ea790ed8e48", x"6ddc267ee1518b28", x"00804180b9c67a57", x"78ca8c0ec876a7f8", x"0f3b81f8536a363b", x"b051eda4e5822062", x"8801da4e08660853");
            when 21926827 => data <= (x"2e08f85cc72e0bc1", x"cdb59fddee5fe7f1", x"b9d02c1df5c25d9d", x"de1d838f8ea097f7", x"48b52b0e062909a8", x"ad8e1f79226671c9", x"e81b3395b5d89d93", x"bdde39436efe8fc9");
            when 12709205 => data <= (x"39d5778c0c803f34", x"6e41d3f5b0d6801e", x"25a44f844d221bbc", x"7adb003cb1518dd2", x"d14a0b2228bd0ba7", x"22078157912b3ced", x"2d838d3680f0f569", x"dad3f17e0a7cc88d");
            when 29558912 => data <= (x"5888bda03fe173d7", x"c6c4712889281296", x"8b19f04a78ff78e1", x"92275d16d5515b55", x"8c67e28208c4b7a6", x"a82d308cea3d528e", x"0c045315a96fe021", x"9a316b4f97a20841");
            when 28573241 => data <= (x"5cf546c418806dda", x"f6b101fba3966653", x"378da7792bf47c25", x"052207dd892d8c56", x"29bb934debbecd97", x"f196c9a7024392d0", x"53176da5b5ef4d1d", x"f751ddd9880856aa");
            when 20131427 => data <= (x"9e1f0334f2bb89dd", x"d90a4c23637e873a", x"b0de66334af10f41", x"0e42fbf6407a3b37", x"6c400e105e26c157", x"e34f4549e4694b57", x"86b6ded4538e9f73", x"f2ce1b298e3d35a8");
            when 5182739 => data <= (x"66f9c60e6108228a", x"a9f081ceab0a8e40", x"31ed6ae60c38335b", x"44f09318d9990bac", x"c707d63f57113da3", x"47e9d27f6b4c9735", x"319c9b4d823d98d7", x"187f8a9d1da9bba0");
            when 24638824 => data <= (x"6bd7356b5209e350", x"46b75dfd05d5bc1b", x"9104a40ad51e5e7b", x"c209daad58212787", x"9e5597663471994e", x"97bd0f1634110a47", x"a2624f577c629a3c", x"515d3f6009d84823");
            when 8301464 => data <= (x"2abd0a2131c04be0", x"5727bd0f4525f332", x"c532d1d4ef15922e", x"e00cf512154c0ae9", x"894a2ce6a40d12ab", x"ada0d43ab07f8aad", x"1505719a26c9249d", x"61f9acc4132bc350");
            when 823880 => data <= (x"4781123952585e52", x"f499bf2b4ff085b6", x"c388bc8b63f0278f", x"37261fb868a9b40a", x"986b35112e6d2ef4", x"7974fc9dfa1f74e2", x"205c33198f13317f", x"d3cdab7a83c2fe66");
            when 33814856 => data <= (x"f014eb586bbfc744", x"a0c4cc164e491c0b", x"6c525e2c2474d62e", x"74b1cb36f703bad5", x"68076a45b8283839", x"24570610903ff186", x"438fa7a3660300ee", x"dd8049d0af247c2a");
            when 9973503 => data <= (x"876ef5a4e24cbe8d", x"1b83d27c9858a7a8", x"52e6c8ad52eab5bf", x"588971be62baa51a", x"951440583b1028e6", x"1bb5fb8d79a906e2", x"e16edd8d2682533c", x"13ddfa6643dc9c16");
            when 14017304 => data <= (x"0cd250cf5d24f2ac", x"5a4177e12038d1c6", x"aa44a024e7ee1754", x"4a5572f42751bbeb", x"57c266992c18e8aa", x"2e6bec94b2df0c0f", x"b4ffb50007c9ab63", x"0139905421ecca3e");
            when 12582484 => data <= (x"40ae1983efb613bb", x"8f1342d1a200bb47", x"e293376dbf14cf1b", x"233731fabf1e1d1e", x"b7e100c38477c167", x"f1490fe9213b7fde", x"fe639c97c642e838", x"29458178de9457df");
            when 4739815 => data <= (x"a5c53e457fa5d793", x"cd121dc1b557fa77", x"06d8c8301213993e", x"a2a282d11b543f6a", x"b8da4470e1fb6764", x"234aa10d946555a1", x"de38e643da143032", x"30f2aac796d5bc6a");
            when 10481616 => data <= (x"5abdc80546e3aeb9", x"8b1fc7019babe1b3", x"d55943033798a91f", x"da11e2d60ef162c3", x"ca7bb593221ff24c", x"0b36bf9b64b5fe61", x"1b945c450afb7eba", x"8967862fd082dea9");
            when 25432539 => data <= (x"39b81955790b94ad", x"67dd1a289e469068", x"8bdd8c3ee9553715", x"8c63a404f17e4a1e", x"d4f41e65b6cda5ec", x"c9832d4d38d7e12c", x"1d545c67094f760e", x"4c43063f23c9fd5b");
            when 23866384 => data <= (x"b061614d18820eca", x"f58330dc1278f5dd", x"edd49e8aa893533e", x"62afe6dbc7667458", x"192df1b95625405b", x"5cf513815701fa3c", x"504401635929debf", x"fe8c24c535d9b8ba");
            when 23120682 => data <= (x"f9dacd7744b4587b", x"61e56d8978b9f5fc", x"2be92967c4bb5f76", x"be21184e4e50b004", x"7ce1d3167e3cb6d6", x"92f0f8a5edb2bd75", x"1a4f5b141bd6e35c", x"2a3669358155a2c2");
            when 33490185 => data <= (x"264a74b3272afbef", x"65806dc66d6fc9d4", x"c5e4b40e18d5508f", x"75ad5308beb795f3", x"e5a3af2023862fb7", x"dce6bcc92c5f8adc", x"e208b7a472ea4822", x"8d400fb45f455ff8");
            when 3984057 => data <= (x"d84d86993e56eda9", x"5ea5a71b3e406337", x"932a8129f7ca6186", x"20aedc39803149f8", x"6ea947cd4f79f236", x"68abf87c7f4cc9b6", x"8f8e75cacd437a72", x"806a886f168a23fa");
            when 2647147 => data <= (x"08dcfaccc0333fee", x"42c0d59fd0a96e4e", x"dbd532e387baf762", x"3de63a7c8ab08d49", x"3bd16db7834c551f", x"56db13da35294e51", x"3f97d03fa6448462", x"ba12353117e3ea39");
            when 28266124 => data <= (x"c9817ad94373bb15", x"f839b17d89979238", x"c74d9f9294fc234e", x"66e912c4c21e5a19", x"f568df9f58b8d439", x"ee7a4595cd23533e", x"1964736c536484f8", x"4a4aad1239b20e19");
            when 12598800 => data <= (x"b4769cc85d8998ed", x"fe5c7b02d98ffaf7", x"4eb7aa6a6058587f", x"dfa47dbefaa56778", x"f77cd4d0169a4e87", x"b732a7f14ba0772d", x"c3c0636b92c03c5d", x"1cf9f8ccd65595b5");
            when 11950533 => data <= (x"08e2d8146129b833", x"51021ab989a4a871", x"b0af4b73e3c91054", x"9a51dbc509deb44a", x"7a73959c70d197f9", x"ea07e5cd7408beec", x"de72519a0b1da658", x"8fda5826180fedf5");
            when 10387400 => data <= (x"93734a68acc57f02", x"a071b7052f1a81bf", x"657abebc7c776b69", x"e864acf0fde265e9", x"ce9ad2b600f8804b", x"af389312564ad93c", x"b5fa48a90b6dea18", x"7025d2efd2a27216");
            when 21174914 => data <= (x"ca8e6bec188d9a24", x"98a714fbd6075f51", x"6eab7b8a1eb7e9f2", x"5c86b9b7e0117873", x"5e2120ef9d89b841", x"3a80ba2ea4f5bf43", x"daca4a23de00cba3", x"16be995d4d35f207");
            when 10965938 => data <= (x"d16d13265702ca7e", x"5edb0fb2db2c490a", x"00decfe67ca51428", x"2995c254457b6fb2", x"d2b3246cd915041b", x"9cfb4b401431d15f", x"d754bb6c2cc3ecd3", x"2b4edceeec4ab94b");
            when 27848216 => data <= (x"463984e95b98b0e9", x"85aa744efc2d4ed4", x"07f603dd10f69bbc", x"e75cc0b04d49e705", x"0bcc9e0ef3239b83", x"4287a2f63178f098", x"2937685be023b357", x"ad19b16d03269ab4");
            when 32299276 => data <= (x"f19c65a1287a7fc8", x"72b080ed113467f7", x"93924641b247fb5d", x"0a4d14f3e7510cbd", x"6a35cc4756cd5172", x"d3e63654fb879b39", x"8623dbf113396bf6", x"6a72747d9962add8");
            when 32320325 => data <= (x"f9e453f252aa90eb", x"9a5df49734416051", x"59f188d8e5d66bc1", x"1b4307dff4d53250", x"7ba0a447e7086f45", x"cff711880de5f102", x"5b718605b99a0fe9", x"2b9a78282cb4c00f");
            when 13375360 => data <= (x"f8faba8c6ce9e697", x"3973019523d4daa3", x"03f5fd9c8484a2eb", x"1b61dd051480a332", x"16c307c1ea0b7c90", x"4fa34ef17d486824", x"0fc7d55c9b59c7de", x"98b6f21735a58d23");
            when 28956067 => data <= (x"afb4c8a7776db20d", x"e1d2eef508a488f0", x"14417e1b43cf1b71", x"d2d052d7915d6804", x"ac015781ebe4a5b4", x"616a94223009deea", x"5dc13fd3c59256fa", x"44196bf28ea13b47");
            when 17972418 => data <= (x"085d9ba11d4adc09", x"ca5f9c2250e520d1", x"940661576f8854df", x"13a07c35bed23aa7", x"ed36e9f54f72123e", x"13ce89ec4b54b6e1", x"fa57c40d36fd411b", x"efc4487bb83cb8da");
            when 12653760 => data <= (x"07c2f0ca3ddf40eb", x"76988122a05329ec", x"88cdd3d8f73774e7", x"c5b5bcca6ffcf1ca", x"af4c3574a54faaef", x"27ce8ba9d8740ef2", x"5c9577da18bd870b", x"d6db083858c7d7b7");
            when 2050657 => data <= (x"11292c127960f7bc", x"7448b4a210d4cc61", x"446034316a72c264", x"eca1a5db61b66b1b", x"cc418730b6a8fa0d", x"9d12c31a1a2ddfd8", x"33cedf255d13d981", x"d3a26dca67bf1155");
            when 28094362 => data <= (x"180181e82f25639d", x"24de670abca25981", x"cddc57f432062904", x"e1ef38a379378317", x"a1fb68040b4a1ea4", x"2504a29ed87a6e77", x"bb5ea5a5d1f8e5bb", x"648fd2b6834f3266");
            when 19393301 => data <= (x"a47ff5acefa21b06", x"bd1a03a0e75c7a25", x"b39370572efeaff1", x"f3d6da7522d1d764", x"d5ad0a9446f2c6d5", x"8c1b82011c11db4c", x"f1808e77bdc79e80", x"cec1449c30d1a76b");
            when 1294544 => data <= (x"ca0bcc8dea63391c", x"67a1be94f2bbca3c", x"d5387236063729d8", x"ab9e4e11b6c1dd58", x"cd5cd9476f8fa5e0", x"9dd6cc530892092a", x"4612be71dcf34c20", x"ef0f3d7050fba8f8");
            when 2091327 => data <= (x"0544dd994146d4b4", x"eaad39d69d046dff", x"aaa2dc6eebd229cd", x"76a9ff6956521553", x"dc701f0ca8079a4c", x"6b75e12283a9ddaa", x"d9694c2f9450a1e6", x"fec00768c7ba2467");
            when 31526774 => data <= (x"5838bf8dc8173c2a", x"386c79f60e96bf77", x"0742b71c7eb5dd76", x"c2885681b48fe9b5", x"a9a9154467d0ef4c", x"313e3e8d9334fabb", x"886f7e77a55c7bab", x"9a5792dbdc794564");
            when 9146755 => data <= (x"3d76f539e91eab0f", x"3eef0b594ba7c5ea", x"4d19ae480859b067", x"3f7071f6e76839da", x"4293c3fdb1cd2cc0", x"58a7840ded923955", x"cf789e305383f474", x"c72f2f6d1ffe295c");
            when 13021352 => data <= (x"da866dcd7e0de1d8", x"66e5b6fa6dbad4c9", x"228dab15edf49f45", x"29d8cb00e2bdb742", x"68a6bc77e7e6ead7", x"2d4b0ea127e4b051", x"b8d7819e89dae4ca", x"887c9f9e2ec961dc");
            when 28281355 => data <= (x"0fdb85e791c12e1f", x"b9dafcf857905a2c", x"9da00323b2735899", x"45a1465d7f1dcdb5", x"d7c65ab06e1bbd61", x"2bec09b240bb2dc3", x"c9d785386d46879f", x"614b3040b4809341");
            when 1960414 => data <= (x"9f56dd04969bcb55", x"b76acd352a39ae61", x"f63c36cc42905072", x"1dac9537fceb285a", x"306af9d525dfd421", x"958c7cae27533762", x"e46cec3d01d69af3", x"a71ff508e3c783d2");
            when 859532 => data <= (x"f0f395ba9d99e6d8", x"eb2ae83e60e8806d", x"004371c02e78174a", x"cc7b2f3ac1378d99", x"faeb354e0033a9cf", x"62bdfa36b4e87926", x"06213085e3e9054f", x"6b609d186bfa18f3");
            when 19230026 => data <= (x"a3a539563a315a31", x"217e6688c19d53b6", x"772b93249fc835e3", x"fdefc4863288a75a", x"3a772ddd15513a7c", x"5d1d436ee824889d", x"66fa88f152b8074f", x"d9da888c58aee40b");
            when 22756933 => data <= (x"d6bae7bb119eb93c", x"600d05767e4ba74a", x"42b8cbdb42a57388", x"901a11a277f7591a", x"7d3b34e751436fe9", x"daf61389193c60fb", x"ca03177738ecf22f", x"89133998cb3942e4");
            when 18422194 => data <= (x"60a1a30dd9a87f58", x"287cbf00ebb9a6d6", x"2334e6c199fa9b22", x"b63b406a2b9f65d8", x"fc6da0273309ec16", x"e954e082d6b33878", x"12f9a12f01f00146", x"e9e8b33cef7dc39c");
            when 33668434 => data <= (x"caa9cca906a33ccd", x"128806be0428b9d9", x"3997892902ade4a1", x"60c2d9cc4532355a", x"423b4b27fbde3da0", x"9281c8d9de9f523e", x"a840c7819a816378", x"b092ec7314b70b60");
            when 7787388 => data <= (x"69682f1f196d18fe", x"ac2557743b04dfcb", x"9ae7c2f36af60756", x"2439d8abb7b40ec4", x"2a268b9ca7f92da9", x"eea620c32a7cd5c8", x"9e6f7b466d4914ac", x"a676108f40a02783");
            when 14800046 => data <= (x"423ae61324e9e81a", x"d391dad4e7c8c661", x"2185dd942883edef", x"7f83e1fe6637beed", x"bae19ff122b92e8b", x"c2b3e254aee0b966", x"e5c210e88a0bf7ce", x"fa21b6e8ba4aace0");
            when 6608315 => data <= (x"354322c5d1a06d77", x"471a760671349598", x"9e5a2502176e83c5", x"58bdd076101ad0cb", x"a5988cb1cb8766d1", x"e7a4d189fe88fa4f", x"70037b18af3de40c", x"f777ff6872234bca");
            when 28041919 => data <= (x"6c7dae64f0d57a6f", x"bfa2633e95fd6966", x"96465afb44bf91a9", x"d9f1ed41d83b8bc6", x"7e539d8e1513ef85", x"df50ebe75282955d", x"2ec6f86454fecad4", x"aea198344d60c09b");
            when 13275020 => data <= (x"2ee9c0ab64887dd7", x"30a110ac86735618", x"1eef4ca6275609fd", x"a34cc1d64063bfd1", x"ed347aba072db221", x"2298692728cf5b4e", x"11dff7bcb8efd846", x"905e139374c863f0");
            when 28507119 => data <= (x"f95a292b79d0c119", x"f2b2b14f3bd9532a", x"4caa92a355c4df61", x"45ee69bc1816f1e5", x"793faca363150d13", x"fb8accde23bd372d", x"ad56472e6e8b4b45", x"26bccda20cb7b012");
            when 11854531 => data <= (x"11644ae0c74d3626", x"71e814d4684f485b", x"20fc10d1210a07c8", x"c79cafb54e1cbeee", x"6c63ffc52de08988", x"b7223f420140181b", x"235cd0c81a763fde", x"686266567cfab50c");
            when 3260447 => data <= (x"0821c975014a8d92", x"71fde432977df78a", x"039e6c76accd1a09", x"c83d11fae09d7900", x"c1bb9e62ed81d96d", x"d1bf54fb6f362c55", x"b80fbabe7aef1ed5", x"b5261e318f851a76");
            when 28778632 => data <= (x"12580640dea915c3", x"fa94a37bd46b9f36", x"852ba249180682fa", x"57ca50b92603a943", x"d93a140c8d92d0ac", x"18b03e5fab7ba8fd", x"d1eb3368aca349de", x"d70b4e6fb2fb8cc1");
            when 9119812 => data <= (x"5efde625c0ddf9db", x"c61a47324012e7ae", x"26e5c7d22b73dfa4", x"88ee2ffcc644a1f0", x"5975951a1ee96e0e", x"fc56d6924ac805f0", x"35d1fc7e21ef45b7", x"d93fb9f02d38a207");
            when 4546868 => data <= (x"c8bc632afbc2f427", x"be70c7ab44a00151", x"d331aa4935d49b5c", x"74b3da5d7de259c6", x"8dcaae346e091448", x"3047a517258df383", x"60390074841d7577", x"766c67d8ce7d1cd8");
            when 22089156 => data <= (x"cc27a5a8e28d6eec", x"57c06f00b98530ca", x"9d06728c13ad5a7b", x"3dd41481fa6eeab1", x"3594271c49dcffb6", x"a04e4165ed5914c1", x"ee73bbad39cb87fd", x"cc80fd5d75e06dff");
            when 6770790 => data <= (x"0df9ec82f335a0a1", x"3c7307b0f82f5cce", x"9513f604455bfa21", x"84e5b56059b7320e", x"d3f9bfdc661acf07", x"0ab4e7f27db7e9f3", x"c043005e88d91d86", x"7f6c8f47fbf2ee14");
            when 4901171 => data <= (x"50613f9ddd76583d", x"caf799975f51aa73", x"0bb7b92488bb2b3b", x"3fa8b8002961c477", x"97879cf29201933d", x"548d7e705ae5939f", x"f76ed5d85ce6ef6b", x"aba07534a0505ad7");
            when 32076372 => data <= (x"623841852f4490aa", x"1ae944b253b82b0f", x"bca89ee58bcd5366", x"7cf6de9dfecc958d", x"5e31dee85c2df71d", x"64bbcb693e04db61", x"5f80e388d6efa584", x"38bf4c924c077741");
            when 1657210 => data <= (x"50f78e07be6c6fa1", x"dcb05a9ff06bb5ce", x"968e915282b72ad2", x"9a89b71ae4522232", x"e388e28fb0d4e5a4", x"0bac18e78ddf2826", x"57035c3279d5ac89", x"decfe83a07e47b2d");
            when 19011373 => data <= (x"9a6ec5cfcf0d8892", x"26ee6b2e52ad68c1", x"f4cd81428c147b94", x"eaccb64ab86e7b06", x"d9d467b50ad45f9d", x"b325143970060042", x"7761c93a63f9f39a", x"62e8accc85e1d9f0");
            when 30795705 => data <= (x"afca29ee55315eb9", x"532d13a7e28f49e7", x"8f66f71296e03ea7", x"3316d21e41992b38", x"53a39297a33e0e45", x"d5213110961363e8", x"3c8b5115a8849327", x"feeb8e2f166a71d8");
            when 30197985 => data <= (x"6a7913aec3f0fa55", x"ec91d2076742bac6", x"b44f5b7e28f2d47c", x"33b72389256a4f30", x"6357fd316a6f2134", x"5172413559284378", x"8dd9e93830038ec7", x"b387e0a219f9826a");
            when 723259 => data <= (x"8a5a69dadb372478", x"5fa8b8c173b3c808", x"6d100e993c1f5ad5", x"df7af1dfecf367a9", x"533d56cf1558fe1e", x"ae301a8a2d349643", x"cba7ba0bd3efe00c", x"a2d04edf28378b23");
            when 562913 => data <= (x"cf157ef9748bbb04", x"5d0ccd1751403710", x"2a83f9eea27625cb", x"e9a87f25e0026dd5", x"f4f2aa4050d9241c", x"86a7781f6d00116e", x"4961267aab38e256", x"8b8cf5286b5ddc68");
            when 31187711 => data <= (x"a3873075c910809e", x"8bce820b45dda7f4", x"b94cdd5282d595b0", x"6c473aececbd96f2", x"22b5636b31553811", x"407f1ceed2726f27", x"5ab3e0e375aea0f2", x"22cbb70fbc5ef8f6");
            when 8156700 => data <= (x"231c2f4c6e6be45a", x"9e718c9bee5bd4df", x"aca48a6b39f2e257", x"44e1ae5bea3c88ec", x"d9bb834fd36b2a08", x"fb69316e36687982", x"1b8f69761f2ca534", x"8155fd2c4b749b00");
            when 23482768 => data <= (x"6f09539ecad3d06a", x"3d20942a390c915a", x"07981bc717b49f37", x"2bf70a4748ffca51", x"5f7eb923a7497f4a", x"eea5426639f9a23c", x"7e71fe66b50f3238", x"e80d2617f4304e4d");
            when 15839428 => data <= (x"ba7f05d867090079", x"4dac1261c44213b8", x"1a3afaf32f250b65", x"377fde5dd51a58b5", x"50517472b5511691", x"da5e50f362fa3990", x"066e8868a93d30db", x"b350682a11d549bf");
            when 24212092 => data <= (x"d71aae1bf4b908ad", x"3b67f75acd239eab", x"219cc3436ede863d", x"d2792235239c025f", x"48b4ae0a5df22375", x"be55b083729f101c", x"3c21ec7f14523a4d", x"ecef380bc477e6a8");
            when 4210229 => data <= (x"087df25d5a045689", x"32b525b02cfcbac7", x"797c92bf95da1cce", x"0aea1f3c05f1e8f5", x"5cf613448afb19d1", x"7bda64787eeedda8", x"cb1ca0ee84f5465d", x"c4d90e473f321969");
            when 29767066 => data <= (x"f981aee51acceed8", x"b9bde30e1275051b", x"6ad4ec3735a17c18", x"78a7471cbd73dffa", x"f5d5c64701c24810", x"c02b211889f7fff5", x"17554fb9d3d440a4", x"e23185f2edf3f97f");
            when 15049411 => data <= (x"a3a7dd92da61b024", x"ae34495ced42290b", x"f86ed50e7d09bd6a", x"eb9bb76773591fdf", x"96199db371231432", x"ae734b887afc468e", x"d180bda6461723da", x"9e1e948634765d14");
            when 22992898 => data <= (x"dc97c4db597ed6f0", x"767d6bc7ecab62e6", x"ad7047c6daca0ca1", x"7c3f924132cffc6e", x"02d62d237fc99f3e", x"fac0f23f957d2f71", x"6c836bc5f6495510", x"a9294b3b4a0cc39d");
            when 15324667 => data <= (x"ccd4b04792b029e5", x"e07bb86eaff01da8", x"aad1b1c70c95ea4f", x"299a597c996d8370", x"be361fe01107e432", x"6876303f373feddd", x"d8101e614ec87127", x"8caf8ecce18abdb1");
            when 20856030 => data <= (x"a5b4bb18506a0508", x"11ab1f7266f8a6a5", x"7b21151ef5f272f1", x"8290117199de94d1", x"11a11aa43ccdf454", x"c5618dcae6a6381c", x"ceee7681edf199a9", x"484b407d59b484e4");
            when 24964057 => data <= (x"e0e1ce78d6e108e2", x"951fad8cf19924b6", x"8623317570e57ac4", x"597fd0f4d045d82f", x"1facb18728f51b60", x"f76fa4232cd541df", x"a6b74e34fced5bf3", x"cbe008b2f74092a6");
            when 18439569 => data <= (x"c73d940ff66fc603", x"edd76cc8e3834f98", x"e8cb2d74128ccef8", x"d156f5b88b7d194a", x"e1a599fa84722a30", x"7ffcd398d6f0f808", x"444c808f8ee37ada", x"dd910c48aedbfd53");
            when 12957440 => data <= (x"8889730fa849483f", x"b478ffb915174bc9", x"049bce2636ea5c4b", x"5cdbde8bc9c9cb6f", x"a72a7b6cc360c2ad", x"eb2d572371270ed9", x"29ac9994ae31d27c", x"cdb7c4affde52895");
            when 31643670 => data <= (x"49749c688209f0c2", x"f1304498c7fc2111", x"6867ef1b4c6a494e", x"840f32fa66edab20", x"07f1fb7b41b338ae", x"90beae5bbfcef75a", x"265123ebd61d51ba", x"e9961e3bf5238440");
            when 17379567 => data <= (x"f2d398c5c66ae306", x"c9aeb6a8748b441c", x"a32ef2e8331e3de2", x"59b4516b87ce3ca7", x"663e2aa89d454c95", x"202d1bf14b9826a1", x"2b920eb706aaae8e", x"e494d7d269e39ee7");
            when 17307522 => data <= (x"f8143e4f7cd92cac", x"852cb38c2e485157", x"7881d603c1456f04", x"1dbb39f98e24c2b5", x"a98d932f3f4af3bb", x"1794a35e513fc745", x"cb4d8c5cc5257926", x"a2635737b1378b5c");
            when 15294290 => data <= (x"761ee59577ce076c", x"7e0a28e53ebb9254", x"98b8970d0d449446", x"519dc5b0a4631b3a", x"7f0a143658ff9d2e", x"0b8e5353d1faa664", x"32ef2b419f204a6c", x"5fe2715f6ee86e55");
            when 23456001 => data <= (x"258084f1362647c3", x"f7edbfbcd020f02c", x"2784b1d66398bad8", x"255132294b07c1fd", x"3d804fa036dd3a19", x"6091703ca5819258", x"63a5d4623f42c6e7", x"3b0e6e634ff59fbc");
            when 16628877 => data <= (x"fde8cd237d2f4cab", x"ca048a981f55e302", x"f4f75773feab6df0", x"838ca6dcf891e45c", x"8f258550f94d7abf", x"ae634eebc048720d", x"5a280752178366ef", x"f7c7aeb11a2162b1");
            when 23947840 => data <= (x"4cc0b4783a7cc125", x"f466cc81e0461000", x"417968dbb835fe02", x"40f7f24e3d27edb5", x"b570b40294872ff6", x"c5413dd9d5ee88fc", x"702111938f866277", x"8a3f30c7f059c142");
            when 1307204 => data <= (x"f810b1debe373105", x"c54c905573e44ae6", x"a9a751c1238280be", x"a0eb356e61ad8f03", x"dbeae03734e7272c", x"4aa6d45b7829d377", x"231ff8064da4fad0", x"b5a99787371ace03");
            when 3700012 => data <= (x"7ac3478867dbe147", x"0ea4f6947cadaa92", x"9493812c5d6b84f6", x"150113840e2f2368", x"2185854fc9919bba", x"98664ac37b1caf1d", x"a62c3e1e6e28a88d", x"9ce2bf1d551453a6");
            when 30500541 => data <= (x"bb0a1d69ebe6d40d", x"29842fd02bb33ec2", x"851ee890801c2468", x"083af3594b3677e4", x"8713c9d001167cca", x"3ab38e8b70c9e56f", x"0f93ba31c57d715a", x"29e3ed0e4b5b4c5f");
            when 4399260 => data <= (x"ec74cc1c07c0ae47", x"7a130f178fccfd06", x"f9f2ab0eaea16d37", x"09663d8cf23728cf", x"2b0eee75572a1e66", x"1098d5cab2335d0a", x"dbfb55a3c78b8a81", x"0b46e1d430eccb93");
            when 16650958 => data <= (x"d1a3ba2c9956f88e", x"243a50d73960f4c5", x"d75ebfd3e1272b67", x"f127c701d77b4208", x"ba840e4c9dfa3a82", x"313a96c43bc0401b", x"2954d070d189350d", x"5b8b4fc836fd16fc");
            when 11137186 => data <= (x"ea67b87f3b0d676c", x"e271ae189cf09381", x"a437377617c61464", x"939ae33e86afe180", x"5e9136b9e5d40e4a", x"f3850a2e3682d82b", x"ba250498dbd92a9b", x"5491855124bfd726");
            when 5422939 => data <= (x"b4a2393150f9fc09", x"6c3622791c682e44", x"6fa9b5f71890a1d4", x"187d0573c3d1e051", x"0f13215de017dbe8", x"852820f2d2aad665", x"ecf922454aa32253", x"55c05a575a54c522");
            when 10013302 => data <= (x"84465ecc44dbc399", x"5d2015459f46adc3", x"1a84400826fea513", x"0df969f5fe356897", x"840d1972ede8a776", x"1a4c7f7190508430", x"94460b8d7e5715f7", x"e4a50f1d7c48a22e");
            when 20552244 => data <= (x"3768f49cf2e9bd8a", x"f8090ebb60b61e30", x"0c2dcb6126774d47", x"fc205e6ceb147079", x"0b3e3e3379973bef", x"e8f4406fd9fb4ef8", x"7dafc9269c3fbd7a", x"9208954a2aa0bec7");
            when 30280769 => data <= (x"552f7359bcaea43b", x"3e203b417389d1fb", x"fc1b20bf4674e080", x"12d7d1b54795bf78", x"1b94a4df6b865f2f", x"d5777e5c300418aa", x"40e506b29d74b3a4", x"0dfc4fdca0f8d498");
            when 3289535 => data <= (x"1e1919cc2b8025c4", x"3a0b091291b62fd8", x"9334a57584854149", x"263d5f8e9507e4ab", x"c69d1ac7ac9180e0", x"497d3dbf1ec8da44", x"45b30ab08d5a3d2d", x"0ca995185ab788e1");
            when 20550820 => data <= (x"33954b506a76c50c", x"72043acc37d75fe2", x"ce7f668bcbf689bf", x"aa97ac93d9e36971", x"cee4b04cd9634887", x"2c9274e2601280a4", x"4a5e35b4f3e2f9f6", x"5ee0fec04d8328d6");
            when 24518323 => data <= (x"4a2fbef56b6143f6", x"23b2252f6a5fc253", x"8105fec10034f6d4", x"42bb3dfacba0f184", x"07adcfd1a3eea279", x"066d841fcb5c91aa", x"0c5b09c677aa6b6d", x"58873fdd86f30886");
            when 12236688 => data <= (x"dfd7960cdf26e427", x"2973f26769479720", x"3a8e6bfb52e11970", x"d3610a704b6a3047", x"0802b19fc7b6a7db", x"4be203115da482c2", x"4fb468d3b62602cb", x"f9bdd90bd569c10c");
            when 11367238 => data <= (x"8b7b9d5d8f84216e", x"697060e3c9888c20", x"069b5758f9ec9fe4", x"478611928fdf0573", x"6e43bd9bc9c3859e", x"581000a0f9b049c7", x"3df6e8ed605cde8b", x"94f642152cce5664");
            when 7409007 => data <= (x"0108113aa2dc5370", x"3f47b60582631b1a", x"ef38b2b661f0e76b", x"ea3a2c5a5669af5a", x"28fa4477b60919c6", x"24cf7af941090ffe", x"de27998f6dd6fefa", x"aff69f7723d3b317");
            when 15861553 => data <= (x"6cfb877832009001", x"c297b1280f40fed1", x"1aa63952b142d679", x"a0a78d51da6a510c", x"85764debb87e085f", x"cedc76a47316227c", x"4bdac59b3b70306d", x"622fd90210832d07");
            when 4178934 => data <= (x"e3919ee33361532a", x"879c9e13083b92cc", x"fc21d3bb9ec403e4", x"e9ee5eb0eaa381a8", x"a19b7c1a539925fe", x"5c5d24641417ffee", x"bcb992c8003b196b", x"d0d3622f0fe7893e");
            when 23785099 => data <= (x"a2c93cd5a03ebb5e", x"c692fe094bc2da42", x"2e4c33193d0e9b91", x"e080aac2ff375fc3", x"2705771b810c1be6", x"9ca86293483acfce", x"36aac217076c9f9e", x"30200eacaf4465af");
            when 9797135 => data <= (x"03904a233d474955", x"564c9000fb5e1188", x"17fe2794a8a6cff2", x"5280758802ef3010", x"0997c4e5011d7928", x"915a45e4b9f8d650", x"86b3ec14a3f23739", x"2f9b2931110a7f9c");
            when 9892828 => data <= (x"fa02f120419005a3", x"e18ad6e803e51883", x"2df419bfb6f9a217", x"dcda17975b0ddbdb", x"11f252f36919a5d8", x"c3e230195f1dc572", x"659426f78ff63a4e", x"e2252a3187eedd10");
            when 12204411 => data <= (x"5525139cf4f505d7", x"bc0a393ec3590f81", x"d80c11f717bd2a35", x"b767594593c8f246", x"2f4f297f88d8ec26", x"99e081e1fbfb2404", x"f0f714bd9feb5adf", x"17b58efee93d5731");
            when 1847704 => data <= (x"e8afb27a20615e8d", x"8688fa063cf1440c", x"ca6f55bd90c39e18", x"8a42111864e7e706", x"4af317df6f3fff62", x"43c2289df245b797", x"8ca71c08f128cd51", x"8be34ddae533d8ef");
            when 24384029 => data <= (x"1afbc2de29664048", x"663be059b224dc71", x"efeeae613173955b", x"413d122b8d89009a", x"bf91c3b3e5e1a3ff", x"ce501e7f07a4a89a", x"b9c5f81dfc0b0fec", x"c9d07cdf87742a44");
            when 25444570 => data <= (x"47007208dbb4b3ce", x"97581b0b2c5e8b6b", x"a4552b97fca62683", x"2f294823a0fb6ed5", x"8d268fe3f7fd01f5", x"a2a4e3f41ce41485", x"115ac082fdde6320", x"47bfd4e89cf0f662");
            when 6371996 => data <= (x"c437ddddc0c078fd", x"8cac49390fc62411", x"03d7bf4dd2c5db76", x"65bd563277e8a862", x"5857ec6d8d556bdc", x"595d0994fd45ecaf", x"061926f65b4fd149", x"66314a1503c4dbc0");
            when 2680878 => data <= (x"11522e164b671ea5", x"b70c5728dfaa5261", x"820304ac6ab2b5b5", x"fd92a70b12cf63b4", x"1092e853b0d58193", x"c5d70195d1c0f863", x"2a52e7db96f394de", x"2743299c61955ac4");
            when 1294935 => data <= (x"ddc2ebb30edda958", x"5f1133d10852c4f5", x"211d2fd30d786adb", x"18b2086559667343", x"c69645eeeb748bf2", x"60c7c6bb40824efb", x"fe67520e7ff7125b", x"df9133f1b3e9a81d");
            when 7724248 => data <= (x"444ac3947f1bb51e", x"9ccb632f501dca4e", x"c6e0fbf76282d073", x"1935ff17fea98dd9", x"a7e9ebbb8b95eac4", x"b5d786cd3bc79932", x"8e9236e57f9b3505", x"657379bcef4c056b");
            when 31904635 => data <= (x"fa4a06eb3bd145ae", x"9e202820708c8071", x"b1279bfd0db4e5ff", x"efdfcd69e3639a88", x"07a5f10e20e39e5a", x"1d55a7dd0b79dd61", x"581f604da133e46e", x"e6343eb25044e22a");
            when 2934902 => data <= (x"884a600a7556ae9b", x"0ee5125951102d6f", x"6952fa61ec337cbc", x"897664f5f3ef06a4", x"a7747efaf92f8900", x"e9bc13bedafe6215", x"fee0be4a6bff1d3f", x"3af4fad80abe86d1");
            when 21673462 => data <= (x"fc8dcb3655b7ebc4", x"625da1ccf3ba44d5", x"31a384acb84811d7", x"558117a791881865", x"7d1525813434bd02", x"7174ff991ccc5416", x"d2f7fed497049776", x"b3f289d1c8b8af39");
            when 6650834 => data <= (x"3f6ad16fa2ceb384", x"263501965f5c0485", x"7e5d45e35e56b1ba", x"774c77248458b63c", x"9dc16053da5c27e6", x"c985676bc776c406", x"b2cf950048d9ced4", x"ca3db6a384d2b6da");
            when 15760246 => data <= (x"e1b8c0700722c22b", x"1d21c09c8ee53027", x"a6bf15aff5972850", x"601f20008e26c1f6", x"ea261258e3d2b717", x"22a0d4df8ed0e6f3", x"52ad48c32d59dc81", x"70ebb0d2d0350c43");
            when 17721166 => data <= (x"264d46d27253a0ac", x"04f4d68fc2154dc0", x"82552b9e43b46a8e", x"1c29e646b90e95b2", x"ddc58e52777702a9", x"4dcd9a1b6f6b4460", x"8e7e65c7c829155e", x"1511252bbffcdca1");
            when 6153422 => data <= (x"f9ad3ecbaf9f3b90", x"242c3d089d375a08", x"42ac090b915fbc40", x"5bbbd443cc1c83cb", x"8852848a593b3346", x"ca00f3f0e50e51c8", x"8b8a8f4aa8e22c54", x"1a5ee98e57229c4f");
            when 23773935 => data <= (x"4edae7bfa885b16e", x"645077077ec5e68a", x"f377d3a8232cf6ad", x"0e63c42801a4a681", x"a8bc7378d8e91d61", x"36d0edbaf2defde1", x"fa3a5de948ceb7af", x"93410ee7350a35bd");
            when 11634333 => data <= (x"435af13fbe121d64", x"6e5f408c13778420", x"6bcd844567f9fe74", x"d08aae3d298e15e3", x"4a1edd0cdadd4aeb", x"8f1ba37007928061", x"ca71ec7a418f6b74", x"741d5aab853ef9d5");
            when 1152561 => data <= (x"5a3f65446d4c265f", x"70df02be8398a6d6", x"5e6f79b779de4f8f", x"7dc9873fbd878eb7", x"8f0f5dd68bcfca5d", x"6c9b140347db5cbb", x"dbdebb6402b8a76b", x"b5d712198a95ead6");
            when 13651462 => data <= (x"a229ce9d3f358627", x"c9b05d2cb2ac142e", x"937f1cb288e3abe3", x"ef21e869a4e30334", x"9510a5fa37ea8d8d", x"64855d0e76fe3c8e", x"3aafd052b509cc0c", x"8d94b80b01e150b1");
            when 14244536 => data <= (x"f695d7370f632d5e", x"5d65c4c011b463bf", x"99e3e335dde3ad69", x"d0c1934896e9d847", x"1c0deedce43ef1e5", x"3d258ee81ea03454", x"9a3e9ee23426cdff", x"7682df724bbbf85e");
            when 27622770 => data <= (x"6090b1a1b6b374d1", x"826b9026661fcacf", x"e36806968ea151b4", x"bda06de2d9aded2c", x"5d54d035e37e68fd", x"e2343336b5a4b1ff", x"44d23009f54fdffb", x"0efa2c96ae208204");
            when 23002198 => data <= (x"aba969af15ecd3e4", x"a737a1b356958db7", x"563cf518908610c2", x"196d76c40a6cc9f8", x"f60f726c98cad390", x"68764ceb9d45f5de", x"f55645add5c17c3b", x"05118840d69ddd17");
            when 25470031 => data <= (x"26d01a61939c8d88", x"6c71b4f04b14eb2f", x"0ba0f3b977ed7eec", x"ccd6650af9f7a6d6", x"8de42fe559d9e703", x"70b135ad623f396b", x"632e93b7f3f0e364", x"958e0cced8baa15e");
            when 21745439 => data <= (x"a30f37c4b512b7a3", x"5baa36223fb59743", x"343c299afaf6f693", x"d6a2e5b03ba7331c", x"fe1cb425a9182299", x"88edfdc3d01733b3", x"581f3d6446d4b532", x"18b2553bb0f8c6d5");
            when 31186840 => data <= (x"fb80d643d25142e2", x"bfe4809813e117dd", x"42d1d72768ba98de", x"e45b6030c179bc6e", x"e5ca0d41cd2ae24f", x"f54e2722c9e7d2a2", x"716185b333823b30", x"23f79d9a7af0c3df");
            when 2913925 => data <= (x"e4befb99f14d9ff3", x"80ce2f1cd8f602c8", x"0332d8a4191508fd", x"70efef851c48248d", x"384ce2763c0af94d", x"1395c19fb9fa694b", x"d6d759b181cecf76", x"e699bf2cbefb7289");
            when 25035243 => data <= (x"e5b9ad3a15ce5ab5", x"50b9a277fc79ffc0", x"7f852d24b70667c6", x"9ac785b97318161c", x"00acf5dba576932e", x"37825b81fea083aa", x"2fbb40648a281426", x"e37b3cdda4fca063");
            when 4857963 => data <= (x"ad2dbeb056c8a084", x"7ad55214ec8bb1e9", x"c1a4c492a238ac0e", x"e4f6e9ee248ac676", x"fa5efb35b1b25308", x"eee597914aed1b1d", x"9839f270efcf0724", x"312d72514f12b403");
            when 19034709 => data <= (x"c42f37cba1935545", x"c46e5a6a6cd0feea", x"92a39cc0ff447832", x"d85418e21de4c9d5", x"4981237a06bb0f5d", x"0b86737c681698ae", x"9ae1f38da05263e2", x"00fd08f8d79b7982");
            when 19929503 => data <= (x"32d493e6c0d294f1", x"2daaddfbdccb7090", x"8751306a41dd6d27", x"3a8bd37f43e70830", x"216bd59a3dfa8147", x"bcfaa4dc0e20caf3", x"edd42925b356c58f", x"dc57f3a458079118");
            when 6475230 => data <= (x"e19357d326a5341b", x"4f1cecfbbf5c5c80", x"2ad52fd548d7a9cc", x"46a9c80dd7dd483d", x"003a81d1ae283889", x"32c59ab29abf2f2f", x"e0eb4eee74a1ef5b", x"b864c57b46f8e1e5");
            when 19466330 => data <= (x"9ab519e4ee8ee07f", x"2bd2c5f8fbe19ac6", x"76d747560c1be226", x"d846bcd7a10d389e", x"265b9a17bdbfc288", x"c8542158b23f6036", x"ac361c710af0c444", x"a420ba87ae595a43");
            when 32662025 => data <= (x"d50a82c3b6d06a1d", x"14cd84728ffb6eb5", x"15e50218b704ee79", x"80cabc2e15788c8e", x"e2d42f857bde04f5", x"a2926843928e2e87", x"4de15c3d5147aba5", x"f69bd5051529a7de");
            when 21546452 => data <= (x"77238b739c3f3b74", x"ada05033fc340fed", x"deea7b87f90d7c3b", x"988c31f437793185", x"3a40bbaefd0a9089", x"5fec23fa2da97631", x"4ac196fdb999c749", x"1ca3a438c5701e73");
            when 27643395 => data <= (x"7e1600b2cd2e5025", x"905c72b14ec21741", x"c34cc39a9d392865", x"f22d0de32d055aed", x"0e04a97888a9e9d0", x"166f35ef7dfe5070", x"d959567cfc4e64ef", x"e125630e80ae175c");
            when 1523429 => data <= (x"46a7f912c3ae69ac", x"20618e2db29e5015", x"88fbe5c3c7c045b3", x"0796797e5e11ecc4", x"bca0e12dd34f959b", x"ae115814c02a1a9f", x"d04c1130b3ea8505", x"c742bfb8b3f2b9ee");
            when 2439580 => data <= (x"864baaa26a683b4c", x"b7e7ab092a76effd", x"7f336608ba9b6e6e", x"3e49022fbd36ee77", x"8fc9343b9ff754c9", x"efd6d15b21b636f3", x"b4cd187f18f18ce3", x"2864e84d5c3141de");
            when 16613695 => data <= (x"ea903e18e5deca03", x"ba64922081933e01", x"7550ca641aa04a2c", x"5bdf517d12ccc247", x"e34330431ce6b7fa", x"f5b2c51f576c087e", x"6080c5127ebe7ec2", x"6698a25132de7d1e");
            when 21989624 => data <= (x"11dd40d26994836f", x"522a4b914c995f5a", x"04d4aa3219e94be4", x"16b61802ae41f4f8", x"af55e088bb9d43e2", x"82d365a3cd391f56", x"0f69eb673f9a2770", x"6a5c076b613a9d21");
            when 15690069 => data <= (x"08fb3d1b73bcd5b7", x"5ca2f2b7fac8e89d", x"41b1bc3382186ae2", x"13534388ccf9744f", x"66cdd91dff012bed", x"392b16d6d58af64a", x"0e2eb2c4b0cfe9bd", x"581639f18f330233");
            when 27318988 => data <= (x"ea54c422ba0da812", x"0b5d675d8e531931", x"40fdf199b0c61a55", x"af40f8e77e6e5b44", x"8d832c8ac90c7061", x"581df68082703fd7", x"58c6f474f5ef2cf1", x"946fbde9c92411ed");
            when 7442379 => data <= (x"e13e5eaf93b9d762", x"cbc83e25292fc4fe", x"1aba6ea2e28e8fb3", x"12ac8f8bd2dd883b", x"172fcf65d46bc42e", x"38508fa2805e0d23", x"12359708f1daf0ef", x"f1989319fbf162c1");
            when 31599598 => data <= (x"3d1fbbc2749cfcaf", x"6672bc3a55e42555", x"eeb46bc510cf8968", x"4250c0468082b19f", x"f4c3b0f859eb4ae8", x"dde50021922f61f6", x"742e761bc88e9fb2", x"93c3f0ec33008b73");
            when 21223256 => data <= (x"c599b6f4cf9f6c45", x"9281cf4bfb83b44b", x"6b8213b0ade47458", x"29637fcaeaad2ede", x"593d0a39f551a76d", x"7bbcbf4630ceb272", x"73d97ac4d6e37577", x"0e2f18b10f037241");
            when 27677866 => data <= (x"fcc2a2fa9e00139a", x"265002a2e02f760f", x"f9ca8456891dbd08", x"20cf16338f8a8d03", x"c8f601df5f5cbdd7", x"51bf097177fde7c4", x"76c5730bb53cef07", x"b84d1b81db4d8918");
            when 2276677 => data <= (x"1f1430db6bf644af", x"862fb20d400278f8", x"be1cd6a7f0f3ebfa", x"8eda23e7b9495557", x"71db48506f0e0d33", x"172fa5b319e12d7c", x"44c2c6aab2349a33", x"6bb430c3468e5f71");
            when 5617988 => data <= (x"95e124a8e25e1800", x"b15d79f87c3096b6", x"b8485cca4736f26e", x"4ed172f741f57045", x"74cb886454f7d864", x"e3ffc2cd4b56a663", x"df0163dd6597b339", x"2a200d0b2846311d");
            when 12618915 => data <= (x"5a553bc152f38c05", x"d4ba9d8c65adff28", x"8a3ee84a16f696fc", x"5eb499207a5476b9", x"b015c21e9b9583f1", x"6d8c5c723920721b", x"84590a6387073f07", x"c1ce2f7539e4bcd7");
            when 21826392 => data <= (x"7870701ad4bb90b1", x"dcf0ba9e6c697d43", x"e3b88095abbf90df", x"e7252a0a6b3f72f2", x"ec78b8f61516f1f0", x"445fbfa93ab44f3a", x"60238f5f63d0ae35", x"86527caefbdb3b90");
            when 21224616 => data <= (x"9aa10d3c7b01382b", x"890e29d8ac9075c5", x"baaf89508a9290a7", x"94582ff3920effc7", x"d3cb153ecf755d1f", x"df856b02f80da225", x"ba27cef8eea66a93", x"8f5cee7ada944bda");
            when 3908258 => data <= (x"e81421d74138396e", x"810bcfb647a09222", x"6f47e3c2412e3cb0", x"2a0d60afc9d52015", x"ecc3c5de6a4d86cd", x"d0cb03fe4820d403", x"806762f7132e1b43", x"7ae3564d90dc5e05");
            when 19660136 => data <= (x"606d879a3ebc8cee", x"4f5c0ca13fa43404", x"df7e39292964bda7", x"03b74abc9ab1c6d5", x"7816799b824b75e6", x"5b7f07512a14380e", x"e193d0ab4017e7ab", x"962577dc1934c8e5");
            when 20976591 => data <= (x"ef5d01e0f76caf1d", x"23ac1137d56600a6", x"d8a4ac1d60df079c", x"09c8cd25a4b80c1d", x"07913b9f5ac12e29", x"96507c17705d89ba", x"b252d19f1d80a66d", x"127ef40ae5a6d931");
            when 30022323 => data <= (x"5f30e2e3b8c6718a", x"d588d58876643205", x"51ec9c06691505dd", x"da27890c47080084", x"948eb8c086b8e276", x"4e5e394198d43eaf", x"d50cd5d3f96e54ac", x"0241afe83ddbbfcd");
            when 24454924 => data <= (x"f0185e2519f88a51", x"2e073b429e6c9768", x"dcd5ca79faf82a84", x"cec2b4bfcfe2dc20", x"1083ab712ff45ec1", x"de99cac89332cd2d", x"71ca6e40919268b6", x"475de9d5db1206fe");
            when 27478972 => data <= (x"69adb955c19c2b34", x"9481d3b60f940684", x"6daab732acc171c0", x"08585f749b7c0cd8", x"6cba3826669d9c1e", x"c4a4363940b5ddb8", x"18122829436faff5", x"179fba6f3dd2278d");
            when 12330081 => data <= (x"e543aa343c3f2172", x"b0d30407dcc9d9d0", x"88bcf1dbe73c510f", x"27c015e34c4bc018", x"7f8bdf560a5a5e75", x"0da4acf6b1dee452", x"2dc85c07618542a0", x"3bfba412b75d681f");
            when 4298304 => data <= (x"e1a57f0275c6a8f5", x"a2aee08cda44949e", x"d5494e56bfa2e89a", x"23c1c3dcf6254822", x"aaf4226512c98ded", x"0cef3b77f86fb2eb", x"50b8da5bce3a1676", x"c078f6597bf2024a");
            when 13020464 => data <= (x"f5db0ce828738aa2", x"2fe743552e6659a0", x"3d814f4430df7de2", x"9cf1e62a41132626", x"904fbb6d7527735c", x"654cd386ab7a6ccf", x"694e097842d035e3", x"209805d59640701f");
            when 33395848 => data <= (x"d35c8df23749b830", x"5cacfadc2f4a87b1", x"9dd69fcf37db0057", x"645142da229f917d", x"eaae3e229f6bbf6c", x"55e20f261be450bb", x"5a1b0b68bbd53e68", x"a65f540c3263132c");
            when 32284484 => data <= (x"eaabdf53a259310f", x"e72e423f7289f2cc", x"fc588be7d40fe262", x"4b2335a0e85f7193", x"e250de269a2b65d1", x"948c9b658a14df0c", x"e6c8abadf374f72b", x"d7ea06886f1d7b72");
            when 8008678 => data <= (x"c43eae164b8d5b75", x"f9dc7cf3fe404528", x"4dcf67e056e02646", x"7445bb3638ae0806", x"803bce7a27a9329d", x"04966ff9230470db", x"58d317d41a3f19c6", x"7ef711cc3b556fd7");
            when 24742361 => data <= (x"3f807ef3a951b65f", x"8d93589a86de3e1a", x"09ff388534e1eaa7", x"dace8fd4b6f3a3a3", x"ef1d43bbd2160268", x"e5cce361b5d460ec", x"657df4d14e3cc4db", x"ef05bb19e605821d");
            when 16836151 => data <= (x"d927c531a04c4c7a", x"881350051e187693", x"dc96dd8819fc3405", x"7bfc7c7c9872be37", x"50c16c990f258d78", x"31244c64850f9a0e", x"bc320b805a737a3b", x"64bf0fb5e2001c80");
            when 15411889 => data <= (x"56b5a4e4664183ce", x"20f54bc35c4a6229", x"55d1d92ad66a0f19", x"32d5bd6fd17b2665", x"1cea46fbe6ff2202", x"93d1356855cc3d13", x"90f189e53b828a00", x"f553b6e8ab609267");
            when 26806388 => data <= (x"edab16974b23a2b4", x"363877a47869be32", x"1726ab497e993504", x"c70069b20ec93887", x"500d6d9833ca73d0", x"d3be225477ff00cd", x"141e3e9bfe72f260", x"2403a6281d8a9a24");
            when 12544892 => data <= (x"e2360607341cd66d", x"d4455ee6b6f2b3df", x"a7cefd9c345fcbe5", x"1b7b89015312a5a8", x"75ada8ddd748695f", x"4fa16043ab36a1a7", x"4afa7110f4cbc4dc", x"b1aaa4c769498b5e");
            when 7433284 => data <= (x"427ab9abc20c8a49", x"dd367fb7940b56cb", x"bc446a15dc7b9dd4", x"eb8f62e7c412ddf0", x"58046e25f6031e7a", x"96a2743c7385bb86", x"c152bdb305645ba1", x"74cbdc13009e0e2e");
            when 10849837 => data <= (x"1c0cb49c7e537d82", x"66e6f7df9b3d140a", x"6390cf679faa5e91", x"37cbdfe48350fa0d", x"7734cd2af0c576b8", x"2743f77bae7e17d8", x"622d497aefb7d737", x"7c5ccaf3c02a3577");
            when 20825739 => data <= (x"a0bd4f7a4b537768", x"f0f64f94b9ca78c3", x"63b0a0b27601e355", x"0ea11e2aa683094f", x"e40d8950dbb49773", x"3eb65889148df362", x"3c69533548bdc846", x"825e2a5fd7f4359d");
            when 8922073 => data <= (x"d00f8a248646e692", x"f10c27bbcfd80f8b", x"da053cea719dd725", x"69174b4cf254341a", x"5e8582087f52eb98", x"d0625f43ffc92fb1", x"372d215d87d79f0b", x"7c7e263c9430b2af");
            when 17728713 => data <= (x"33199da82628d687", x"cc6b59b2e9ccc8bd", x"c85f62067a6ed035", x"23fb70b256af256a", x"918a8e3c44e10b77", x"172f04e2e294f411", x"a31ed6043fc2fdc7", x"1a4fc988828b780c");
            when 10976179 => data <= (x"9bbd87a06bcaee2e", x"3c179d42100b6944", x"711a861d11a34dbc", x"92b9d3f1b7ffe636", x"c20c465209967fe9", x"0e21e2b4ccea01f5", x"90ad01fa7dbc371e", x"a571a5034ce2801f");
            when 4818250 => data <= (x"8ff912bd05fdc167", x"64bda6fc9eea5592", x"298e1ec7156aec59", x"9b142c4512379269", x"be9b25f1cd8b5686", x"27405f760f7e277c", x"30fb341279d1c278", x"fe751f464b83714c");
            when 399642 => data <= (x"6626cbd803f6d77f", x"717cd001919e3d18", x"1951738f04bb1fe1", x"350f497f49c52642", x"7dbbd4e782964552", x"acab973ac971416a", x"23252f560691833a", x"0ff2443c38323c70");
            when 4465486 => data <= (x"0cfab395cb0ca79f", x"4b5e76968cdb75fe", x"b25612c160dd1173", x"006e1fbdedc61eeb", x"bd201cedc6c7bc4e", x"62db83079b35fcb6", x"973ca378f36f0940", x"a6646d33270a82a7");
            when 30557815 => data <= (x"6e346b70780e0bb0", x"dd865445dbf8d777", x"d222b8eea0f36873", x"1f367143f50da3ff", x"5fe96baa04f41ae9", x"d8bfcd5b78169547", x"51c0482d8faf9610", x"68f8faaebd5319b6");
            when 16048707 => data <= (x"d16b69aa308ad5f2", x"ad4fccb7124b509c", x"e1f30578a8a5d690", x"1d559fd2d027dcc2", x"fbd585fbdbb7b018", x"597b5cc6baa9fe62", x"ae2afa511a832ba2", x"0c6f6d1a90c29470");
            when 3011333 => data <= (x"df4ab1dec6f42fe4", x"84a35b2eb0ab71fe", x"287db16ced327485", x"fea717fa214b5ee1", x"8c4c6fb5edb968de", x"6f271294b16848e6", x"7cdfe4aa598961c2", x"11c0bd4b47a06496");
            when 20989632 => data <= (x"7e885f69cd4301db", x"dc2d5c880bb72451", x"db7b710d8141af97", x"5fc931e01731af91", x"a653c394b68c6cba", x"a718de236c29f3d4", x"40ccc5bef383ed7d", x"bd3c4ee49b05177d");
            when 17598218 => data <= (x"d97f7a9f112ac9c0", x"fd66588ab0c16297", x"244b0fa71ec90250", x"ad6c1c61d6960017", x"4ab0830fdeddd326", x"00b3cdd1077809b9", x"9de6f1ad79369e2d", x"87d43e3b07e0345b");
            when 17139383 => data <= (x"e850a13c7c71e7b2", x"7c6eec1864b9ff3b", x"a6eb698976e91676", x"6a3f3cb40794fbee", x"f7690f160eb90fd7", x"4a43a704a351c325", x"9f0b768104311d33", x"c6868cbf8e33f6c7");
            when 22085673 => data <= (x"1fdaffa20689bbef", x"6a11c51ec7ac9dc9", x"92f7fe73283dc371", x"2a70c6504882b1fa", x"568d14260d3c0ea2", x"26c8de12b621f23a", x"8d93580d3d61f84a", x"628d716f14483d79");
            when 21514830 => data <= (x"e7a521cd1f4d488e", x"097047b0888f4cab", x"5c40c91de82350b6", x"42d50decbfe1bbd8", x"b1b816a2d116c222", x"f100d7e5921bc2c7", x"1f67e0ec5ea4ee8a", x"923276bfb57be10a");
            when 11648357 => data <= (x"ed63605974bf4076", x"6ace395b803e26aa", x"71c1192df4198bf9", x"8221280aa05cd41a", x"0ba7d5ed67211864", x"4cf27955038422df", x"f9f3dc4fb66e1f2b", x"7bdde5d8d55eb887");
            when 3463958 => data <= (x"ade24a6d6ae926a1", x"a29f8cf0a99554e6", x"dc045f76fec4cdd4", x"83c1866b49542f7f", x"f43ea33aa64ef9ef", x"d083532e35d59193", x"908352c60f18c6aa", x"6923ed79c0a1bd25");
            when 5536125 => data <= (x"95c8140a9cc5a42f", x"6cab6f403c2b3e62", x"5099a677f2ed7413", x"eb12c957699a5246", x"e4c1eadcea9fac10", x"f2cba5ba742fd220", x"36034da6706cac14", x"d39d8a2c862732b0");
            when 21053738 => data <= (x"87e53ce52293e9f3", x"2fd07c05d0602a16", x"017b8845454c1b00", x"0efb916e7244aba9", x"2bc59d95cc5b3883", x"79e91e7cd9479f46", x"c5a38a8b80135e2b", x"e41cac46651a3375");
            when 22745056 => data <= (x"62bab6af633e57e3", x"cf5f802b07b1bd78", x"94cabcccb261a7cc", x"7bfcb7742518ea84", x"dbb776b89233401b", x"73d2f33f72c2f5c5", x"c070b56c17dbffa6", x"5030f5b8fa2a211c");
            when 3160912 => data <= (x"314529dd2636ef24", x"748af1e80c8a7b3a", x"38a137153ca51c4f", x"dddc2fd7dd7bcda2", x"a9088ddd97f04595", x"7ec827eac98640c8", x"fbfd1287fd78028a", x"eea34e75d4f3b083");
            when 33655204 => data <= (x"56934eae745b5af6", x"942fa5335b074486", x"02fc5a45f4c4a2ec", x"d5f6483e9d05222c", x"b37c266fdb1ce88f", x"747e39c24dfb8f72", x"180149934518845b", x"f5dce8517cc35e60");
            when 25263246 => data <= (x"03a0a55f9241236d", x"03c2afe8387346d8", x"12cd2534d7bb299d", x"9996075f0037245c", x"00cefc3eab1283ae", x"b9be82c78b7f1898", x"fd4f66ffb16f10bc", x"f18ce27d0246f48e");
            when 28570813 => data <= (x"1ea64122df4cf3a8", x"b09eb938eb8941de", x"41b01bed86438832", x"5bfe7d2718e0f9a3", x"a13fd786ed9cb423", x"61aa75f805bb1502", x"fabbd024a44a0501", x"efd2e78da303b0a7");
            when 31438698 => data <= (x"0f0ecb083a18e92e", x"bc36bee2fb248dcd", x"03839cc8f14cd42a", x"618c92aee6962120", x"2494f237b8b29824", x"4a2f91306343c6d5", x"28a8680733da678e", x"14eff1f2e9335092");
            when 32259388 => data <= (x"d0369152f4c8c914", x"ec88450796ccddcb", x"7e772a6ca6f24e55", x"7a926351d8b4a908", x"065b5213ae926e65", x"0b92c433cca332fe", x"108751bdc12bcac4", x"3871b1b6863c9da9");
            when 13363361 => data <= (x"a69ec15ec122c73a", x"53f828a6fc1dc72c", x"d3d2e3da5763d25e", x"c19f3cd3a78dbb46", x"7145b5c0fe2affea", x"e34f90a32cf13bc1", x"26c605f780bb204f", x"42b832d9d29f7430");
            when 13592045 => data <= (x"441ddd167b808c70", x"f65714f57d8595cc", x"ba186b12903810fc", x"91679f51480d2414", x"29e1d82b22110e01", x"676d022abf760635", x"233dcc7627467849", x"6e488f8fc7bfe9c3");
            when 23051613 => data <= (x"a411147a90f98910", x"37288f0b754d0b2d", x"dcdc539c6be3e5ac", x"81467a3706e803be", x"3638c4217d299871", x"1473da3a382afdeb", x"4a760a67909d51a3", x"03c2fa028367a0e7");
            when 9416058 => data <= (x"5643968b894feb6e", x"28805347d8609def", x"65384fd49cc9a19c", x"2e13fd531088ae02", x"2dbb01c3da9ac26a", x"2a6d072d64dd8b5d", x"6dc222680b49c336", x"4a82176e6a3dd17c");
            when 24526343 => data <= (x"699fdef1ae6337b3", x"f424167e5974c9bf", x"f45583aa00fe633a", x"f7cc6077ca71f53f", x"df6a23c3734b51d7", x"ff1fe535a27adf57", x"d5f125fe1a0aba2a", x"e7032e933011290f");
            when 20643344 => data <= (x"267ce3ae884b7a05", x"4b6725c1cb5ee8b3", x"17ba7b55de3e1d4a", x"5192e683aa376e95", x"33e155e10977ac15", x"f9eb76ac1e54c733", x"4914e9055d4c6c8c", x"b79b2415d67c6b39");
            when 32296945 => data <= (x"eb5737cb2be18e9e", x"f9ea6f5e95a6362a", x"34edc5e4a224e5d6", x"42d5c2a536e6b6f9", x"c980ce79abad8ad6", x"7c3ce4433a5e8e77", x"794c7aee8e4efacb", x"84de35e2d86a937e");
            when 12002784 => data <= (x"1338e1c33172121a", x"46ccbf795d59c483", x"a1cec78e16d06e71", x"7e86289a288f88ba", x"f6643a1d3145d8af", x"226a22e09a27177c", x"dc3de3c2537db10f", x"24632c96b4a114c9");
            when 1835876 => data <= (x"deff0e86448b9645", x"f0d3ec56be0fd2f3", x"fcadc8b0bb53d872", x"314929ead0117695", x"d2e6c4aca27511ec", x"49f5c285648b8c12", x"29828537a99c6cba", x"7e87631fef8a7b4a");
            when 22654018 => data <= (x"34b489aaa78af419", x"e76b130f7b6dfbdc", x"36c7d5a96058b1a5", x"c45d77c76974c60e", x"7f8713769b9922d6", x"272ac17e0d996d64", x"08eeb484702952a7", x"7966a3763631e2d2");
            when 20362042 => data <= (x"00e09ed454d19b31", x"7b7267f9ad3b16cf", x"f0b82c13faf5cb10", x"bc6a22a38bc573ed", x"58ac3f7a74dd0781", x"12eefbe16c6b9794", x"2d6df4b8b5de0bb6", x"e15b2f718946db9f");
            when 22718699 => data <= (x"682fdaaf8d110e88", x"b4fed3ca9ba86688", x"0f0cc7420556cb43", x"11e4725e7c309ca6", x"0442a8ca3901c412", x"9607ef432f48a403", x"71e36939ebb4031a", x"f64e0e07319445da");
            when 20136921 => data <= (x"e214f49f286fc8e1", x"7dbd74d692047fde", x"9f1581f8d57d6847", x"0731be53ee349c79", x"696bdc331aff6a7d", x"32ccfb948c6a78a9", x"53c4db4634ef05f5", x"5435387fe13f5994");
            when 18624344 => data <= (x"5f8a4b99bac443cb", x"f7845f564c59bb58", x"3991f931a8636b09", x"ad5b510661969678", x"48ae8d7bdae38d0c", x"9da40a7e1cd8c6cb", x"43a5a61bb8fc8295", x"3b2046f9e1bc2bed");
            when 13227954 => data <= (x"8eed450800e1a2e5", x"4280193968767b54", x"d72e2aa71f3e3757", x"7022b5a601eb9c20", x"7884fce3d9ac3e38", x"d3b916ceaaae9e0e", x"2b3f2a9077184986", x"830391a6d2528e9c");
            when 16960967 => data <= (x"724d6fb4f3f8af2d", x"1afb97044a70c51f", x"25522c17580866cd", x"3066bfb068164faa", x"e608fb24b5accc7f", x"93a7ed25869ef698", x"513c1d57658db4bf", x"a1eabf5fc01abe44");
            when 1339236 => data <= (x"0a32dabe9f8f59de", x"8812b6a7e1217d5e", x"894c51a338024a5e", x"1fa75a0ea9b05d97", x"5c66996411583fa5", x"e6ce05e7d79c7ade", x"a5a6edea041e69fa", x"d7d453dd8dbca16a");
            when 11633661 => data <= (x"dce20e4b8df4fce5", x"2d13c67304299f3d", x"883904991b40bb88", x"fdae427b1358ba90", x"a634a03d42c174e5", x"deab5ff71d7f66a5", x"95e5dc1c6579b06c", x"2cb2e3bba5a12d57");
            when 28725300 => data <= (x"08d94c926127a67b", x"f483c6e525895bb8", x"93d4beb15cd4ef87", x"e11ed7aa6fb96b37", x"593f9a8d7ac2aec4", x"08cd4dc0c0e0b7e5", x"9a0ec6b89aa4b8b1", x"d5796b551c10d7c2");
            when 5514964 => data <= (x"dac69b0acd4e6540", x"ab6436fce09400eb", x"552e9b96fc08e369", x"fff3ad938b37a48c", x"ad3b46208d595284", x"26eda5ccdff44dfa", x"a3d91838ab542d25", x"b2aeb61dbd39f3ab");
            when 20281608 => data <= (x"7052606debabb75a", x"0cc12a3228e2562d", x"795fce759772058d", x"f573108618784969", x"fb484f58c6fc4b0e", x"27834ce53f1ec980", x"9fb46e5f7e3c5e2d", x"724747dce8670a51");
            when 27120886 => data <= (x"aa58a9aa74573cde", x"cd36352b07d2d7df", x"ca689c566cc4b426", x"a98cd1c258b5922d", x"b18280d040d4e193", x"1dfe2f2be727decc", x"5d6412f90715fdc0", x"84e3089efea66637");
            when 24053474 => data <= (x"c0689ff66b8208c2", x"112cb087ce822192", x"09cb1eb8357e34e3", x"a220ef7a8783a581", x"d30ca3d4e81ddae0", x"79d798be3d16d1f3", x"63851208afeff40c", x"b6e92abf368cfeaf");
            when 5420769 => data <= (x"b3a74b56ca6a5d3a", x"fd8be559827b4537", x"fd5acd5c9c438750", x"390e257e17662e89", x"786d0746365362af", x"d914f90d888e3056", x"fd8d14523dbb5a8b", x"f2479602f9c15b38");
            when 859677 => data <= (x"ccc08e511a905603", x"5993b433ef799ea7", x"580bd1e32937aba2", x"fc9c55d29052c1a6", x"03d2d7c354833eb9", x"0746b989357021b1", x"0e6918dbbef008c5", x"efffaa248f7a7e4e");
            when 24687481 => data <= (x"a93c287f3b02f200", x"4d6e257afc908c84", x"ddfff476e3c01242", x"c907616fc61e9575", x"48d991573f892ce8", x"361a1a5d302c7d0c", x"a7df0fda355d8e46", x"1351c5f6a0c4db05");
            when 20357107 => data <= (x"614b1164cf3e42f5", x"bfb2e832a8ef1f9d", x"43a1d219414fefc5", x"556a48dd173035b5", x"090d083518eb0535", x"7576b8dccf7c1c3a", x"92472874914b233e", x"aaa8302df253780f");
            when 3353394 => data <= (x"1bb8901da0a75191", x"f54a840af180bd20", x"9e74876136cb7c98", x"103bd7c003fb44ee", x"2aad834b1dc06583", x"09769e8d6dfd857e", x"47f71b2995de0e84", x"98a764ff90b3a82e");
            when 32842234 => data <= (x"85c372336184dae5", x"0ed5b20c87a75414", x"85be0fbca5131825", x"f9843b010811561c", x"6d09d3fe251d8f79", x"0d4cf62901d942f7", x"89fe9d5e91802b48", x"cb0a8188c2bb424b");
            when 15144426 => data <= (x"3ffb91b7680afd32", x"0fcad8dcf67c7db2", x"4e425228768f1ae0", x"ebb3d20aa7bb3528", x"f2b15bfbe261cc40", x"e49af3466c02da6f", x"fa387881023b6c4e", x"4a0dcf468caee37f");
            when 17795210 => data <= (x"973acbac6d7d2afa", x"9ed5fde1991cbead", x"a0b5bca8bdc31b40", x"85df81c6898dc828", x"cc53de60bcf85cf1", x"3131ffd03becca3d", x"0a235c8c350021ca", x"555f195eb57fc80f");
            when 20736444 => data <= (x"684c4f4427fda135", x"f0be13ee38bb0af4", x"00abc3d208d305dc", x"0b78d902ac2cde0f", x"49f4e7b8513cc13d", x"1ed6261746d5d41f", x"0709c78c7312c497", x"b81095d68fe9428c");
            when 23223941 => data <= (x"c96b96f1699ad080", x"f01ca0d63630de7a", x"998a07cd415fd166", x"180f9021c7c6933e", x"4783a68a22f9ce58", x"5f325c318b465f1b", x"2e9948132631f8df", x"ce2ade64dc0d4fda");
            when 6401540 => data <= (x"2674d7e6084e89da", x"d5585b85d4008cf6", x"574994949bfd4825", x"9da0169bed829d5a", x"4a2be153ba40c6c1", x"6ca73c35245e0b50", x"095b964144040dbd", x"bb040802c3a3b7c4");
            when 26097197 => data <= (x"3dc262963d8f6363", x"13d2d4b5c7f526f9", x"60a842eb34b2e517", x"18fcfe26fcc19cb8", x"93849b0c9b573a40", x"a170890a45aa5d23", x"8afdbd42aed42781", x"fe6303c5028e3629");
            when 19099735 => data <= (x"8158642462963150", x"bc71e15a555f0647", x"232b18d99ac77fb1", x"0d6ab3f447db004f", x"f001624abd0be5b3", x"960cc89be3ec4efd", x"60eac6db18c253eb", x"10d8867283b2a129");
            when 33225675 => data <= (x"e735d8932ed90f23", x"b25aa912462b18ce", x"47b4b3da8b3f0965", x"df3466494aac3926", x"c2b5bc35c81a1ed7", x"a9b1a330933a0138", x"be7ab714cefaddba", x"7e76941f5635239b");
            when 26927935 => data <= (x"099647544cfe970c", x"9482a412a5cb5b5d", x"75a0cb7e51297071", x"74cb0a17a07e2f72", x"8787aaed8c269e2d", x"1ba047d3b81a340b", x"b6fd48c3f3445efa", x"ed8c132534989eda");
            when 28110006 => data <= (x"df84c193df7af7b2", x"1fb8eb7a937499b7", x"2e33df2373c61ee3", x"435c79d71acc5dad", x"2e8cdc94e8ef152f", x"93b03730206973fd", x"f421c6af838ee303", x"4e7b887748f06c93");
            when 33669930 => data <= (x"ac5ad106e77bdbbf", x"af2d7ce6bc37e041", x"e794ae2a8fa61adf", x"59d3f9ea1d3fd804", x"a6a9b61eb295d484", x"7a752ca60a75068c", x"98de8b6c620dfe70", x"e1558b0555d274d8");
            when 23920545 => data <= (x"a3f2ae357572a4be", x"5a8e50550ee80808", x"60c6a6342f15eecb", x"fd5d03fed118487c", x"9e923a4b7685edb0", x"d3fd5acb83210104", x"6831d7f3c43df594", x"a4ad9ae360e78867");
            when 503503 => data <= (x"bce4988b61e78fff", x"a6cbdbc330102edc", x"077e209ebe9cf150", x"caa5d00f8e4f6102", x"9e6406d6dc2307bc", x"dc1535d830cbc3f2", x"9a4a40b844d34058", x"b77ee102eff0168d");
            when 15045164 => data <= (x"433410c3b5f983a9", x"fe5c878f450a2fc7", x"7d472ee0cbe3d8e8", x"399ad5df07a9e1fd", x"b69ac34035e23036", x"bed27e9ea9adb021", x"93609fe4e57f9f3d", x"aa935546c77997cf");
            when 16985594 => data <= (x"fb3099c0937fc440", x"c3e34c0095914211", x"9e83bf271cc14171", x"f1f8a3e721af1c6a", x"a8ed8c75aafb13eb", x"42a8bdb049cc635a", x"a16f9c6877ca999f", x"a4d94eecaf8314f5");
            when 1578751 => data <= (x"8de146dc9068d06c", x"145e78c2c1ecb0ab", x"5315f5e436a991f6", x"0f589e01624b9c81", x"08f6403ef81dec46", x"786302e5d58cc68b", x"91266827ecf0ab34", x"6c0a4c0bc18c871b");
            when 18860380 => data <= (x"98c2b6b94e3a5766", x"638387ddaedd5461", x"945a00a4f6fc7c56", x"808250740ed97a51", x"24070b57bfe109eb", x"c6f5c64e4c1acdf9", x"3e34b7bc81b8ff40", x"3b42a8b6acd6881e");
            when 32064377 => data <= (x"5c13b7c69decd144", x"6d273b4ab3a701c6", x"0aa360f1f051b12e", x"615a1f0165dd84de", x"b93d1f676fdecd4c", x"65422f123f8d811b", x"0bab1fabe17d3999", x"8098100ad6b52139");
            when 31641532 => data <= (x"13d73174ca0a4ab6", x"4f55906eda42613d", x"5be863f250362fc8", x"0a8cd12bfa214474", x"2358443a88d478c2", x"b7141b806bfb0281", x"5cbed5b8c5815f99", x"d2b054dd061d017c");
            when 7311839 => data <= (x"d334f465a1b456b7", x"fb3e4707af94acf5", x"32ffb9fde7d3c49c", x"ae4503cbec8ebfb2", x"59bd7ed3a5c8ad8c", x"9923b2fac95be82b", x"660b4d160403d448", x"8a72dc8a08b5d493");
            when 19362386 => data <= (x"af4cbc2d89e2752d", x"0c3750903ae97692", x"04400965fb562f94", x"d7e645e950322ed6", x"f4c345aef96d371f", x"3ec724be8e1a6230", x"aaf1a46227c11ea2", x"085b8fe3062c925f");
            when 16249463 => data <= (x"1842c84435e5cd2b", x"bfe1d655e0ac73c2", x"89b8f032d0e26860", x"808a6f3d84a543b5", x"f7e7c1d884c2334c", x"f04054bdf73ce75f", x"ede6bc7c7b304f9f", x"c286d368d2d15fb7");
            when 13555927 => data <= (x"ca011be4b7f940ef", x"731e9b1ffcc57881", x"3e670096a3df932e", x"e9dae3859452a0ca", x"48a59c2e029f75f7", x"3527419d997983f6", x"78286da8588b2c62", x"84300d3929e064ea");
            when 8809724 => data <= (x"0808685a271501bf", x"c00b2f4348ec2590", x"4586742f8b35f78f", x"fce124bb5954eeb5", x"b5ade88edbd1d1ef", x"1508e8169ffb9cbf", x"5e677baaf20083a1", x"88d0a843cf6965e9");
            when 22219554 => data <= (x"7a8ada13bf56fe73", x"2ae36ca1a0fb7c0f", x"856adfabfc6e5ad1", x"48ba73b2c87b9f5c", x"75cd99fb46e51386", x"4db0cd588218bfa7", x"79fbef939471e860", x"607b6e4ced68ee4d");
            when 14547059 => data <= (x"4b3fdb69db8840a6", x"ef1c1b6bc318ac13", x"8d5244b0d7dca340", x"53465918d1570fc7", x"74e6fc402deeab4d", x"6bec2e857d2d93c5", x"4230b485ab43f06f", x"8a5d25e4df84af49");
            when 13688711 => data <= (x"be4f994413b6aee5", x"0b8b1839c1146308", x"16e036bb3e868638", x"7a9016f24ba33d0b", x"77b953699a19c214", x"e09ecbb73aeea725", x"f0eb05dfcee310b5", x"8b8ee2a91dee549b");
            when 23562383 => data <= (x"d36489833cf52dec", x"2807a0feda91c54f", x"be214a61af4c145d", x"109762847b88e523", x"53f3cd51f629b6c5", x"f05d553341f2c14c", x"1c5f017c0cb677a9", x"1e1128152dc73635");
            when 17436513 => data <= (x"51bd072324a1214a", x"290e0364a1ad4b70", x"6e9a2e795d2b3cb5", x"c41bd8702d1a21e7", x"14a1a79d0ae2529c", x"b9be03a5cebcea4a", x"f154eb831258a5d1", x"356746198a4c985b");
            when 23608401 => data <= (x"584e26aee543491b", x"01c1678d559f6295", x"060638974d979860", x"dc4191bc44ad6bf9", x"93b5839a06ee82b3", x"80135bfa1bdfe903", x"062cbf3e65a61a34", x"c3ee52b547789205");
            when 17275165 => data <= (x"d554cbecc4b0547c", x"2fc83af4db0c0bfd", x"8297cb87e262f9a2", x"17090cd5b8a8a95e", x"57882fabee3ca6aa", x"c2d376ab8bc8bde2", x"6ba33b8ddaaa339e", x"c2c3244f02d04143");
            when 33196483 => data <= (x"2f1f09d70d35e7c7", x"920c30d95f83adfe", x"1d5f8a5b6a1e3aee", x"02a19996b44dbd33", x"ef596f5065a67879", x"7bd9c7916d9c73ae", x"f40b69e8ef6c1850", x"ab7a8a368a3abad6");
            when 24350509 => data <= (x"352fb2d5f5cd5c88", x"63ffbc7ddd75f9be", x"39cfb57da11858d7", x"0f669bf381cfb5a0", x"e9663a607f033c2a", x"4d50460613a298e0", x"c359a54dd6e76682", x"c3a3910022257b42");
            when 4482145 => data <= (x"2195ff52ae5902a3", x"0d261fc52eb404a1", x"9f516f92cfe32806", x"d13c8e2d06792b85", x"f157e7cf650ecb60", x"9d1205b8b37e2908", x"fd83785869aac20b", x"e62a1c8d64ef0640");
            when 25712098 => data <= (x"d820f1b558e0f118", x"6d1ef4fd33b9d274", x"d5f64e61f8f95d0c", x"c80f7cef6382ea2e", x"832668a3a03420e9", x"9d5d1fca93bde0d8", x"4f13f0d8be746e92", x"b1e962ff33231225");
            when 33174253 => data <= (x"608cb4a56b6b9b7a", x"5e1f9daa8c0f149a", x"35661613d722b590", x"09d3732b1ec31848", x"afb4a47798533f24", x"2a6608e3f0403fcc", x"a0e5c7e2dec3019a", x"c15dd97161f2e18c");
            when 31594720 => data <= (x"68f62422de257903", x"c2af2b8b262ec8f6", x"a2e1f620a4786d32", x"5fa54e3fb6cfafd5", x"184dbc1d1a40599f", x"8dac89bc10630513", x"908eb02a006b940e", x"228ca61eeef71203");
            when 2101106 => data <= (x"0e1b0e6028a50c59", x"640d157fd9a1e4ff", x"409ab13ed55d99cb", x"cd1771c4b1d334c7", x"490b889a23679dd1", x"bb66b93abdc00577", x"e7246570fe287495", x"d24c1d03e87ec623");
            when 32023211 => data <= (x"8fab19ed63fb6d8e", x"e9a7e83534435099", x"d16a99836525365f", x"ccf678f71dd84933", x"6232a7b458643def", x"a854aed2e26611bd", x"dde196e81f4a183f", x"07aa79784603ad1a");
            when 2234093 => data <= (x"8c781a192ee8fd7b", x"984202bc09588feb", x"c4d4a27e9510f40b", x"7d4308d07ce81676", x"d7b60ae49faa4852", x"aa90a331a775023d", x"2c6ef5c1a62c82fc", x"2b16235d018276ea");
            when 3477454 => data <= (x"5d52a9ce0db6c1c8", x"5f6c21a8eba37c7f", x"ba27d65157d96142", x"dc684f41014d6a17", x"ffd28981c3d885d5", x"2ad75e641a78de26", x"91f949284237b967", x"9eb496bad9486e1f");
            when 15011353 => data <= (x"f6855d51b56802db", x"2c92b79a974e5827", x"97e53a7fe2bc7ef3", x"3ed8158d7b7e8bdc", x"aa8305f040c65740", x"09fbd9c9d2d320da", x"247a36a661f7d610", x"b9391da2533fa802");
            when 31621796 => data <= (x"a1f120ccfcd8741e", x"4ca1e727a89fe135", x"efdf15663d1e69be", x"22cb9f5e7e846059", x"c6a5fa719b55e963", x"bb295767e2456dd2", x"ce3f0479b7bd410f", x"9a403db534988f02");
            when 19837404 => data <= (x"804f1573ccf17aa4", x"849b0be92694ce74", x"3fa09573b467a2c2", x"8b23f7b612a2d07a", x"58d2e2fcf895d12c", x"8f526d9b064f769d", x"1a6130830f5e5e04", x"c27ff0b117ba913b");
            when 26919918 => data <= (x"837c2ff2b039d1d0", x"e48536c1419d7ab3", x"34b13ab352b9d6d2", x"c0f4228ed911c2ab", x"2da44e881f15c18f", x"a78a64c96b596b7a", x"7d6d23e87599a39f", x"a760f032ef16e057");
            when 18169554 => data <= (x"391cb5b31a67cea1", x"2679d0a4034613ea", x"7d712be51d8a108e", x"f35b07b4a8b68ea5", x"82aeffb053d40734", x"37191eedd7410302", x"f6ed9b171fdcc52d", x"7de4bd8d4cb85abe");
            when 10527463 => data <= (x"485dbdd84b023854", x"b7f207e00631e8c7", x"4b8c5b7f107d847a", x"49a7cda87fe29f8f", x"f42bb0918b85fe60", x"1359d1495e46674e", x"cfbf0d8ac82ec857", x"d3cbfb622a7d6da3");
            when 22142663 => data <= (x"c37eacb6c4254ed0", x"a28db4bf58be1c06", x"9417bb8afff9ac3e", x"6d51d35e9e54bea6", x"61eb680fa380e387", x"e8d1bce5325cfd66", x"1acc0f7c89c8459f", x"a3e62999c9e057b4");
            when 17202629 => data <= (x"62f61c01576454c6", x"94845f07d27d3298", x"d2a490cfb7e10639", x"4fb4e0884eb55b45", x"24d78d7b3004f717", x"0a95b15fa2a14021", x"2d65499cdf307fec", x"ab117350d1ee9946");
            when 19634577 => data <= (x"fe731ae13f349bac", x"1cdd00202271cd1b", x"c00ed8add9c23681", x"069e989f008ded95", x"8cde27edb383c90c", x"d2b95aaa63c01fe7", x"f44ae6a77370693b", x"be1df913fc42e5dd");
            when 27350728 => data <= (x"d68b4d4ab5c150ef", x"5acbb0fbdc879a38", x"30c631b3b72817b8", x"a47441d81e51fd13", x"c67c27aa5d5d7db9", x"2fbf702d7930c0bb", x"c1396c1e78ef6e8a", x"21f650b2fe4a7b37");
            when 14385522 => data <= (x"9d025667602aa15f", x"a261d754e94f5ed8", x"005830f090fb29fc", x"3c6155337a9d347d", x"14f413c9100a903f", x"d03107a91e08e1ed", x"b1200ffa964b9cf9", x"542dbf2dd5b7c350");
            when 25180887 => data <= (x"f64090eed72cf594", x"bb8495b0a0ed4877", x"0e48629c404d501f", x"ad4b00673417dc26", x"864e0ecd588835ec", x"471d6e843b31bdcc", x"6d1cac9dac0c8973", x"71b6721e2dcec291");
            when 26827029 => data <= (x"291a415445ffeb91", x"fd17186097174398", x"3a3fb87cb7e2edfe", x"b8cebaf9939ae3d9", x"a60c304711a7790d", x"f75abc1f4a01a197", x"0388ca99edb7f8a1", x"82cc0439a25f9994");
            when 27942531 => data <= (x"39119de87431cc60", x"f9c2572171e6fdf0", x"d523bdbb3f0210d1", x"87049b867c333782", x"f420dedc06c284c4", x"144e8f7fd07f55ef", x"8f2cc9b92e6cde09", x"c7e15d9dfa1bfd4b");
            when 7957989 => data <= (x"b6d369f8261bee35", x"5bc79d13e0f45ea6", x"b4fb0b95b1eb4cc9", x"ec3ff8cb98e0d575", x"d25f03d86751b619", x"7b8ef726f1269e40", x"2968e7eb5837b864", x"50260f5f6da38790");
            when 17933410 => data <= (x"534b884383bf04c1", x"dc429c1cf80af52a", x"67944d21d215c746", x"074a8a10aef13830", x"3b3436a0714ec96a", x"e0a67016d50d5b1f", x"666a4962dd5e5a6d", x"810841416f92aead");
            when 13265107 => data <= (x"76bb5fd48e8f3742", x"877a95eddfb67be2", x"bad085478b75e9d2", x"c285d94df75a9d83", x"3712cd869b171e24", x"c536416f16fb5e5b", x"8f85b815455fbca0", x"dcc756d557a10d10");
            when 27104760 => data <= (x"16b7a08fbde85195", x"d9043a0768451399", x"56d5ea84ebb5a29b", x"46edcea53955b89d", x"6b8dbecb806fc6d3", x"d911b947b91a1dc7", x"f7edd271c94e98a6", x"e635cb58533d2842");
            when 29111114 => data <= (x"680070e1042fda12", x"a18915113c78a3f7", x"7dae4fcba1896ec8", x"994645a973d2240a", x"121ee33722ec86d1", x"617f25b51ccff3a0", x"ad0b3d4ee2d447ea", x"ff0a5345f6c028f2");
            when 25273128 => data <= (x"f139c92a67b48ef9", x"930c7520e72c69ba", x"bbba04007b510131", x"f7e9a5b082e3d3ca", x"5a43aba400083f3a", x"19f3c3a4240cea7e", x"c69b4fad9fcc468a", x"29f299120a1ccdd7");
            when 27667497 => data <= (x"cede7a66b0bf1307", x"f5f412b2e04d3f32", x"e4fa3f7059ce71b1", x"6bc3dee147ab6c2c", x"748ece322703ab2d", x"bb707877cc9c2dae", x"0c153077effef634", x"160cc23ed86c984b");
            when 5083918 => data <= (x"29aa71f64c773fa9", x"1df2b29b8faa3b34", x"214fee1401d7a0fc", x"923aea3b79861cfa", x"a1458690386fe08e", x"3111ae85ff796872", x"94011b9ddff71a78", x"db46364314d8dba2");
            when 5216245 => data <= (x"9fb2f88b3f5ba511", x"ec690de0c43db1b4", x"f5d424cfc71e91ba", x"56d0783da342b155", x"b0368f010b2bfe5e", x"0414ee90ebcb5398", x"ea1504c252fa3927", x"4c6e1148b8ca28dd");
            when 3719493 => data <= (x"ef7800dc7327fd80", x"a2593f2686a9c3b6", x"5b61f520ac0d9a8d", x"51a649d205334224", x"534170c2efb7011f", x"2bdbc425aa83f968", x"a87619af72439e47", x"f4a755f44c6e0fc3");
            when 18964605 => data <= (x"d40451fd0a771904", x"e8beb1dfacff2b67", x"fa962a9adeedc855", x"13963fefcba37aea", x"bf8a4465138dda5b", x"2daac707a6050474", x"822ca81d544de054", x"a1fb0c46d44d3bbf");
            when 5331231 => data <= (x"826dcfe195fd93f7", x"45f26c80d8ff38ea", x"ad08fe7f8b4c9989", x"6e02fc882d597217", x"de542a4761101875", x"a7fb8afebbd669f8", x"53da84a80d086a33", x"2b05119764212638");
            when 24351521 => data <= (x"a56b93b3683d6981", x"2048085003495112", x"b2ac339959113219", x"20f43a4dae982b3c", x"d7f02e9632db8f7d", x"ab7b3b15c6793276", x"8c12e0e23726b0ec", x"ffa305f58f205302");
            when 10115425 => data <= (x"dbf660195aeef09b", x"9e3072ab3d2ab9ff", x"57442ad2e29e4961", x"3869f3d010532f4b", x"d5a141640f4723de", x"42f8b92f0738a562", x"6d75ccdbfae30922", x"0eb47d426d991f5c");
            when 6452675 => data <= (x"2cfe483f97a1385b", x"8885c68840b0b27c", x"0a1cb144f822fb71", x"6586370e7046356d", x"797ab0041c5bdb79", x"9b110deedc786b96", x"9f880758971118d8", x"dd6097c6924ae936");
            when 10984835 => data <= (x"dc7ac8b5459ce691", x"d05753297dc19051", x"c311f55ea1a23825", x"e9a9541b049a4769", x"ab3e877fee98cb74", x"7e3dcbdb5c5d4951", x"136e3b12968f8331", x"b2ccedb5d1cf8e91");
            when 22332393 => data <= (x"e72f9aaa81bb1f55", x"5d49f925a2f3d7d2", x"eeea55233fd8f3c4", x"955bf6694dcbbc0e", x"cc572a1388ab62a8", x"34a369f28f0c7bfb", x"ebdd44df00ed8344", x"d6e948e5ce8c4c83");
            when 22859723 => data <= (x"ac31165bff8cbc34", x"f3b68ec0646e9c7d", x"f7264f83a7fc2b13", x"d990abf881e997dc", x"b5c0572e0b40e0bd", x"4cf61e75b3ebbcfc", x"a668f2b5e435ad16", x"ff46c2e6d1d5614a");
            when 33752636 => data <= (x"95065c3b4d2b5328", x"23c62512b978e097", x"60332daf31855935", x"f5b8ceb4bb670a9a", x"906ce68ed2ca03d9", x"9df8f4f8110b2ffb", x"0db7a110796c9322", x"1e6fa4b58fb2114a");
            when 15057614 => data <= (x"01739f82c689070b", x"73f6793f2053f0b6", x"84fc3ec591f98fc3", x"850e5a975d5d72e1", x"f0aefd51bd80d8e2", x"637e0cb3afdd0051", x"756985b182fca26a", x"751ff50c405c137f");
            when 10610846 => data <= (x"4a400affac5a564f", x"4d8244b680e72bf9", x"7cecf54fcb6ed432", x"311ddba69ddf27f1", x"e0cae1f77dc7bd44", x"02bb37f0b0f3a79e", x"a5935b8765f501c1", x"55f25eaed9c68b92");
            when 5150263 => data <= (x"02c231710d27b0a5", x"721ec62e6f5e3bc2", x"90effd5107cbd022", x"05ed945b9fa978c0", x"651f71203ecd5e2e", x"5723a8fd0d81bb8c", x"5ff6b5deea8809d4", x"9c55889e94264470");
            when 3370490 => data <= (x"57b0069f4cb5575b", x"502d948ef7813ef4", x"442fbacd43e839bf", x"03de0e8ad815b2e6", x"7be0fbd0d85065f3", x"1c79a680eddfb64a", x"263d541c64c730c5", x"5a2bd80138bd3e2a");
            when 1783443 => data <= (x"501fe2cc2063f0e9", x"f135bbf2797982c0", x"737c4c05ce1ad93a", x"9174634cd408af52", x"f8f04e872fdfe19d", x"fb827df6c4f35076", x"6d9917fed5bcab70", x"66a45449e91dee80");
            when 14326932 => data <= (x"00bab098590911b5", x"614ba083c2a782de", x"bad18e59c2a37cd0", x"683b15c65b40d069", x"5e77a11ce6eb7ffb", x"52f6faf735b7d878", x"09f31dc1a368ac6a", x"19fdedfa86cc90d0");
            when 26982962 => data <= (x"c5a2ddc5db6cf61e", x"8b30ec4661d1f9c6", x"3a7d28c21198b27f", x"0b7b13cbd549bf9a", x"557bc3ae32d4b702", x"bf48fe42e903c72e", x"31a21e2cf7fdb7ac", x"8d5153e0044a54cf");
            when 30126866 => data <= (x"634b0bed90ba2ef1", x"2218a64548653ef4", x"29e8096f56fde58b", x"3be485375c739b49", x"995a7d8993d1c8e6", x"1d675555af2108c1", x"c86264e9c4138acf", x"c6c88177128f56da");
            when 10882845 => data <= (x"813cb4f934bbd40b", x"f917897a355196eb", x"fd8e65429f2ae74b", x"bd065ae0300a8d9f", x"db312d0f989f5560", x"d66893b54060dc61", x"ea74313032617636", x"dafd199803c19258");
            when 3112696 => data <= (x"9ed1d48b7e36cab8", x"cf8d337cd7723b38", x"7cf8ca0e84484ee5", x"853b8332a1c89178", x"5d840db95416cf96", x"d5bdd321e929d7d2", x"2759a1132e0a365b", x"85b2fed710318b8a");
            when 18716854 => data <= (x"52de34167b9ad718", x"ca16fd1739f1e5c6", x"9aa4789d3e4ae87b", x"857e83a2518e2b2e", x"62741a1f53b4ada4", x"1dfeeef86b5dd4fd", x"787316c1e467f057", x"648428d4b192261a");
            when 30348865 => data <= (x"1a3541823fa0a75a", x"fea317d139f53df7", x"38113effcb1b1acb", x"e6076f6a1ba2f71e", x"090ff2bb2464747f", x"b66f3b608417abdf", x"d0ff1325dfe8b201", x"f40cb4401158fb29");
            when 4589093 => data <= (x"d7fcb0c884fd3021", x"ce5e0bf7a5f85d95", x"d7a544cb6188dbaa", x"d0a31dc4c5a344ef", x"81aab9219f27144b", x"12edbf7348f70caa", x"28a0dd9e843c8480", x"648cfbb67d7707f7");
            when 29868674 => data <= (x"e17b86d7150dcdb4", x"579b764ad22882e4", x"1714c4a6c1017ce8", x"7c27db6ec142569b", x"91a75df2fb9fc51b", x"5247db8afaf282fd", x"b73a8d5acc2eaee3", x"77140b5cb191561e");
            when 31430875 => data <= (x"db4df5b1da1d050c", x"00ee1f7a1b155a47", x"727a3a4fc435b9e9", x"f802099d8a30215b", x"b9cb516239bfe2d0", x"a48221f581cbd02d", x"fd709b3deebede70", x"91b2701becca9faf");
            when 13561834 => data <= (x"57acc486782e6c25", x"5c67295af4b8df55", x"2dba73347e7b908a", x"c042e00b82ea3eb6", x"d1fa1daf064688e0", x"da68cd991d462d04", x"d4dafbecc8c231f1", x"999cec8adc4a2501");
            when 31336479 => data <= (x"c39ed1465ff9a5a6", x"1eaa7e0bcb04332f", x"5ead02adad506d9a", x"29c32e9e8fcb03ed", x"d17b3c600e7fabae", x"424f6e082cb3a720", x"6b3d169e4f7482cf", x"c585cd89e58df3b6");
            when 15924143 => data <= (x"6f1e6c8383e532d1", x"8861a3dd1a44d07d", x"d7ac1f77c8b72f10", x"7328b2d5bb135b5a", x"a769bdfb0c814707", x"897f5f7b09e2d24d", x"30f0640bdd67cafc", x"86fb650affa998ed");
            when 12549374 => data <= (x"dec303feff0a7ae0", x"d3555e46f8ebc019", x"32270035251b289e", x"a9d2488f42333924", x"e516cea394027832", x"808587cc40e2d90a", x"b1b3698c62cff331", x"03a0122ee7dc6c70");
            when 31477867 => data <= (x"1b7731ca9cad09df", x"7c294788a609553d", x"a69e4e4069fb6f19", x"65e3d72b039915cd", x"652345c5d4f32c91", x"7066cc6e4a4d1725", x"ca56f93f13368a3f", x"05c50f44d2000486");
            when 32844907 => data <= (x"bb58d9678bf0e4c5", x"2bfc62bd3660577f", x"adc3648d8355c0d7", x"e412e19769d4a2de", x"d35032c15378146e", x"e3e212e70616583e", x"38b0db9745126871", x"08976f2819d4f21f");
            when 2558601 => data <= (x"f746c47590b44c37", x"c754427654d53f81", x"94a66b57db4d7e52", x"c7021eb3279cb44a", x"7cc81a90e888dafa", x"e43f0bdf08ee3a56", x"edbf5155d8147d75", x"1cc59e4ee36c5104");
            when 30213537 => data <= (x"264e6c4c4950d4ec", x"131287b072951358", x"4199231dc8d36a9c", x"224d121340aa3e77", x"c3cfc5890b9a7b42", x"206fa0c7015d2115", x"6ae124b7557514ba", x"9fa08d69873d2794");
            when 29005865 => data <= (x"657091482360851c", x"9b2ae16c7ca6693c", x"b2734ba79d6e1720", x"6684d24a1cddaa30", x"3d5ad6d690bfd9ad", x"00e8a3dae23d4ba8", x"79dca296f9b65cfe", x"50cf782990ab7602");
            when 8850987 => data <= (x"18493fabe80fbd96", x"e23239631c6478bf", x"b0d53f7231a0ea75", x"ba853f036e0f1831", x"04a32f67ae56a6d1", x"58340874e22a6e47", x"74f4b608d95e5861", x"3b03109a32accc1b");
            when 28290147 => data <= (x"82a5eaf9fd42283c", x"10e3d0268c300736", x"773e5eefadbd7dab", x"110f8858c3a8981d", x"0ae4c9e3a6416b04", x"cbb02f6dc8bf0970", x"eb0009c027725ee7", x"6047496d357c2202");
            when 3770997 => data <= (x"07737016c2a280e7", x"5a6e4e42d996ad1e", x"78f3743667738a84", x"600f1ae461b99650", x"e9f40bd3d077b87a", x"58620d24f534bcc2", x"7fc7af421c42e54e", x"382ddb11928c1818");
            when 3670659 => data <= (x"a37697073b4dce26", x"c77faceac3611fef", x"5f4bcd2854d0f5fb", x"0311d74e88635665", x"b6d7296d1019a975", x"a3983bab68292b08", x"53c9e00a38cc78c4", x"762b73a4677c2a36");
            when 15353521 => data <= (x"9fdf6de51d33599b", x"d953b09b109fda7d", x"3d309a617658ce9a", x"18abf2e3fa368a8a", x"290b178a549c1ca9", x"904a14f7f4a7ad0f", x"feae32c7025e24da", x"b79cd9fe1bd8fefa");
            when 26013827 => data <= (x"8e9c424c3f69e6f6", x"d9e1067140232aed", x"1dfbcccdf25b2e45", x"3a5b949c971fefd2", x"ffed3355ec4ef125", x"a200e745ecd74b43", x"bdf98dd8941b899b", x"d60d5bee2da7008a");
            when 14555716 => data <= (x"de17e4ed5c6040fa", x"e2873557e18e18b6", x"c23fcde72c070124", x"e50acd24abbe861e", x"4d0d638c7d4478d6", x"3a3daa7e162753c2", x"431cbabc5c95e13c", x"eaa2f6fd1c854741");
            when 31537389 => data <= (x"21030afd4f9240a9", x"27da2338c378d19f", x"d1a219e91dcace23", x"87587c29724c27da", x"60132d628e4457eb", x"389da63b77f6f323", x"8925545f3cdb48c1", x"0e1c00d1760b4b99");
            when 6139385 => data <= (x"c31e50a94de7c9cc", x"a5d567f19b14bd29", x"1a5a6f2052b6400d", x"e05b2cafcaa34964", x"0c99aaf63263c4ca", x"d59fc2a6aa68a683", x"a46bfe03a97ea0ef", x"5110e3fbafb22e54");
            when 25064831 => data <= (x"1d06e4edb8ae6176", x"ed39416b6d3ba957", x"380d876bd459dedf", x"e1f23cd7f206f9d6", x"5a91210dbe538f3d", x"e3e15d13e3ff45e7", x"17f94e531a33f014", x"ef0709149327dff8");
            when 23796764 => data <= (x"3e776bd71f72a03f", x"6bf6e7d5bc3cc9b7", x"8468090d0bccdbc7", x"14366bb3819d7b4a", x"cc408ae002a087a8", x"0cda9d2e44e7dcf8", x"4364d8d99c526484", x"15fa80d6850c5079");
            when 16282447 => data <= (x"f6ea61ba9f9f208a", x"926ec09129b0a2ff", x"742ff132b965e7c7", x"50d5b5f072a20e9f", x"682c594577bb86f7", x"4b823f2ae90c953b", x"ccb64f9227e982d4", x"06333b23ad8200e3");
            when 27955102 => data <= (x"fa3418886a3970b3", x"8c5e547e6e4c6258", x"0b6c531ba36428c1", x"ae8ca03ce781b6d0", x"fee815a57754c418", x"d30f4cad8784309e", x"0c0a373e87c2329b", x"c2eff103b1bb3caf");
            when 22641833 => data <= (x"a4522f1018436e69", x"25b97c820f11e092", x"aacb26971c3b45c2", x"4fb36e47131fbbbb", x"fd3becf0285c253b", x"da297707cc194139", x"f7a7ef3b2652330c", x"fe5efb175156db2c");
            when 22816744 => data <= (x"119520e114dcd850", x"b7eb886a4d1102b8", x"332cda7e61203f71", x"aeb1c0faf257e0f6", x"faa263fbbcf377e6", x"d8e9d2b76a98e01d", x"1740aa6fc4583ad5", x"c2abccaaba025416");
            when 15383129 => data <= (x"1e69bf326053f826", x"f39e34850bf2bcca", x"a355c06c834a36c5", x"7597abc719ba3df3", x"e1a2cc81de628e8f", x"89c3c38a23c4bd2f", x"4974745225c97484", x"5cf991b9f3a5e38e");
            when 26737765 => data <= (x"cb977f8ffb9ddf58", x"77af084ce1d33678", x"0fc706f26ffdcf73", x"79456205c038a781", x"8f78fa238547c0c4", x"c508b63507d57f81", x"77a7c423f8514a3e", x"7694f35da777762f");
            when 11040404 => data <= (x"5f40bd5dcec6e4b8", x"db4218820537ea0f", x"6719245fc256af13", x"0ba3024428dc0193", x"996605f986794388", x"1e18facd0313fd53", x"70f01a31818fde4d", x"a73f33430d796012");
            when 16257956 => data <= (x"c94d201c47e73338", x"850a34d02963a222", x"77042e06fa82b598", x"eac20971c5e47dfc", x"bbc93d2a53c12c0a", x"573b50099eaca01c", x"572a276a169510e9", x"6304d70b098c2939");
            when 11984969 => data <= (x"9a277f444667b3fe", x"a5b225c90c1a74f6", x"e9bf6bc7fb069543", x"f4c542cc8888c5f2", x"5b85a4177d106aa8", x"5a406f71ce7ebe0f", x"f03558924030a8cc", x"db0fadbad9954477");
            when 32994772 => data <= (x"e8b1692957e6628a", x"c6993ba630869904", x"f4c3e69fecef8a1f", x"0c61d19b037dbf66", x"32004457e03da730", x"5d4e71c1a698eb90", x"a716667299f8fbd6", x"44716d7e721fccae");
            when 19412676 => data <= (x"5782b285512eb74f", x"0860e6583a12bbee", x"dd3e7a1ea0ae8203", x"2dfd6fdf1ef2a0a9", x"34f45b2df28e3e57", x"f715393f437f9da3", x"d09f7dee8352edc0", x"18663e3114622d2e");
            when 31970888 => data <= (x"db662c2a8b37c999", x"4d1c4bcd70835acc", x"218255718aa2670d", x"ec0f441474add00b", x"675f1b9ece06d68f", x"ac8a2b9097ee4929", x"3d042bfec50b0d83", x"41f07e4f6449b61c");
            when 19748908 => data <= (x"c982945eb8200ddd", x"ec4562e3cc6e550d", x"027c3728716272a3", x"9a7e61f8fa648a69", x"1f5e94d18907d4a7", x"2363c6a7e8f1f28b", x"de2682da0c53c53a", x"ec39d3b7b710fa95");
            when 25978491 => data <= (x"6c183098e03df29c", x"acbaefca5abc04e6", x"7f7178a44b10cf65", x"5e637f558f9dd73b", x"9fff758071e7f5e4", x"2e99ccde97b5042f", x"fdcb8237d1e0b73c", x"9a3c4f6f926b1765");
            when 25984320 => data <= (x"635bd7f807bce0ea", x"1387e5657733218e", x"2297172d91f338a2", x"f929250738cd789f", x"917ec9cda7d6a0cf", x"b544d2b913f58079", x"a4ff5099e2887a97", x"83b2344f7dc210c8");
            when 31667050 => data <= (x"96381d548a049639", x"bbdc8e98e28b9477", x"a3be60970528b03a", x"e70c3acc85e384e9", x"ed574ac57a5a2894", x"5e80d66240d989e8", x"c9a43b80c085fbbe", x"b118f2d6ac769424");
            when 31708322 => data <= (x"2e4a6a322fe08920", x"3ad345a1c8caf51e", x"74e8cb0ebee2ba5e", x"dc1677001b0c28a4", x"df1874092d953769", x"150250840b04f904", x"c8a4a50fc0750381", x"d86df6e473ae7d6d");
            when 30593587 => data <= (x"47f0317e8075152f", x"b005b823c17f6c22", x"a4ce00ad929a92c4", x"17d75aa032b16fbd", x"ee6e957533ddbb9b", x"84459f7069be3d8b", x"f8e86f509c45bd34", x"627e9a912cf92a86");
            when 13261430 => data <= (x"cb86f15e5d7c4f60", x"5384d259b9397859", x"f5ba0b6f2e1c1f0a", x"3b7ec7afe8e1493c", x"8dd383e509ff67c7", x"b88e40326bf39762", x"a0d756bba9baf212", x"25455b99114d8d27");
            when 10320469 => data <= (x"a416aa8d2dac8ed2", x"3fd94128d43ec072", x"7d380c274dba477e", x"7b2a0511d5929c5d", x"d9056af798a32502", x"0ffee5433add2e32", x"101ad3df43c10b7d", x"c7ee48aa388f84b3");
            when 33414646 => data <= (x"a260327d1aceedd1", x"dd89bbff137fa495", x"7401d9bc5e59c9a4", x"93b35979187138c1", x"695d9c266bd797c6", x"3ef05c693a39948d", x"77bc730e177c6255", x"090231b292e85152");
            when 23280979 => data <= (x"57e1904f09495386", x"2f1f5ee579831a71", x"a8cb9f907f3a5ea5", x"0b75b61cb3327ccb", x"8a4b815d90348602", x"212b13273011fa69", x"e656089b0aa6e677", x"54aa3a448c05ab22");
            when 13794619 => data <= (x"efb32c91626aed92", x"7e8995e9712b2589", x"d413f44268e4843f", x"124292509771a26d", x"40a3171281b1f1b4", x"6511b35ab0ba848f", x"77117f940a5d24e3", x"05cc0626851743cc");
            when 10847021 => data <= (x"f1e1b115c00e5fe9", x"ed5b7a740180cb79", x"d79ea164e148e728", x"26c72604111ef74a", x"f242eaa76800d41a", x"1277c893e091cdc5", x"da71aca2f81986cc", x"87ae9a3dac9aa836");
            when 10808781 => data <= (x"127e9c9172a16004", x"0da55d4642f474ea", x"07350ade186f2b56", x"5e30255cdb0714b9", x"e469083beaf31867", x"72b5c1dd891ab823", x"5fb39126abe1a354", x"9c024a8857bed9bd");
            when 4502211 => data <= (x"eb21d2117d7e990c", x"7a6dc7dbd43e7671", x"fa21acb83cdf991f", x"054ca49382556736", x"6f27074122b311ca", x"6485feba5294acdd", x"9da25dd967c15a88", x"401c0e63f2a95717");
            when 2330425 => data <= (x"c7019cbb476fd3e9", x"caa30592acc20213", x"eff01d2d14a6148c", x"4145bcc68eee1230", x"cff6543911215932", x"8639ab50837edfe8", x"1e39c86bc4b60f5d", x"8caa447e4954e3de");
            when 4418045 => data <= (x"4bb03b7fc194d34e", x"bbe9be423be9450f", x"bf3e708e1b97564e", x"dbefffaf21f14d56", x"55c1c1ab4551a2be", x"3ed079bb58137e9b", x"c58a3abcb29ad9a2", x"bbf43d8ec9c7bd34");
            when 13896077 => data <= (x"e8dfd21485798340", x"93551eecaebeea13", x"c54d5882a21d7af1", x"e6eb72b0c9cf342f", x"61b3224be96e16a5", x"0bbf84f8b8819745", x"eb67d4d97a4800dc", x"b8ff9d18c6694820");
            when 15741089 => data <= (x"f2272c51107cc1ad", x"77e56ada306f9058", x"8944b808b615d028", x"a75d71c3d8bb49bc", x"e4039dccd0264858", x"7125075ec0545445", x"34b997d17478156a", x"f8bd4eff2be98b5d");
            when 26996940 => data <= (x"4323b7f1b1982e35", x"270b9236497891d4", x"1284c67d10238296", x"b3b701495dd0ff43", x"90d40c3fbbf92558", x"8b0ee16cdd8500fd", x"8833de3e1e0b2552", x"6e206b4f74487dd0");
            when 21869217 => data <= (x"14896f15267e9643", x"4b4aa566563e1bd3", x"58308e8a50739303", x"3e05ff2431265181", x"885bc3eec20dd112", x"dcd1bab5fa665ea5", x"875ab2e6cb49d1e8", x"057894ecfa4c041e");
            when 2260420 => data <= (x"40fb311de18af3da", x"feb46b29d6ca1bf5", x"959cc43529454898", x"315cdaf4ae558966", x"1e61e6cddcb2a596", x"f7526308e1208cbd", x"e027c45037d569cf", x"753342c543ffb68c");
            when 31706615 => data <= (x"62028d610a209b1c", x"d63541fbf566c62a", x"34c224b5125267c9", x"a03779537607c5b5", x"fd0fa9e9c5d471c5", x"7d3606b8210eb190", x"e58e560ad9396726", x"4812139c242e3bc5");
            when 9738756 => data <= (x"0b6871716951598c", x"9fdf21dbed9bc276", x"cc40932b2932d70d", x"2cb5850d720e1b10", x"325981930bfc5183", x"2cf85decb62d7081", x"7ebd386d57f4b0cb", x"8dd0546bfc1cd869");
            when 33298855 => data <= (x"fdfe5087f1913f97", x"72c5da0f714e493e", x"a09c19f8933dcf40", x"5e249012817d6303", x"59f527b813c09529", x"f6312daa9bfb61d2", x"696cd8910fc5da9b", x"64b9c292263d99e2");
            when 30679441 => data <= (x"e325ceb1b63a76bc", x"baf95ffffb86d74d", x"08e860f44708153b", x"439ae077f99ab52d", x"ceaf4c7878090c2d", x"5f90f6b1e87b4c56", x"c1938f311be2d86a", x"6bdc7ad744424f1a");
            when 13754632 => data <= (x"d96b90d693f6493d", x"9dad19cafc200f90", x"979d10ea27985530", x"433351781519a074", x"abdb08148d2640e1", x"b07415955886f4d7", x"3211495b4e5bb7da", x"de7bc3a47270fa8c");
            when 32554718 => data <= (x"f332b065953fea71", x"4f881de003059f74", x"a93cbac183c530f7", x"81d17bc737aa7da3", x"727f3ad4157bd70d", x"9ccf5cf579b6384c", x"220c5f5723add1cd", x"e1b91e8d1ee9644e");
            when 10933289 => data <= (x"6355d62e0d551d6b", x"00c75061924aee27", x"6845a5d60ad9391b", x"dfe5b6775cbc4c92", x"db9768e745b86c91", x"36925f67cc0604e0", x"793719307e1492a0", x"bb7475d13f3de55e");
            when 8832620 => data <= (x"96a7d597b7e575ee", x"17ab3736650f47e6", x"fa3a60d4d8f6783b", x"a669c74376700b9b", x"b1d7cae8ade037b0", x"fc2aa2ec77e4f000", x"5a488c434c8eab4e", x"b0cb544f169ba69f");
            when 24342815 => data <= (x"53d2479a402f71eb", x"53e6edb4f9e0d65f", x"620a0db562dadba3", x"44aee0d1bed8ea80", x"1f7fb1f9f99c264f", x"5c997858c99cada8", x"5318b43a0533b78f", x"b9c79325032849d3");
            when 7172086 => data <= (x"e68a640b0e60a515", x"6355d333b3811147", x"9ca6133354f799da", x"4db113815c036096", x"90313a928f084936", x"f9553a0165236926", x"375cb0060ddf4e6a", x"7313fc6e43ebe741");
            when 26128860 => data <= (x"fc755f120323e370", x"b8ae3ffbd73f9e6d", x"31d1dfecf5bfff4a", x"6d47da565d78676b", x"0f01c387e3c9587f", x"bbd6d74971c228de", x"f04a68fee62e7861", x"2a7175f1be66ce69");
            when 25867443 => data <= (x"4d5ee14675de7660", x"5568f8b1aadbca7e", x"a5053ee7719501b5", x"e89d30ac26ef5d29", x"c7bcb161ce610bc8", x"1d1314fb6b168213", x"42e04a6edd55f0ac", x"0010135786a9a0f2");
            when 11755940 => data <= (x"6b436982e26dcaec", x"fd77d7722f0c6b22", x"b6552bd3cf8378fe", x"cd789a95f8b17459", x"8f69a41a09693800", x"96403f7c625335e4", x"8bbaac9756bba3ab", x"862d478535d94eac");
            when 13183226 => data <= (x"4db1ae82486218aa", x"80bb545e8635a4a9", x"e457e3ed3cc0bf0a", x"d0482fe5acfd6084", x"f3aec1c4613da0cf", x"2de574431d274cf0", x"d08138317a695db6", x"1fe84ae23b9b3cbf");
            when 17564415 => data <= (x"77612bf62ae65c11", x"e5648a392c90c270", x"cf0c397a4e749307", x"e707149f906e988e", x"07e05507b9b2970a", x"9c34fe434b0cd2d3", x"55e04a4ed46df902", x"c67afc2d0b32bb1b");
            when 18671483 => data <= (x"6ce90dd78d0f82cf", x"14a72a99185b7fb1", x"9574521ab82cdce3", x"5f650d220f109fdb", x"43741f452dec1a23", x"5aec1ebd8ae2e2a0", x"aea660ada2fd8845", x"7019685a847db7c5");
            when 5196556 => data <= (x"a97562d3fd4dc68a", x"1b57cf5f155e522f", x"dd36c055475b27e5", x"42b9d89dfbf69fe1", x"bbeae16e58efe00c", x"4094a72482c77bff", x"31c953448343f4d0", x"74fbbeea66678b92");
            when 5545320 => data <= (x"c1075db217e2dd0c", x"56985340f4058b88", x"c7919418f2f4e0e9", x"5980eab13aa241f0", x"66cb9715ef582807", x"ddf49ac04673f999", x"b5b3a3af9897c848", x"13607309db1230a5");
            when 29741650 => data <= (x"588cf4b96cb961a6", x"6a0cedbf9a369132", x"59876daa51087f3e", x"b9c78d35e46a9bf8", x"f6615d52712e4444", x"39708b124864134a", x"1d076bb565f138cc", x"e02cb0cee9e2d9e0");
            when 20466324 => data <= (x"c692a1b445296a61", x"c02a6f2b29ad6a99", x"79ebb08b1ea45aed", x"7f6a9efcf4ac8773", x"6ce697c100b1698c", x"2ebc4a7f3369c151", x"eb130d80d011309a", x"0ce439d1e55db592");
            when 14724762 => data <= (x"02fcf3205cf6bbc7", x"e7e8bfa23f28eed1", x"8d06a07d1d81c449", x"66c3713358239772", x"adbdad4457bf7475", x"2f9613d8294258b3", x"8bb60a706b066831", x"65440262a91f94a4");
            when 33421409 => data <= (x"c36ffef4d40de845", x"455c1a55e5011dbb", x"96866c7157de0eda", x"063ffe68ac4a7e83", x"338d9af1c91668d8", x"04d72caf42ee3c62", x"9b97280b457a13b5", x"e4a598451a9ec6ea");
            when 5998747 => data <= (x"7a6c8ad1e187ff3c", x"b03bb1424abfeebc", x"dcd24a15dc927ff6", x"e41e8256ee1051ab", x"561d3fb3a4cf54eb", x"8b72249eb43fd846", x"ec41a4db93a527a7", x"662bcbdfb8987345");
            when 27036625 => data <= (x"81e924eee68d1193", x"18644cddbfb28253", x"e4b530e387b8408c", x"da3aa2cf41ed6942", x"226ce48ae5636d54", x"b68e4c0f4936773a", x"a1ddc0786902edd3", x"c94c31b8e0fabfe4");
            when 19819700 => data <= (x"d8eb0360e4773edc", x"2e364894eba9fe2f", x"1d775592fa7e9b68", x"df620f0007a475b6", x"e042bc4bc33e7365", x"266a045115eaec62", x"40afaf4f8fd12c15", x"64d7e79044e899e8");
            when 27892886 => data <= (x"cad4aea7950f003c", x"dab5918ab2c171d2", x"7d4d7dd285a7efcd", x"8f9cc24d951c17e8", x"df3052090d7afe0c", x"784278a543f77f60", x"dec70b98b997ab5c", x"d725fc8d790b77b1");
            when 17921692 => data <= (x"d929083678178b51", x"972ac3452abd4714", x"58b65671acaac3a2", x"ba3447575d5c4fbe", x"f67d1f375fc43761", x"c9aaedab6173cbb7", x"04998e80c66e1e7d", x"84386e943b31d184");
            when 3579382 => data <= (x"c670c56e8b1d3a51", x"d653f50bd875c055", x"74bb916bb9cf0b0c", x"9a275daf3d50cea5", x"9bf82dfb1a612fa9", x"571437c6c19e1466", x"779cc08ff6971478", x"184eea2efa524ef1");
            when 17407250 => data <= (x"6466ccd9c7a5f326", x"452a3a2b1ed0c1db", x"47558ca22b667665", x"3850fd8601659a01", x"7bcb549273951f30", x"e8f0a5ca13160e06", x"51b2cb7ca93a8e77", x"cbb03f9e35224242");
            when 17863336 => data <= (x"a29a866f3789d1d7", x"23d397d2353332ea", x"732b122df38deeb1", x"9a739cf0a4c84507", x"335c34ecaab1f116", x"8b52c2049f590666", x"fd9661cc59843690", x"7d5f1281a746fa0d");
            when 25393867 => data <= (x"7fb71d80464d9149", x"2eb45c7843543d48", x"af98c3c970e7762e", x"07f5df3379746a14", x"d2d7594056ff3013", x"508fb544a2554053", x"9c2e6318014dc5b6", x"c97d0850ee1499c8");
            when 13393174 => data <= (x"b10f9e18179218d4", x"921d1aba37c32a66", x"e28f8f646505ea29", x"0258110dbfe52379", x"3929ba05590a49c8", x"b7cf632ccd7b40d9", x"3df679ea3bd188b3", x"58f8a482537ff212");
            when 15963419 => data <= (x"35d4268e0c74d554", x"1619f99b0fb12bfc", x"df5538eea0d7e00e", x"19c4da3b84b9751e", x"c1bfa0dfa751c032", x"1624104e897298fe", x"a710d47bba5e47a1", x"79475aa1a8629084");
            when 15611463 => data <= (x"177622e55cd9a597", x"a5e0db39fa0e7f17", x"59bd63c8371603b1", x"fdd132f11534be40", x"2a739dae4c2ec07e", x"3342c631bb245850", x"9836ff184e5a6583", x"c3dcbd543e1528da");
            when 28560466 => data <= (x"97d33620a57bd3e5", x"0587395d8907c56a", x"4330821a10ef876b", x"476c5ac83747fbcc", x"f7ab3a645353a8f3", x"c8b097d7076ad4d9", x"c4c108e7e83a3327", x"1a856525a2048a76");
            when 26935801 => data <= (x"418fe4812d5914d3", x"94eb5bc1d6239ef4", x"bf4aa1cba3152825", x"77294e1e8341c95b", x"c24247a9d066880a", x"cffa63f01239d1f1", x"76858c02379ea598", x"6bfddd7499a1da4f");
            when 15755665 => data <= (x"17b9c5171b7ce39e", x"d285bac29a0c3ffc", x"f4156101d3c4c377", x"469471e4fad84907", x"5de0283dda239088", x"f27c363b9f01a80e", x"a596fb8cd4c820ae", x"05e0993d892bb8ec");
            when 3306813 => data <= (x"d83ce65d2fd10b2e", x"c5a1d065c52e1e9e", x"b11a1976635cb438", x"462f5f121825dd88", x"9b51af7c2d1c90ea", x"d1d2572d67ed93b6", x"cf75951b18d47514", x"fae4c7d7c88d63dd");
            when 1618545 => data <= (x"80b0279848cc487b", x"e7a7a28a2dbdf539", x"4fa369536a46749f", x"ca1a577854b1de31", x"edeb5396382c57a1", x"27c45fe970094441", x"ca5c74644001bb6e", x"1800802a3c0cd03d");
            when 11493754 => data <= (x"f7cfc4f052cb70e3", x"7ca03a1a2e00f1e5", x"a094dd8a4dc6899d", x"34bccd4f3e76c189", x"880d761890251c99", x"ae19402c4973c032", x"34759c591a9ef150", x"8a9e22cf7fcbfc23");
            when 15247195 => data <= (x"7dfabd3e58059e3e", x"b0a9188a6abfdac9", x"0b9cacbd9651ba87", x"7617bc0ba5156923", x"677450114b00e690", x"72a47630412f5c7d", x"6ffc227e9baf264a", x"228190c59f65b294");
            when 20247010 => data <= (x"fec1b3cc42fa0ebe", x"017a52652b61b863", x"a4c3b6b65416e624", x"5150b4a989b4a863", x"55d2811c43668ff9", x"ace070dcddd1946b", x"668694d4e14ecaa1", x"11901bbd776dd86a");
            when 12663394 => data <= (x"7daf692fd26ef55e", x"69a974384c915dcf", x"982decaf2274cc68", x"6ba494659eef61d6", x"4f137759ce37d87c", x"ac8590c533899eb3", x"d0cb7dd2dff9981e", x"a4378ba35400342a");
            when 23817156 => data <= (x"dfcd7bae03488780", x"70a1946dce1a9fe1", x"e544eb8e23c2dbb5", x"6be60e5d3448751d", x"fa8a31cdf4ae32ac", x"a570f2f5011be280", x"39872c4c75cdd104", x"64451ce2a6f39321");
            when 4582517 => data <= (x"2ea60a4ce3d70b5a", x"7a80b8a955b470d1", x"e9892fe425576aff", x"bfdca4146688cf3c", x"2f7ddb22cbdef32c", x"94131f7720bc0ff5", x"f0c5db9a03c4da63", x"e301bc4eae28f021");
            when 4084829 => data <= (x"b1a1319a24636418", x"9dece9eefa4ab290", x"16078213f0b86a7c", x"928e1327f0fbe15b", x"192eb25f837452ce", x"b4e0182b5b688036", x"c5feba428d35464f", x"30380a5cffc48cae");
            when 4499979 => data <= (x"a466ad76a8ca491a", x"a6825a6758f515a7", x"706b8e4379bcc163", x"3289bfcabc7940a9", x"7a85b4beb6d70ea6", x"903e7f6e0b81db62", x"32111aa62e754d30", x"0f78f20f84af8fb8");
            when 9862518 => data <= (x"1bc93130d072c152", x"159ee7518fa10b91", x"b240b4fc5eb70e61", x"c96aaa336072a1dc", x"74209d2e04e0cbe0", x"1268e5f73a8f16bb", x"0047135473956d4e", x"5ce85cb15819a975");
            when 20181517 => data <= (x"fb5abe34bf623888", x"65fcfb0cc8c01ec9", x"5e6c8575a719c2ff", x"c79a6ddf70377071", x"fbe4fe7af132089d", x"1e5b2842fc07b188", x"2a012afd0ddded83", x"e01f9c5b48bf733b");
            when 20684715 => data <= (x"5dc5dd9659508a59", x"9325d0c20c5a4194", x"c8aeff33c3c7c266", x"ccda70491fa39881", x"7672b83d719d6b35", x"194c491b79a377a9", x"62e787e8517190e7", x"59162dd38df99d3b");
            when 10276630 => data <= (x"a299e9b16285490b", x"2fe145ce6829bfbe", x"115c2a6564fd35a6", x"1f54be6d6ea34392", x"55670a09c0658224", x"504fcd57e99122d2", x"80d16c3192be7961", x"010a3109ab8db42b");
            when 23104596 => data <= (x"50982da6d0e422a7", x"eb2da6168da8a13d", x"ab36a73feaba54d0", x"a627787015c2ea7b", x"15caca5d8bb1732c", x"f92b2088b4a0e1c6", x"e554798342b315b7", x"4326e522f46bcebe");
            when 2533832 => data <= (x"5cdbd349a44b6cc9", x"42db476b775de349", x"df7033fe5735b8f7", x"bd6b981925ae6b34", x"fd14a0e85a259cb6", x"0cab5380d429a3c1", x"813350e16fd69437", x"c2b85e7562c09ee7");
            when 16483250 => data <= (x"26ba8c1c690b06d6", x"480d116f9e9d9fc5", x"a6cfab0bf43d7e27", x"f1b8ba9710a0d25f", x"113723c4cda48313", x"d1ea6b26a20236ca", x"ec1d7a7670b7c581", x"4dfbbbdd42c14f3b");
            when 27758876 => data <= (x"6cad48d40cfdc23d", x"661f4aff1a7616ef", x"489b8e26edd9937c", x"99db7e78bd862e0d", x"5ca39d8a6965a860", x"818442be86f2daef", x"043c1ede60140d13", x"c42fb83f973b492c");
            when 20673907 => data <= (x"d43629d94949ee92", x"2bbbe7724a4f0ab2", x"e748b47463f8a4ae", x"9211d603c7c9135c", x"d89fddd41a9b2ef2", x"21aca9a024a5f2e0", x"e05dfedb9b44e7dd", x"166c3bf0ebd18c25");
            when 8014457 => data <= (x"77bddf70ed88065d", x"70cf253fbc31bf7b", x"cd30c6f52379b447", x"da051606bed5d83c", x"bbb3b1dc5d726825", x"6fe41673695f44aa", x"737055d0ed591c79", x"398412ad29dcc4fa");
            when 12185597 => data <= (x"c935ab92c33eed65", x"5683af54d45d3bc3", x"b5aa8c36a39d3b81", x"7c85d07a6c5533a6", x"738dee8ef6cfc7fc", x"bf21dcb8de19e2cf", x"961b84e4ea981054", x"47f46b14f30d652f");
            when 33697596 => data <= (x"5359caa8584c4353", x"73407e7c3d3cb76c", x"5afd92c9acf6e324", x"9f1dd762a046a47f", x"6016b318838e8a4a", x"93cf940c2ad2c27d", x"dee0d6ded8901287", x"3b9cec70d23fd07a");
            when 18514490 => data <= (x"4b815be707f6f4c2", x"263fe51f65f16525", x"f642519923b7001f", x"510888ac77c268b2", x"930905dd3979acf0", x"e31856cd8feba15a", x"d0eecc1326fab78d", x"5f7f1fbe861bf834");
            when 18756840 => data <= (x"0f1ca49abaaad49c", x"68f08e260d31a881", x"adf8a739643f5e93", x"9e189a902f08c247", x"cf8e32772cf329b2", x"269dcae1eb088a2e", x"70f3e1843161d285", x"c6908d2465de9d76");
            when 10910950 => data <= (x"a2f33decac6cf788", x"ab15936757f1545f", x"b43b2cdd46ae178e", x"b39b84a4b00e5284", x"72b545017de37da4", x"7a72ec14d3ea864f", x"b78bd83b109690b7", x"90cd260a100db42e");
            when 20879395 => data <= (x"7c2e1a6911406e7a", x"f4c744fa6d2650fc", x"43ab91c840c60160", x"a1bc35e6bd72dbf2", x"b40c682815ca2daa", x"0c3469ed8ac1aaca", x"5b2a8a7b752be670", x"9403edaf0864b063");
            when 21615246 => data <= (x"aa60f7bcb7420164", x"248d1e96d66fd6d6", x"a72c2f231af82b1c", x"4fec45ee9412d3fc", x"73f3314f3b99743f", x"90d95a49003c19b8", x"d7649d4d358e1756", x"fa1c8ae8fb5bab3b");
            when 9351071 => data <= (x"8c7cfb8070975963", x"5f663a0c1863f998", x"23d21199ff7bc3ec", x"f7e53afd35d9bf43", x"33f90abbe6911ef5", x"e5cafeb7436eaceb", x"40a23d593d295a6b", x"a68b1739372fceeb");
            when 8582628 => data <= (x"2704797c56f84de0", x"40dad1b4d2a87217", x"7b14213a37457ce1", x"20f4e0e9a59c446c", x"8537c3947aaa7934", x"1c9dc9d433097dd5", x"56f3ebd75ae9b35f", x"d2272996ebc84121");
            when 5716524 => data <= (x"35976825ae4f5348", x"d8ff23936017ad1e", x"c285c3216e75cbd8", x"06bc4e680dc33b3d", x"433a0e71a27166b2", x"e4408c5b4ba19ce0", x"a9a2a9b53fc97544", x"2d8d7b8bb50cbbb3");
            when 14350073 => data <= (x"1b9b55e4d094d53e", x"e0605975f26b351a", x"98fba07075e2b3fd", x"b0ba54114c1e876c", x"4d676ac3d564f6b1", x"739784ddcb29149a", x"ce1fd92fad78ddba", x"8b3979c5354e17b9");
            when 25264507 => data <= (x"213095370168bad9", x"899f636a780cdc8e", x"5d88b95e76cad9fe", x"bec01fe6914d58ef", x"002acd2e74b191dd", x"65133436a0a807b6", x"fa42f04578d6cb53", x"6f120f89dbb09389");
            when 16082544 => data <= (x"632d1102ed86a4aa", x"ef35282a677c2bf0", x"0192200bbc865a98", x"9105dcc31c65768d", x"861d063f58c420f8", x"8f3b2666b8daf1c1", x"e239050402c0238d", x"7305c3f5b5b131bf");
            when 8770793 => data <= (x"79880608fd0553c8", x"19f361b5d0e074c0", x"1a317dc3f12a872a", x"dc35368b30031edc", x"97349dbea9c74544", x"e51998d95d70fd4d", x"2f3183f79ca4e0f5", x"58c918f8d8e54d6e");
            when 22368368 => data <= (x"1b718ac989f5e6d2", x"9b7584cf3dfc2307", x"39c0c784edde913d", x"b06a75476327260a", x"67abd3fa4e09825b", x"51662633c83eebbf", x"1a6f446d5a50ade8", x"6abe0428b0d8aa79");
            when 2440733 => data <= (x"c82041769af7b76b", x"6d2757bff2fa2ac3", x"65ebaa2a33c88a1a", x"9e9ee2efce085c64", x"b6ab39a59d98cb4f", x"9b755d6be8e81a42", x"ca3ba95f55846ac4", x"745bffc90d64f328");
            when 1255069 => data <= (x"0d4766a82b7ff845", x"f5817d00042df828", x"89f82fa4b32645e4", x"56face216effe7e6", x"1360deb05d64ef2e", x"25ada380201d0405", x"88c1764ae18e2012", x"dcc6a035dc94cd7e");
            when 27847717 => data <= (x"4cecb1dbef0996a6", x"594bfbb49d4e4bed", x"e4b2e9594eeaef4a", x"c6dfd2bf4a486691", x"0d85745c9feee303", x"d143e0ce43a53d89", x"44368d59c5c8ceb5", x"d8188020d06968d2");
            when 21068383 => data <= (x"9cc75ce8ee72b612", x"f40c26f58665387c", x"b481076f05e3ec8d", x"cbff66e0297aa7d7", x"e8a3eb21938d42db", x"e26924fc00dc06e2", x"d748ba058b52ffdb", x"cdfae2d96c5781df");
            when 6153824 => data <= (x"c16580c21877ad64", x"d4261b55408a86dd", x"e8bd4895b4305850", x"d95a48275efc7356", x"fac1782d9f3fa7db", x"472e1ff59030e4ed", x"37f697f165a2dcaf", x"9f79c46a04310117");
            when 25671854 => data <= (x"83044915bc7aacf9", x"ad30afec173a7ea1", x"2e58796a31895ae8", x"f9a313c7196c8a48", x"4a2f9508774c195c", x"1a4bd4acd7da3b4c", x"6e43da62d3b01953", x"72a1318d19f6ceb2");
            when 28695160 => data <= (x"2062187d75a8543b", x"c48f33a036a2c74c", x"5d2ead4fdbe30128", x"c67b372581cff739", x"5e2674939df4b212", x"51aa08f5c174a76f", x"f524fcbbccf2f2ea", x"0cc217e11be117f7");
            when 19627051 => data <= (x"50820ed4e6c25378", x"c2b9e93e7f32c00d", x"bac01c9f851fac2a", x"b6da8d5a51b38416", x"9e343dff09336fbe", x"c3c02db45110b22e", x"ed7d32f9ca8d9c88", x"1a76c9df6bcf3c66");
            when 8860642 => data <= (x"c4478aea0f5969e4", x"b2c5f7db7e0735f8", x"3d416e7e6b08d9a2", x"f44435b4030bc8d3", x"57e24b7b38b99932", x"1fa5e5ef0b5e650e", x"c246559490631779", x"249b740f3f2bc2e6");
            when 499062 => data <= (x"1a425bda249202b1", x"66745869551e1826", x"57f9aba876e2c596", x"bea08d35ad9212d9", x"399c3152a757d5bd", x"ce6c5c5a772c67e1", x"b310edfec0e90775", x"ed9d6f42290119e2");
            when 13482554 => data <= (x"b1f7bcb88602a462", x"46ce0414ffa97cdc", x"15a2ffd71e63c2e2", x"b4f8acb0ce425bc7", x"76a004991adebf13", x"d25f4cde6a640f0f", x"1cc9cd1dbe591ef2", x"cf0b9f23940c3892");
            when 22439064 => data <= (x"cdb8c593902f213d", x"e11c224e4259e7a8", x"260023638dd733b7", x"8a66bee6745385e1", x"9f108532cb0196fc", x"e91b11272c394d87", x"addf82fddb7f22c3", x"4aaed2fc96d14aa2");
            when 13164891 => data <= (x"154e0e4747b22e8d", x"c9ed66bce41d2d25", x"13a442b8355bb14c", x"efa08f4cff631443", x"4c65b14032548b07", x"bc709105dc8c7071", x"669103aa263318a2", x"622eba5abd3653e5");
            when 30487683 => data <= (x"2f5fa8ca70cd1bf4", x"6810af44fd41e9f7", x"09191f1b89532e0c", x"ad0c15adbb4ebbdc", x"228838830f55aed6", x"094d8ee61ec3705c", x"474abcef4589a68a", x"a0aa7adfe56f6f8e");
            when 11363517 => data <= (x"aac0abc2992d2b65", x"cffacb1de6839f2a", x"f24e7fc5a76ffa89", x"cc4dd842175bc38f", x"a64f7aee03d56373", x"3e6c68174aad134a", x"ecc983b83abb9443", x"49d45580d3fadecf");
            when 16347258 => data <= (x"c986b545c91b5894", x"c07be98b3c12d905", x"24a7ea20a0c39a6d", x"e1482a58871921b9", x"e8f1422ba1fdca70", x"05facd5245b38b3c", x"37832bd55a875d6f", x"948523d7ca4f974e");
            when 30933716 => data <= (x"08750fa299b424b0", x"f321bac1fd8db7e0", x"b33c52045c0e124d", x"af55a0cdfa1970f2", x"14c6caeacb159b75", x"991d4bd29a4b66d1", x"9b1f69dcd72e9137", x"ca2e6929e9026de5");
            when 29669546 => data <= (x"9ea9c7f1e60b5a9a", x"f3794be574b5bc76", x"0b7e5a509296b8bf", x"f1a8d8567d6b79e5", x"9fcdb8a250906e28", x"70231513dc3727ed", x"1987c784fb9c4eda", x"1c110f29f1d6b225");
            when 13788454 => data <= (x"c3bf8accd7fefd59", x"3ceda78461c42bf2", x"d1b0f1f2cddd15f5", x"8942efd8a25f2fe8", x"b0143489c872017d", x"cbb5f6c63f1c4390", x"d77c8a240848398a", x"01bbbfda5616fa3f");
            when 5768439 => data <= (x"4916d89cf1c8badb", x"b2752cc2f9c7f507", x"898423755870360a", x"cdbccf5623cfe610", x"24dad9a4779870d0", x"145f0fe7c67702e0", x"4459ab6e7dfcae26", x"eb5c63d57bf0cf67");
            when 30890024 => data <= (x"8da377f5de1b22ed", x"c652481485a00448", x"5fab82a92e0a84b2", x"68ca05a0e66a299d", x"608eaead739d72b5", x"44fbdc0b0cd28edd", x"21098128962a0366", x"9da5905842141f6a");
            when 10792413 => data <= (x"92680a5121a88e9a", x"4c6bd297f4acb4bc", x"441e8626be3f2de7", x"a142dbbd669583fd", x"3c4ee8557eca7d59", x"ac3d7d6d9c34fa05", x"5028efb1401c57b3", x"edf98a1febc00088");
            when 1416828 => data <= (x"9d3a978e6977af03", x"b00007d62d3b834c", x"b6a3c5ccd18517a0", x"6e6b7d94d5cd54a6", x"43a39d46f76537f7", x"cfe2494bceb7a593", x"8c3f0fdb11572afa", x"9baf0d68a65bddb0");
            when 14953067 => data <= (x"c3f80160fa49986d", x"c30389e5ec75efdc", x"b86b95ba6d9c16bc", x"5ca2d878ce10b448", x"c62df91f62d5fae6", x"36b3d1736621fc37", x"163207512aa053bf", x"a147ec53824828bf");
            when 10102048 => data <= (x"06d2893d13d4e35f", x"205b76838e9efd69", x"df9672ca3c2e0326", x"d1aa2c3d21307078", x"84e9e80a4bdb49af", x"bc386463d5d8c716", x"ea83c4646338d268", x"7190e82fe5725dab");
            when 28284330 => data <= (x"ad00311c86d72271", x"daba8c9819be5771", x"036c006b366c150e", x"4c422b5226b31e13", x"ea4496b95c5d6a6a", x"6024cb29d73c5db5", x"000ef48e33a8b10c", x"611f4c66b2b70ea0");
            when 25580524 => data <= (x"d1ca271d8c16b814", x"a22435ae34c78deb", x"b7ce72b33c416b0e", x"5bb50b12909927a2", x"ff13e0e4290fc7aa", x"42204a8499f8eb36", x"d8bbc54a98d8e04d", x"671fa6164279e830");
            when 22105524 => data <= (x"f500c368ee984316", x"c66c424a186d1f58", x"d3ca3a66961437e5", x"f6e23efdd2ae0001", x"900a3925ea33df05", x"893d0d26c783f007", x"9c8557d3aaf15deb", x"61149a2fabe71371");
            when 26025782 => data <= (x"6b0b474f4d707824", x"bc6da1344571d9e0", x"a61a47a301e6a733", x"27c8ae06572a4ad0", x"1a4829fafdb53dd6", x"815ac612e4e28a61", x"f261b9619352da6f", x"aa2dc44e44a0f927");
            when 32711055 => data <= (x"0d410aa4bb351246", x"44e41a15ff55a416", x"02a89cbc91ced5eb", x"1cabac039f12be22", x"c927dba0846abf1a", x"102bfde115be13be", x"9542b2c7c40b924f", x"71497909e87030df");
            when 357539 => data <= (x"005a6fd32d4f8a7b", x"047fa9a5fddfacdc", x"3eb8c1f51a1a4743", x"38675df5416128fe", x"474369aba88bc48e", x"511da64ab9617f64", x"1edee1db232aeba4", x"5843a88102a5b74d");
            when 33553389 => data <= (x"e785d232fc01430c", x"38f43209871cecc5", x"b829192fa289ce7c", x"2636c1f9f9b3520e", x"e77dee22ed001e80", x"413c946d4375004a", x"db777beb7c27ecb1", x"78d1ff1eb531172f");
            when 28301712 => data <= (x"9193f6560709b80c", x"225782dbd74a424d", x"c606e9d188d3dc71", x"fd1f4f81adc4bca1", x"1c56e87d5d1e8e63", x"e7c8959bd6b162b1", x"f663459f97af0828", x"c1478273e8c3b1a1");
            when 371468 => data <= (x"e8eb0034782e0eb4", x"b3f48350a1231da9", x"a350d6fbea79f9ec", x"e5a0074a894df863", x"ebe7657bace223ad", x"4d217319b897c37d", x"91ce8ef1adba82e2", x"40cb640ebe61558c");
            when 27639507 => data <= (x"c8bc23d9339785ed", x"a44254124dcb7162", x"cd6c128905260c2e", x"0648cb63d8f01f1a", x"32161ce5ec83b43f", x"5586dac567f80904", x"00d50d61f969e192", x"e2a1a17ab4acf322");
            when 21686565 => data <= (x"d2bb3d4f54fae14a", x"369ad4105c601746", x"ec7a171b1b1e0325", x"6f3b21677debe61b", x"addffb3863c96ee4", x"7e7b4060d3de776f", x"e205d95dde973c78", x"24a0df908ef20209");
            when 10870307 => data <= (x"011a42083c4e00c5", x"2ea64594670b33b8", x"d89b66667dd28c90", x"1c8250518fda6f9a", x"51f445412fb1aff8", x"5aa09f35f47918c1", x"54afebb2c52b8e26", x"f4a06037eb158faf");
            when 11311539 => data <= (x"0797e11467b62565", x"85b0980bdcc8c888", x"59b8c46c410024e8", x"4cab7bf2a5458b86", x"c009f696130d32b4", x"0a20a9e676fdfe43", x"2cc7c8d3f2051b04", x"40c8f3a67b1c33a3");
            when 33003159 => data <= (x"f7deb4d1a8587c70", x"ba5c83332ea8bf0d", x"e44978cd5faf2c46", x"07b5834783970265", x"492c28c542ab1c61", x"4a3388a1b7e33499", x"924fd746a1ae456d", x"e8b9edd679c438ed");
            when 30530109 => data <= (x"77a9198e7e1802ce", x"b6e50541d5503757", x"63349e770ed6a33a", x"b5abf75bbb4cc10f", x"6706c9117746532f", x"d18be13da07216ea", x"00c3cb5960a31aa3", x"5f0c5eeb2387e5c7");
            when 7729574 => data <= (x"134690a59c752170", x"654cb6cf0b2cce85", x"e6f374170487c0f2", x"2cbe62895d2fe953", x"7515c581a00d9180", x"93236e83dff780d2", x"bdcf124397b9de52", x"1dcf5baf1e78fce0");
            when 7695669 => data <= (x"9adaa405a4fe0a28", x"2f0a4f2d0524dbff", x"581de6cd3c222d99", x"ad6deab5f50e7f3c", x"0e2ce52f473cc4fc", x"5e776896c7297686", x"cbd525c0f14765d0", x"62176b971210fb97");
            when 3051922 => data <= (x"141069783945e455", x"1fe667beb62ba569", x"8d0d4f291efbbadd", x"82b9c57b2391acf8", x"067878d9f24f3171", x"1eed6b02b033820e", x"fe20275402aa1e03", x"f357b453afa0f7ed");
            when 3166129 => data <= (x"d38ed946cabf637d", x"f1bd48e90d24874d", x"19ab0eeecf5d96be", x"c99569ecb25959a5", x"80b9a51c04cea1a6", x"7fb2b7069ad6c3ee", x"b501580b596f8699", x"61237c99f1a35e41");
            when 32116986 => data <= (x"3cd15ab1c370790a", x"823c956a2b86355a", x"05e43263152e803f", x"83e03ee7d16aa6c6", x"ed2584d668b66516", x"19043b4f647d6b1a", x"8c882552e5c428d3", x"720925d92b4c77d1");
            when 19819810 => data <= (x"1e62e8645ab6cc71", x"c77575dc484184b9", x"c0807bcb62d0169c", x"aacfd60d807ced9f", x"4168e88c7ef528a0", x"8b5e1713ce87656d", x"f9b05ed196305e10", x"794e13c588111ba7");
            when 16619228 => data <= (x"8db60b6b475df88c", x"dc3c3923379b0ba5", x"3cc077e78e9f0d58", x"16bd1190d1fc9b07", x"e70c0fd3d3618ef8", x"b56606d73134df56", x"a6f1a78a60dd8b79", x"b731a6bf631865f2");
            when 27330603 => data <= (x"677404bcac3ee41b", x"4a39c837bba959d2", x"c27f781432d5b00a", x"a6792d59caabaa6e", x"4f7a0b3ce7ec6b65", x"615fb01c6a1f32de", x"1a2f45353eda7cd6", x"62c4e1980ef39821");
            when 10093128 => data <= (x"b223941d872ea8f2", x"971c1b9656292de0", x"ef39be746ade0e42", x"cff418a2bd5ea8c7", x"0be3cf2aeb932deb", x"cebf42e1fedb4458", x"3e428299333ed29f", x"657307ed830ca25f");
            when 12731918 => data <= (x"746ea0a258eb215a", x"8a64ce9da4970cb3", x"b938b5f6b778a166", x"5f6a9bb8fea7bc41", x"d7780719a5ab70f6", x"5e95921938e80ff6", x"c508254d2125fdd3", x"707a2934fdf98378");
            when 8152289 => data <= (x"b8d66e3462510244", x"f84eba4003fe8b01", x"4a480f222701a31e", x"48264935aa201c3d", x"f2cd2735fa2a67b0", x"94dd7f3b5f81fdff", x"ac4ab93201fe292a", x"6865ad3a54b9e131");
            when 27016235 => data <= (x"3d4b53d8e2925ae0", x"d5c35fcf4671db61", x"6afb1f8e20386826", x"73df8d34ae20f719", x"f641f5fa6cf4b3b0", x"cea8bf575cc4da31", x"d5d9e57ccc3bc4b3", x"123171b7c459bcb6");
            when 1142334 => data <= (x"687c83d09b178c4a", x"f4b0b53503c31d0d", x"81f3000f1cd9617a", x"c15d1b6a6cb0f41c", x"6d7ca7b15c9c48c0", x"b469d535cede314b", x"db4bf6308c1c9545", x"4613365dd7f9c2a8");
            when 32392637 => data <= (x"e0e7d04467b502fe", x"6764d7a09ba3c4de", x"f57d176521144733", x"7b42870b6785d5b3", x"72c39cb8c9c019c6", x"21c7f82098c2ffca", x"7a284c99458b77dc", x"98e02ddada983387");
            when 30289438 => data <= (x"38809792d2601871", x"f45d3b351efcd57b", x"f87ac3ad06791d5a", x"5e83c4458b8a9c20", x"fa71eb6d2674e0bf", x"bc9047dbb6a430a0", x"d2a0e7a73c80377e", x"7827101f8bc5d186");
            when 8354960 => data <= (x"05a90f84b79cb522", x"01fa157236ad9f4d", x"1a2719ae49415f03", x"dc1b9027d7f44af9", x"8a60ba8414b001a5", x"eb7fbbb194328045", x"fd56820545a4e3dd", x"ccd8573880474688");
            when 26916792 => data <= (x"512b0061f01077ef", x"f4fe32b6cd424143", x"0c7ac8aefc814b7f", x"366ee200354bd0ea", x"d2127b587eb3a580", x"92b7450f13e629e1", x"7579181b86ff4dd2", x"1ded24c1b5115251");
            when 15712880 => data <= (x"55b7608273d8b594", x"84e498a8cd84894b", x"2c3ee35d3239bd3a", x"d80c3fe1e0b9369c", x"02f2ec13c1dfa510", x"b993e4a09517b89b", x"3188ecad4e6f574b", x"2c4ba31a3c19d22c");
            when 15487447 => data <= (x"e837a372be1abdc0", x"4525a13b1d759173", x"01892303185a4c8f", x"5fe0c94a3f58a2a7", x"9ff2d99b55dbfbed", x"f53e8874a7448778", x"17fce393c3bc1150", x"03f9a68a1fa27c1d");
            when 11125807 => data <= (x"9e9632b33fb11932", x"76bbbff52547b5fa", x"365d17bb56fa3374", x"2f2f8e7248d9742e", x"acb0c111f42fc081", x"a683b7df9edfee50", x"730fd4e09dfbdb46", x"2439333cb1d3c227");
            when 19247866 => data <= (x"5398e50580dffb47", x"da938b506cc9e121", x"9c0b20928650a449", x"acafff1ab0dfa293", x"b224965385da6ddc", x"96117ddb4d8d7ca3", x"3ca31e796a1581cd", x"fb88e447922045bb");
            when 5014336 => data <= (x"c02910cefa4fefb5", x"22188079e579f9ef", x"81604d390673ad76", x"70201344d4892915", x"a903bf7f2a4ed72c", x"7f651ae1b8a83d21", x"22dc6edc15d1ad5c", x"24888fef870f946c");
            when 17968679 => data <= (x"a7ddeedea93f2616", x"a57437f235780c2e", x"aa3f2a375863ca00", x"40d5992653811a8d", x"e5e62fb4c0b13e4c", x"406dc3a8de60995d", x"0eddd75192f59021", x"789cb9aa7ca5545c");
            when 28253500 => data <= (x"1ec3daaeb553cdee", x"babb0b4fdf8e9091", x"b53072599c6791ea", x"8f89b728934c2e74", x"088ac36edfc1af29", x"18647bf816c441e4", x"728a08d56fe1b263", x"37cb1a5224968478");
            when 29930068 => data <= (x"16820adab5e6d1ce", x"d3dadc984d74ede6", x"5eb633d568b0dc62", x"913d9f9e33ee6701", x"8a8be02dd01cb060", x"bd9c50a255060398", x"dec2d0d571b85fb6", x"3f2456e77fe76048");
            when 13647418 => data <= (x"f6037fd4c6f8e1d2", x"6e4b323815f3e4e6", x"388e338815e855cd", x"1792fd695f88154d", x"cedd9b15d679f93b", x"4eaa03efbe4d93cb", x"ddfc698d502bb0de", x"cca1d0b845b0a6f9");
            when 761426 => data <= (x"5476763d2a2d73ab", x"1598fa9fe744448b", x"cc6a07a7eb8a879a", x"06d4d1f4fba0678e", x"4f12a1edd62c18b3", x"e4fab2ba83488408", x"c4faee1e0df3951d", x"f350b42da8d1a58c");
            when 15414088 => data <= (x"1c315a49ba7e2c87", x"6cf9b95646674396", x"65d1622846263595", x"44a39e3fde828783", x"622a56ffd7b98a98", x"ef44212974b57803", x"bce25a3de3e3682f", x"01c1471ae9cb3d98");
            when 1824820 => data <= (x"091901f66e294f8c", x"81641ab06573017e", x"93d977a81096d7a1", x"871a2e24349271c9", x"e6ab400de04133dd", x"fc44dd0858b58a21", x"5559286d06cd45f3", x"409705e61518d70b");
            when 26417332 => data <= (x"5384e727efdea7ca", x"dbe625f8facb3162", x"d1ca5542b22f48d4", x"54e96a0d860fb338", x"93bc0d457f987fa0", x"4a8a47bd86c009f1", x"f7e65b53273b59c1", x"b24f31f091aab306");
            when 394607 => data <= (x"39f5862448358e68", x"f17d1b104d7ce0f2", x"4513d85ed5520e9b", x"ceca909d378998ed", x"a4c55bce2fb62940", x"e54c8acf36692f3d", x"808737eb8dbd33f6", x"b84b44032a81ec5b");
            when 15357460 => data <= (x"f1a978e8de298478", x"64d5d483d8feb673", x"0eb43d3beaee451e", x"5d1fbbca51a88e2f", x"7a063b070ed5f3a0", x"996ddc4c0cf2c4b9", x"f602b2e8e459ee39", x"1c2fc19b12002260");
            when 13979505 => data <= (x"ae2e4f8f0f934905", x"9d51ef18d9164699", x"5fab253bf93cffdd", x"c4170e0f5bd2a259", x"4f085ac332a820c8", x"20dd908ae59351c7", x"f0a88c75b34e8ff9", x"dec557d050601c12");
            when 14887976 => data <= (x"e981982746b3c9a7", x"16cade0f7156cc5a", x"813d0ded35019cee", x"f8d2287108441017", x"6ea198563799ee32", x"400eaf17f00755b5", x"0a55947e5b33f713", x"74c42b0bfd80bfea");
            when 33646534 => data <= (x"b78197264dc6f894", x"1a2f46570e324077", x"3febdbb6a2f03d58", x"fd37988b108a850c", x"d60c2e11b9f13219", x"9bde02aa9fc8a1c2", x"2509cd9a03b135d8", x"7fe82fec09590597");
            when 32059870 => data <= (x"9015e60d0607ba15", x"563e2f1a4295cec2", x"67f2d5f22e6521f8", x"352b10dc1ac48b38", x"023cef9fe34231fc", x"8ca88e5409442597", x"5fec9bbccbde6e95", x"92b3797c48554eca");
            when 12298975 => data <= (x"196b86b56ce8b966", x"738d97dcb00e34af", x"6bacf6e8342cd797", x"e6d84d95ccadad22", x"8674f0caedeb1719", x"9457e0039e1e558d", x"5a4712d8730042bb", x"0f74e374fda13072");
            when 17863559 => data <= (x"ca04d64eaa36b112", x"546099e0b9c26d15", x"a394cc094db340e8", x"c026e19d2b265f11", x"649552a96cd13b15", x"853d7722b8fc8b0e", x"eba21f04231c4eef", x"ccaa3844a8690df1");
            when 6416779 => data <= (x"d53ae59d018c9abc", x"35c43d14b5bda3a0", x"b1d9276388fb6b0d", x"a5bcb62a85545a92", x"8349c09c47aa87f4", x"8594f808b6fa64ae", x"f7d02b284d19b9e2", x"f3a0edb4e3e05b30");
            when 25107346 => data <= (x"08642780f9bad437", x"9d65c6272e268b15", x"1fac3096cf7ed39d", x"dd274fc9a803bb9b", x"53c18dc491814993", x"3d4ca68c993b58a3", x"635affe859e9510d", x"7a77fc37cb3d0d2f");
            when 16111360 => data <= (x"3964c33acf52ec55", x"a2129e7c007b16d3", x"7e6bb2d83243a167", x"0f75a4850a618259", x"249063d285c28553", x"d7980bb29d8c0652", x"08aa47256a552fed", x"195ab1bc9c9930e6");
            when 8131708 => data <= (x"21d4d7b991a9017d", x"4e559dec458cafcf", x"59ada275e72134f9", x"3c6a87b03cd4afbb", x"a430f08a12cea4c2", x"ffd9f1dbd9ed40f0", x"2a7b861828f4772f", x"48ed8261f27aceb2");
            when 11966661 => data <= (x"c11b327661eb290a", x"7b04a47cb5f1cd7a", x"f50bcc1c727e2da5", x"a62b02d9859cbb05", x"0cf2f6e9a9aecf29", x"9ce9be5aaff5d957", x"54c5897748b5be7d", x"9d842f4edcae9d09");
            when 6140720 => data <= (x"dc28ef2d88742379", x"f8b6fe0f7fae2ebd", x"56689cc7a36ddde0", x"0414b2b8d227dd5e", x"1af82413381130fa", x"45d189ddf1ca5ea3", x"50832d18246b32b7", x"727ef1df18482d40");
            when 6685859 => data <= (x"d9d46fc9803eac0e", x"d2ca5a42905a41ae", x"74cdd31290e0e894", x"31759e9d7c3b2a7b", x"9170578b7dc67fdd", x"8857f0c43259c7a1", x"99b3dbc218d51440", x"dc325c2d8096ff70");
            when 16142886 => data <= (x"1fc88c6ff5e6017c", x"7e204318ba7b9ae8", x"55e398dd6f288ce2", x"cc9dc79a9852077d", x"e972627f8e93546c", x"c4f392381efa30ef", x"849be06d2ffcd490", x"e024de7f694c2fa0");
            when 24726042 => data <= (x"dea72321f75c4cc4", x"5288ccf207df48c6", x"40fe2dd50a315660", x"be04ef8023ec34d9", x"4a0245af5410dac2", x"007205cab88bdb68", x"25e8da10237463f7", x"882b5f0a72f85390");
            when 33477343 => data <= (x"33e84d5d592b93f6", x"8ae2af3e5ec57f22", x"44000a0f97a4c87f", x"6b6f7eeab0bd9c83", x"a867dcf61b7e46bf", x"00b7c102112b0b68", x"6464ab3e53a3be72", x"4e43e3d53fa8dabf");
            when 1943608 => data <= (x"b4c52c25fb4cbade", x"ec986760bbc0af1c", x"28c424341310b923", x"91eca17dcc01ee62", x"e4a2d0b59ce08cbf", x"0fe6b9c38003dc99", x"1f617a479bc77601", x"96af80f0c8f1ee35");
            when 12224532 => data <= (x"cf42769bbe12a1fd", x"167c23f43f462f59", x"c8677fca50494030", x"b07b6d2c908d59ff", x"af76c3a6a9a42299", x"cc69586da933ae07", x"ad1653329de09b47", x"1ba7191952583c59");
            when 25553529 => data <= (x"6e3764aae97b7d14", x"fa5dc186130f9966", x"e89b0c3176f04f5c", x"48823d1f9405242d", x"5820b8804d03d81b", x"c0d1025a59d748c0", x"fe26dcde7cb75c0f", x"35fdb227546d4bf5");
            when 32586863 => data <= (x"f3b9f622c758aeff", x"31197091b6e4adef", x"b745461b9a1c2337", x"85ca1f18f5af8389", x"13b63be5a973e769", x"257aae7f50a6a2e7", x"4cb28a57d1e3f83c", x"a18df90b4c6e2637");
            when 10343804 => data <= (x"b863ab5b5fa9f388", x"24ea4461a0ae176a", x"b5b1b787ea7b5c1a", x"e946fb6235441b29", x"5932e5c8e8d65ecf", x"150141bfe62d3d32", x"79e648da3be8ebb8", x"41961b0b029d44b9");
            when 669276 => data <= (x"d02aa5d517368f1f", x"427ead9cf01aa607", x"c39f196db8017739", x"149eaadffe22878d", x"bbe1393d3f762d01", x"2ee3c6f63a8987c6", x"e41b0d9658737002", x"f66986f1abd106d8");
            when 24580551 => data <= (x"9671bd3e2a158446", x"969ef8c195e1f867", x"7ee4f8a0b535e708", x"e740100a0bf62c6f", x"b228091787eff072", x"3a24b51cc9e52eab", x"5ff1e071a60f6783", x"bb432bb8723f7ea4");
            when 15940869 => data <= (x"6f7dd8fb9cfaf475", x"57af91b4446dfce8", x"6aee3c77ce1429b4", x"1ad8dac37481a6da", x"cd98b4df68640b8b", x"e8623f57baf2dab2", x"a5c13a5fefafc40a", x"aa43271637e6c862");
            when 8208066 => data <= (x"505d415c2f295c45", x"28eb73ee73750ca1", x"eec18193200322a0", x"70c3bb7b9f657517", x"acf556885a5ace00", x"ecc89bda4cd88581", x"a55990f84391b574", x"c76944fe61a4f772");
            when 32521752 => data <= (x"f7f57cff02967246", x"19d06bd35af1fd2d", x"d8024b8c5820b01c", x"fb6f240a430f485b", x"62572afc8de52365", x"b699fe538e712905", x"981508b2ef0af8b3", x"e451bc60244d9bcc");
            when 21274836 => data <= (x"372282365e63f37f", x"c9690a983233e3e9", x"5826e1ea456a16c8", x"51be49223df8a4aa", x"4149834c199b7a09", x"4e9a7ff42c66b574", x"ed82757a6a78a47e", x"fa3a4560d6226760");
            when 22076976 => data <= (x"7aa7889086b457f5", x"a38ea842ced756e5", x"ccb711bddfc5395d", x"3067dcbb018ad65f", x"862cb2f16697f3f1", x"d3b4c23550c0a069", x"3b16ab2c91d64f71", x"36ccbc6cc8961b2e");
            when 3489855 => data <= (x"6b4583ab0807d520", x"b37e9149ee3e3a67", x"f55911b6b2bf177f", x"2af79094ad374cd9", x"5c35d734a5c73915", x"4bedbdc92e186a5b", x"0ce24295092963fe", x"e26d21f026de7592");
            when 24619781 => data <= (x"73634515d9ec1d6e", x"2357eec2d075508f", x"2d2a142404ae35a0", x"73074361847ad092", x"56eb1eea1fde9dec", x"63970a4ae5fdbe65", x"89f03e6423793607", x"782d0fec3614f02e");
            when 32717899 => data <= (x"f71728b3c566cffc", x"e4e587bb6a7582c3", x"7e4bb86665b0e56c", x"153a427dda707fff", x"7912cc4b12fae187", x"4ccf11f71430f732", x"6bf75042b58273b9", x"baf6613705f76048");
            when 19936705 => data <= (x"b71482051b8410d4", x"9632625ee9d7a54c", x"11ec18d0ee5aa1c0", x"4bcaa92d8d00d85c", x"149a49ec3d1d5c70", x"68caba75d5f22a6e", x"d82f6484424ce4bd", x"8a22d6b17ae6a8e6");
            when 32405909 => data <= (x"839bb1aa13c421ab", x"a0964a4fb9f9246e", x"455c0787f24a4a1f", x"8c89485da8fe90a6", x"ab319585b69b086b", x"bae67201a8430e99", x"7a4f7be1092b90d6", x"e3e34884eb695ca3");
            when 29031103 => data <= (x"2c9a22d96a67e204", x"bd6ea6fe25d2aa00", x"a7210487a0a3af5a", x"b45ce779495e5f4b", x"119f674318066ea1", x"fa61fcdbb302e199", x"684cc6bc0092cfd4", x"f546b4448791ea1e");
            when 366189 => data <= (x"635ff4f8f4c3e3b0", x"cea7dcb2b42f6b24", x"ccd8e328363fc159", x"78b6436e9334ed45", x"33ff6db58b3de49e", x"14284bf58ea8e82a", x"0fbf4137df8082a8", x"717975ddf12a65f9");
            when 31862788 => data <= (x"47cffc64ac272333", x"09599b5503ec9b01", x"e0daf731b3ac5a3d", x"71023b5d47fd43cf", x"cacf7ea963ad4364", x"5b23f3347cd5c9a0", x"d2bd41b8f13a6425", x"b637ec5ef50a923b");
            when 25659307 => data <= (x"9c9d3fd479d40b98", x"9063ba9b8d679884", x"1ca51498a5b02032", x"0efb1a5a06edc974", x"e017acf0b270c25b", x"2038c6d53f8b4dee", x"de1e8c87cdbdd33c", x"a1bf576359f07956");
            when 13355483 => data <= (x"7e378ed44d1ef433", x"caf383fa41d4a8ba", x"7941f0ba93c02954", x"41a11b49aea65b2f", x"f772c1d7e9da5201", x"e275a56990d3cb71", x"5e9636aca042b4e2", x"2c4da21822e0415a");
            when 32722421 => data <= (x"c6e88b5bcfd213c6", x"eab5616e6040af5b", x"ebac115622ee9084", x"6c181d98dd692c85", x"17aeaaf794820780", x"5e9e526b144f7f37", x"ddc5a63fb2190bd6", x"4dd381b1f2d34eac");
            when 22011845 => data <= (x"f129e5f969021bb9", x"cb122c6e6bbbd4f3", x"355a1f934301f743", x"28a1f72d16274726", x"e642846e7fa04217", x"0ec815a59d5c97b3", x"2406d0775c614933", x"1425f1f5a7b98eba");
            when 30954120 => data <= (x"e7ac107034ee9727", x"a3d38806d686947d", x"f2ba86a6080e58bd", x"26093f28f335e04b", x"12b502457314cb64", x"0e9904f610fdce24", x"5f9635778e3366bb", x"f816097740882edd");
            when 28127766 => data <= (x"6264b57bb761356d", x"e2fb4989b9290e05", x"372be2ddf99dce4b", x"6c63d098577b7830", x"4e7539a9dc94d963", x"4fe17d561ccc68ad", x"c331d27238c3f2ba", x"30ad6ef6339d0d01");
            when 23862741 => data <= (x"b7ac0a34b01bfe3d", x"05a011f7a5a8f81d", x"bf02403f7c6d96eb", x"946bdc7a66e9adbf", x"6e367dccde604e7e", x"2daee4c3b43fc95e", x"48237f7e80dcafbf", x"a606ec5b987ce1ef");
            when 6390520 => data <= (x"251000f626bb13b4", x"33357d2d1e146472", x"486d070d7f3a327d", x"2d8eec12f7ad7f3b", x"b089057777efc41e", x"b293b2f55d4cad57", x"757ba895eeda2921", x"8d82ad387ad29fc5");
            when 811287 => data <= (x"4ec3a45d7bbb859f", x"bc4b873bbc552029", x"78f3cc55c6da3e71", x"0b173dcf7a6151ba", x"09e30a63fa6193e0", x"c34264a60a90ba42", x"42880b9dab494607", x"5ef1018dca78819c");
            when 15995585 => data <= (x"8ab5538a110eca26", x"0f4f3090cd5b0371", x"b1fbf54d3b664bbd", x"e531795dece0245c", x"6e8ade5377569469", x"9ba2d4475570f8b4", x"49b61e1cfe7c76a5", x"b9bf3f8ebdd38e8f");
            when 30094659 => data <= (x"217f1d0863675bd0", x"a6bbf189f3ec2dbd", x"e3de149631db9e2d", x"51e7b46ed178786f", x"dedbbb215e8a4b0d", x"c2f9fbf74a7b2841", x"60555846f449b395", x"c9e87dd4be04cde9");
            when 33412224 => data <= (x"e620db85e33e5d3e", x"3b7e95e364b3e626", x"b584f0e587ef4846", x"f0919684f283afc7", x"fe7f63efcba2aeb3", x"298825d8e4773eda", x"ff139e3350ac7a32", x"8bfa275b63eafa1b");
            when 14830831 => data <= (x"f0dc023c43c9adc0", x"b67532a9794bc780", x"50fa945989a08f4e", x"3ed95678d6a09be1", x"06a42e66f5dc2e65", x"4867ee8eacea5712", x"667c1ded7e7faa9a", x"230e1c77e980deac");
            when 14652004 => data <= (x"2b2a294bd65dc282", x"3fa7896b94f18db2", x"3274d00c38792140", x"7b388e9247a99daf", x"aa5581d211c13458", x"40cfc7c7bd41b945", x"81083a851127b272", x"ee2149692df95e66");
            when 6741739 => data <= (x"41b7e53e2770903b", x"4ed67e53a3ba773a", x"a8a35bdcf5e39350", x"a73e5c5194da560c", x"dc8f8a97bee5b88c", x"74339378d71fb428", x"1bc00a608860e7d5", x"83fe85dceb21b9e3");
            when 19820345 => data <= (x"3fd4d2093bf26908", x"7c1ce1a7542e4968", x"d8ce8b56cb7a89db", x"3dcf4f34590a2973", x"677ce1beaf202ebb", x"deffb35ab00e4f7a", x"2705211c6dbf875e", x"733ceb946bf2cf18");
            when 17078654 => data <= (x"2378d98c735abb7b", x"78e2f4ace053f9ea", x"7d318b6b229c4219", x"f2a9e9a014ae7707", x"186a741fdacf460e", x"3d71ae4ccd253fc8", x"aa8f745389eb7737", x"a44b32a15e67ee93");
            when 29263255 => data <= (x"7f8529a7aeedce06", x"475418792abcd58d", x"a5dba656427e4959", x"7a0ee2d56bf8eee0", x"3238b93633312425", x"b84bc9bd27c76f15", x"6fb0c97ff4b1fd77", x"bf22c1554f1595ba");
            when 32919796 => data <= (x"a5340e645f6499ac", x"86f12a6f5ef0411b", x"fc05c3009a0e88d9", x"f4b2380f10adf932", x"db92ef8a59c63c81", x"0bda1059f2eb046f", x"60e88691ec4b4324", x"2c448f27b6585bfd");
            when 28563865 => data <= (x"613dd346e2771800", x"9d53ebd31b74c545", x"91d4fdc9fda15e12", x"a8b18f56af71d917", x"03ff07f039121116", x"8ab976565f5b7abf", x"44798b0430d6885c", x"9af3b8aab90ae427");
            when 22166492 => data <= (x"195261b79afe8f06", x"436abc1e78067825", x"34a2ea5e61b01669", x"474d489ec9751832", x"2203a24601e0dbeb", x"aec7983c881bdd2f", x"2f8bc9148e890d07", x"4e7fce0e012f5c4b");
            when 15134543 => data <= (x"65174d6c673a045a", x"228bffc03e6fe13d", x"342adfa0e3e70b95", x"4247c0e382b2dc13", x"129d04c6dac68d57", x"a51f061b3cee3cef", x"e5e135521c6a1f47", x"7c5b589e5d2e870d");
            when 20498559 => data <= (x"08bafc253be55ac7", x"c004880dcae4e872", x"252aba9dcf638b00", x"7da6476710133b44", x"764c437d14c8097b", x"a49de7bf03dc8131", x"dadbe10261abbe3d", x"7a982be93bb57621");
            when 4076599 => data <= (x"4062a2c0597e781b", x"38b4788d8d0810c5", x"ddcd7512b1d371cb", x"22d98b6d2381afc7", x"e41c69e86c4922ba", x"ba045c87e10d24c6", x"c30c31b9af868573", x"a8f416ffb3e4d1be");
            when 2849265 => data <= (x"be33b9d590385a25", x"e1b04c78c6193b4d", x"6775aa685277e4df", x"745526e6aa1c0902", x"0a25c51b216a681f", x"aa90828b9b2b78cd", x"a976627c35cb9013", x"551eac5e926519c8");
            when 7893018 => data <= (x"626a4f2b31341a67", x"9359aea9c6f6ea9b", x"1683817cac9156c2", x"24e4a13c11939ef2", x"2db1212fb1e6f3b5", x"ceeaa3f5619bb739", x"b410397251cb03ba", x"e7029e140021c342");
            when 18529385 => data <= (x"8d93da0e210930b7", x"124be401ae7e1202", x"c325785f4137bedc", x"679fd1d694470b33", x"8215788fec9295ae", x"01f546cf4c38f6d8", x"267a9d6a2ba9537b", x"ed82b29e5b4c216f");
            when 10198435 => data <= (x"2adcefac44cf7831", x"eb52179767c503c6", x"c43b385adaa4e1a8", x"40f2e481d396ae7d", x"0890d77601b6b6ad", x"0d44f0d4d1dd3f34", x"a311cebf08593baf", x"27cd1bffc44e0500");
            when 27085045 => data <= (x"a98a0e8d8f81e4f5", x"65e797fdc4da8460", x"56e825da8d1a84f4", x"0a3815675ecfda12", x"eddb3bdb239daa44", x"bc5c46a3c243e920", x"0c3997d88dc9e655", x"86f38cb46a30bd25");
            when 22222886 => data <= (x"d5d13cd42a311634", x"a633522939f67bc7", x"c4debe5ed5860bac", x"7363d1308035ac5d", x"496fa8c0d2af4f25", x"e7a7382a6e460b08", x"fa829385d3ada88e", x"6a73975c1248df18");
            when 5751568 => data <= (x"9cadc016cbf6e592", x"7464b42f56392c64", x"10e54573e5ce0f14", x"a72538199c68aac3", x"1412c4e7e25f0dc0", x"72d34a21cd2ad9d8", x"f6d1b190db3a064a", x"dd2ed7dd1e00ae6f");
            when 7609231 => data <= (x"c5c7dc2a7b8a9e6a", x"44af1fc6b19b777e", x"ef5fa9ff11a584e4", x"b53d348a1333f34b", x"b92d382edad52644", x"7dabf51d548ccda7", x"f2dd2f22efaece32", x"0c3952eb292a396e");
            when 2551998 => data <= (x"6d0f90b1e743cac7", x"fac561d4c8330690", x"a9bf1f332658da39", x"e9f05d0d29c7dddc", x"b09cf27e591bd662", x"f670d19f449b28b1", x"b52436d1e8bc8831", x"fbf0298933149036");
            when 7080755 => data <= (x"65f9ded0fb274ac2", x"a7017039ab3a5e20", x"5e96144b96083733", x"00f5c4cee06711e5", x"302a9282ac330c06", x"6a817344425d260e", x"8d698378308f8c94", x"e5a6bf89ed29a888");
            when 5147270 => data <= (x"c3f024738fc8faad", x"e1239e07595984a4", x"a1467472195f975e", x"3f940d710db124fa", x"2c991ef3f7061a1f", x"37116dfd27dd5a53", x"f4464a6e46401999", x"29d918211daa8bf9");
            when 33768253 => data <= (x"64334b8189b179b3", x"ff89d4f7eb89f56a", x"add6137b79174ba6", x"0d1d7227acb06da3", x"3c439bcb23b95268", x"5a54271172ae5acf", x"521cae28ccdb7547", x"f15d16f63ed6c755");
            when 7652908 => data <= (x"73b922753b3a924a", x"ef3f470a4cd987a1", x"94bdd22d8200776b", x"840c7f382f923df4", x"ddb66488051d670c", x"e2cb58f917575039", x"262474325805b918", x"a5776763fb1acd0e");
            when 28554949 => data <= (x"eb35f477c4458743", x"4d0694ad8527362f", x"f8f5fc8a719f8687", x"70513f81da150ca6", x"47b3c90fb818e5bd", x"a44246e4aa204d3c", x"7fbbffb9a6078e48", x"c82809f12666da2b");
            when 1719537 => data <= (x"6672047fe1ec2163", x"4e16093e8906c659", x"599c7532990b1bbe", x"65a50180da61b2f0", x"9f84dc272ba08b0c", x"e016168a3e70ed3c", x"94d561d2261baadf", x"08e2a3fabb976990");
            when 2759589 => data <= (x"88c4e375d6650458", x"bf7a9c3cc5a4159a", x"33b53a299fc12f77", x"0f5c2f9792bc964a", x"9093718444b44021", x"2b73efd34e87bcab", x"0f905bc47520b61d", x"498bfed085e41294");
            when 30270467 => data <= (x"e1f2e587ad3b0b7e", x"9f289293798b866e", x"8aa89bf3d7fc1b66", x"11b540a2816a7c0e", x"8e06075edeb481d4", x"07bab9ee0ddbe886", x"b55c2790de05cc77", x"a2ae469d9b7d8b8b");
            when 10522887 => data <= (x"9592349c4df61aa3", x"095b022a8ec55cf5", x"77d5835bb12a82c6", x"818f47c0b72b9b2b", x"0237ff31ea3dfaa3", x"d1278dc87ab28ef2", x"111b3f759dd068dd", x"fd31bb3616e664ea");
            when 22289683 => data <= (x"eb6e39da81eb0255", x"803fb06e1838bcbe", x"7c07b3729026d008", x"bf3e36c799b62b70", x"ae42e34441143903", x"cda941a2b56bce24", x"05b5342deb906b91", x"eb303f593ad192bd");
            when 16946726 => data <= (x"d0383452c89aacf5", x"570143c1690c338c", x"c529bd7c56f3612d", x"00c2c7f75717d44a", x"994b1cedca96f8d6", x"2092543d47ca4125", x"27781f8ca1c72488", x"9e417b63867d536f");
            when 20909344 => data <= (x"111d44d517dde092", x"3f1eb15e5dcc5f72", x"9a0a4764cfed3690", x"e6955ff3c100b383", x"b4c9e0769a6fb79f", x"48eaa407327b55d3", x"2efa68e69c518524", x"3e77039dd43078e8");
            when 10509681 => data <= (x"24d3bc32817df1cb", x"06cbbd825a8bf92b", x"5b82149a7049d84d", x"5347ee06f996a0ff", x"5df36d2bde2a9e21", x"7c1a59ec5d0631b0", x"2b1a462f79809f20", x"8e27fc341d61d8e3");
            when 6076394 => data <= (x"69a6ffce52735610", x"634c0e11b8d21d52", x"027b9f4664d47168", x"6d4b64e993a09dc4", x"f9268cd6c3c7906e", x"b88dd97ae8ff78d8", x"8d6695409da7f8bd", x"4e7bef40cc2277f8");
            when 26448688 => data <= (x"da05c818202e107e", x"2aba41d0f3edd536", x"f972521aa03fbcfc", x"74b42eac64f9b323", x"085243e3394f1b30", x"e2083b3422ba9abe", x"0e2203c17d92f211", x"1c2d7faef6e60727");
            when 32697736 => data <= (x"ae74210833fc39de", x"b3a274c3060e9413", x"a19d905d5e8290de", x"5fd5ca231007e43a", x"ea49fe778b2096cf", x"c45558a17da40f6d", x"8d4bfdf123a1f399", x"22b83f1b46526e91");
            when 22045292 => data <= (x"341173f328608e21", x"f35bc0d568eaf923", x"36f43ceb3845e4ed", x"91a34b7d4b85c8ef", x"15d9bc0f47899b68", x"cb8070b9299e86f1", x"62518e4dbce75694", x"90cf7b8f94d4a2f4");
            when 31648186 => data <= (x"10e92ec58e414943", x"ea6f5f7c9466a73d", x"b9722507dba7c590", x"45074fbba290a10e", x"dbaebb40b734c706", x"75ea0a1e0f0c94d2", x"5f5d70610defb1aa", x"aa4a7e4411f67fbc");
            when 31604941 => data <= (x"503d993ca79247d4", x"57cae7b0dd516f90", x"3267655fcaaaf09e", x"6937051266f21941", x"aa8cfdd1c73eaf34", x"b70b5b19797ce9ba", x"d0859c579d86501a", x"83676d8e5987a783");
            when 31925009 => data <= (x"7a23f5887e4ed53c", x"7e77c773c748bd85", x"4788b6dfa058541f", x"4da7f5631aa5ce97", x"e7d3de6ad73e4091", x"ff63387e1c32a6af", x"2db306c5b2d4c6cb", x"0157e39e0048a7e2");
            when 13532630 => data <= (x"ad013ea220c75d9f", x"79c284f4d8e71c99", x"fe95de2221c27704", x"32d47cb1fd93f73b", x"4ccc50924da0bdbd", x"a986af3da5e329f3", x"6b1acf93dd968e9f", x"3e8e1a89e8bc024f");
            when 13244882 => data <= (x"a0cf09cc3599c049", x"0acbf14a92b7fca5", x"ed1925e3595199c8", x"4ec0f6e2f09fd341", x"38788b710eeccc7c", x"294adf554a9ef588", x"9602aa26a78acf8f", x"e71ba31cf21e402f");
            when 14986678 => data <= (x"7a3744615d9d22e5", x"8d607205be008994", x"860031f77bfdb945", x"6abca30cfeac272e", x"4b6700395608ac89", x"57e5573116ec65c3", x"decb2db09a92a6c4", x"2276a61312e18262");
            when 32128671 => data <= (x"acd1f0a06d93559b", x"fcca29eb1c03e7c4", x"547af66edf8a887e", x"da7dd3c11e4be63e", x"d698d4fca7422860", x"e1c1fd3637b6cd6e", x"92dfb24a15d653da", x"dedb0648252d66de");
            when 8251055 => data <= (x"db0b08318fbd9ef7", x"78aa85686d9a4a15", x"a787df1defe6a369", x"97686cca8629043f", x"110a487720dada1c", x"4521016c37103d1c", x"1ce24c82da6264c7", x"a855162545dbc477");
            when 30476709 => data <= (x"eb77ec88d6886779", x"8efaa78ffe06a852", x"17198ce20062c65a", x"c08a6472fe7aacef", x"761af18567a49df6", x"61906b07f0fe2608", x"9f2fc85c1ddddaab", x"17ba7ed504b32f50");
            when 24454626 => data <= (x"14b6f37e4226b9d7", x"9fda31ef263bd382", x"b794037efc4fde20", x"d977b6a9b201d904", x"51a398045d181152", x"ae2d47b0f61bb28f", x"023dfec7cc9cca27", x"00291a429d1c39cd");
            when 32964534 => data <= (x"d3552f3f0de13cc9", x"b26a84536834b199", x"95e171b748047dc7", x"5cb8e812f3e8d578", x"27b32921ea2f859c", x"b1260f1e36555b2a", x"793f87b1b0e91c5c", x"cf3cceddad657062");
            when 17580972 => data <= (x"925f50e40dfa44c0", x"e24c612a181b8c7e", x"62e75ce16f86fe55", x"01ff229a4053c72d", x"9742cb0c46bef8f5", x"9a26d5049f174c7d", x"52eb83a0e3aa56ef", x"700091910427d580");
            when 29732127 => data <= (x"93832a6a010b8b31", x"7cf6c8f1d94f603a", x"6b86c22cc146c2f2", x"a08c1fe04094fab5", x"f72d5eff181fdccd", x"6a05726a45d962e3", x"311e79acf5c99b13", x"f164678f2e29dd03");
            when 28008891 => data <= (x"6e4ac1db1a66f2f4", x"16859d61a2827bc8", x"6131445f9a83519a", x"a35dde1fe4c8c70f", x"81f9232ac7c5abb5", x"ce4bfb3c186a0c83", x"13f488a881bdf86b", x"2f8f20071c95d63b");
            when 23221235 => data <= (x"1d7f3232a8d07d6e", x"88b72d175a52ad97", x"2c1ccb37aacaae38", x"65f46b5029f3e2cd", x"0df90c3cb5dc345e", x"65d260a48e51157f", x"c0472578acda0522", x"54bdcc45c8cd257b");
            when 20757557 => data <= (x"d54e4cd318a7d1f2", x"70d42e2ea2f1e18a", x"785afd16d20348e4", x"237857950507aa9d", x"4fe4e0fb3231bb9d", x"b9554af05c206d0b", x"d027123a455f1627", x"8f9cadc563ffbc0f");
            when 4696943 => data <= (x"bc869ff09b732367", x"4bfbcdac1417cbbf", x"ae94cbbfdb98349e", x"cc728fdb4ca82a53", x"ea211513c742b625", x"fbb3f07d16594d49", x"1388975dee8bb572", x"f1e4dab787b7f830");
            when 29539349 => data <= (x"ec963f5befda8ffb", x"d0b656424cf644a5", x"5e72521e151a34dc", x"e6e6f7f1a4817bcb", x"4674e517a3438132", x"b492852296b74c2c", x"c99e6472f48a1644", x"c57066de31d5c3a4");
            when 20918490 => data <= (x"6b4b126d31295125", x"c962aa8601147e76", x"f66e8b1d86a35f46", x"c204248407789447", x"1ddd4b0533c1cc6a", x"1db1385da99b74b8", x"7f324408844c8b5e", x"8487d04974566a89");
            when 14760365 => data <= (x"a33e53b1f34ee85d", x"82aa540409bc3b4d", x"965862f105f999dc", x"823263d8578d8693", x"2cccdd2e50d568c8", x"15341277b592e636", x"5178a5ba95495701", x"0d55fd08a4fccc27");
            when 12758964 => data <= (x"7357e8e2875ae688", x"2c8f54decb8b667a", x"8a50ce0472095c20", x"85c38cf978d7fffa", x"7f501c4729e97291", x"8c78d0c78aecae33", x"9b7d88f5a2d153e4", x"6853d7a65d88b2d9");
            when 910873 => data <= (x"885de1a572ebe98f", x"a13cf763aa8e9975", x"6380796d868618c8", x"4b2eaa6384e2c348", x"6e5e982309b55a55", x"f00c9f2f6fbe812e", x"366483eb7e3ca7f7", x"918b8db78e3ef64f");
            when 20907980 => data <= (x"5b9f08d9f443c34f", x"c9aad697b1ecd135", x"6b3d21bb3657fc30", x"764002910c0a36fe", x"658adb166e96a2d3", x"67dd91b1133c37c6", x"7b09bd0f3dc596e0", x"2c6e4cbb5779c9d5");
            when 7843411 => data <= (x"f8b404c3e549c2f4", x"76fbf98ea5b53f22", x"5d6572f18fb18cbb", x"85b1a2684b47d363", x"608fabb34a1675c6", x"6701b73275aa836b", x"5489a70e93bc92a0", x"276c55f4a5646577");
            when 8252609 => data <= (x"a47d06ec309c96d0", x"0202435e5b9844a5", x"71328d51b315f826", x"29db58159821d2f1", x"f3b1c9f06b5773d5", x"3231f544f0f95aa6", x"7afec14d4a3a35f5", x"9b906fdc614dadd5");
            when 32833669 => data <= (x"dd2dbae0e9aaaacd", x"32f31d32116c8d89", x"132d3c4cd933b49c", x"0881dbbe59c0ec55", x"bf640cb17d702b31", x"fc8594b790702df3", x"27ddee75ae504c90", x"c6385b90cca904b8");
            when 3061408 => data <= (x"da64f88257a51c63", x"bd3c6633eb9907a5", x"4ec3cc816534f6c7", x"a4061d2ead626d69", x"44a3bb42c2b043ce", x"655e23343b700a64", x"66964029945d60af", x"1704d8dbc978b8e2");
            when 20642731 => data <= (x"e892f58a630cf41e", x"0e7ee11f1ba0d9d6", x"1bf051a2baf3b0a3", x"1cc0d649f9ce315f", x"1cc8d0b236d3c715", x"c5c6da40523fba22", x"18d8a8dddcc18d9d", x"3b7b3ce169c97e3c");
            when 21417883 => data <= (x"10223186e880780a", x"9670ed2d7e2c5b1f", x"325d523e2c51de5c", x"0ef5c47922179495", x"72671f3db9b8caad", x"b338a72715e9a313", x"edb5660396d3c6d8", x"2ae2308dd74bacef");
            when 10891595 => data <= (x"a436dcfff0063be1", x"661d767d57f7c438", x"307e00866508c996", x"e17559810b325562", x"52f76c7e5f1366d9", x"b5de239ed2611ff2", x"5d3f480c23ca3224", x"f2302e2970ccb43d");
            when 7415408 => data <= (x"174399c8c0382c7b", x"6e0c4771433ec02a", x"74aab9e5e595e72f", x"fd2a002a25178666", x"a97bdbd5efa6a564", x"a061f405235e096c", x"b18eac82704aa5f1", x"e6840f3393bf9931");
            when 24711261 => data <= (x"d8b241d6ba016eaa", x"9904a210cb520813", x"b277797b9df27fec", x"7c5a79ad66e36c88", x"4825089a6121e53a", x"f44bf86b11127304", x"1973c97d99cdd04f", x"b0d293aa8e69e8bc");
            when 31626855 => data <= (x"59b36509c212dfaf", x"74b29451affb2353", x"882fa5af6e86a190", x"89c8fd81a794f17f", x"1572b28766328ae3", x"a7e823afe705899a", x"de9b632b880032b0", x"147bb78adf16f1bf");
            when 2336116 => data <= (x"35c9aed90001ee6b", x"44843b743a3468b5", x"ab065037b1fa4d1a", x"78c9cd94a9d78201", x"ac5ad8cca2722abb", x"c0bb971f14ea8c5e", x"fa768b9ffad78a86", x"fbf5ed4b672a973c");
            when 21868964 => data <= (x"b28bf3025da191eb", x"1c7229680495b9ed", x"c13d4c88c15aba47", x"e8e357dc92c475ed", x"7ab55351cb26cb03", x"a5898de628fcf11b", x"331c0075035e15f2", x"3e291f4544ee26d1");
            when 22220815 => data <= (x"fc976e856d3dbc9f", x"52e8fb70b39bdcba", x"85860a3e438977a5", x"c0e7fe3766dc127e", x"abd58f4bc3bf0fce", x"21ec7ae7c452bed5", x"7c502c09932640b5", x"bf2834643f5e037e");
            when 25187565 => data <= (x"0034b7879bc81870", x"a1775cd436940bf6", x"f987fd5162a851f3", x"b0dbbc2abed2f32d", x"3cdbaec5a4a136f4", x"2911e4b59bc146ba", x"ffa6c854d543b71c", x"a3aafeb94e19e91a");
            when 32085612 => data <= (x"9c7096dc18f04ae3", x"c1878fb9f15672d1", x"1128d7a6f4dd89c3", x"ce5177989311de94", x"9e48ecb147a33bc4", x"d53601f98afdc85c", x"f49cf9ab6e2cb609", x"8c26cbd586ab399c");
            when 25790767 => data <= (x"8d20c22029438c45", x"34767de9d21fb2c6", x"ce790d7f04d5f460", x"0dfb5daab0a087e6", x"b21acc7657645a8d", x"1bfeb14073649c47", x"5fb643059fb8a063", x"659b7e7a75bd6115");
            when 7231820 => data <= (x"0daf8b3757d6c466", x"3140ceac87d9916d", x"b06922a55a81b90f", x"aab7a04bb4f57bf6", x"97206f56cb03871f", x"6aa6da1e632574b4", x"77c69842ad398011", x"a299da1a15df0e9e");
            when 18862166 => data <= (x"16d7b4e11cdd23f4", x"78902c8ff5c765c8", x"72a052ec3e9ebce6", x"11944821b873fbe8", x"187263b69dd84301", x"8632e597bf50ef4f", x"dcf458acce71b553", x"40a9e4f5b9c077d5");
            when 10931111 => data <= (x"531e739f539ac27b", x"f35e81dafe3d58b4", x"7a5ee393b953b7b6", x"f97150851b069cbf", x"5c0a5c49b17e7705", x"bce58356418ddc48", x"55a91b1c7a9249c2", x"f6af3a0b5859f851");
            when 12734116 => data <= (x"49f158ea3a8784fc", x"575260dafb1b7f99", x"d2c8099c3fe361e5", x"68a4be4cfa7f68b9", x"63d17270ea57deb7", x"822a1d9f33161be4", x"43e8a392c2ba02b7", x"ad1ebe6cd2808dcf");
            when 14914969 => data <= (x"3beeaf4c19cb99a7", x"6261a29e370ffbf1", x"9898368fbacc2ce2", x"315a1905f8ab3fff", x"46c61726a4033f70", x"c599793f88a2a8bf", x"71fd3ce44ba0091f", x"7438a3d76911261f");
            when 18061069 => data <= (x"7c90d32d4fd4d749", x"e80162e62d73a29a", x"6cf492747946de30", x"a6f54ff335759998", x"90b53f2e45ff2a20", x"4c6ffde2a5fb1e97", x"97db19858c4d9617", x"fe801601da4bee1f");
            when 14936603 => data <= (x"d39b61cfb094d6e0", x"d8306f627e15319e", x"8d3e054c4651b5cd", x"814630059414405d", x"d98727a751a560d0", x"6bf022a964da249e", x"f595f65577c57a11", x"0374372fc2810511");
            when 22530803 => data <= (x"ea02bedfea135c70", x"c37b72f78b034b29", x"1e55863f5aee8b3c", x"cb92fb486f830dd8", x"432fd2c24d3e26b3", x"aed6d02cddc6a881", x"0ea0118d468041d0", x"8befdae9face7457");
            when 14721494 => data <= (x"80626539a9b6205e", x"2d7f8e67a397ab79", x"f74cba8a50afe481", x"314a130e7762ea86", x"985598c4aaa72396", x"348487c90f5d44b1", x"f75bf66a7e04544b", x"54e0eba92198d046");
            when 10052632 => data <= (x"3a1f63c7d379f39a", x"47cf012be1465014", x"d1fcc3d9f8c9ca83", x"f9b840548f08e204", x"f8ff56837b6d14ad", x"12624f52e4e78bca", x"7f15bff550d8447f", x"f9103239af19aac9");
            when 32817487 => data <= (x"3512094f9a22a378", x"54798e2034a1ea0f", x"26c0d8782b0d57fc", x"45c9e85cdeb947e4", x"75078f060dfaad9e", x"a0cc671a5c3905ba", x"e01c621ebd380fb5", x"9f1c6f7ea5ee5c6d");
            when 686915 => data <= (x"995128ec1aa91fbe", x"5a2285bacb4f23a1", x"63578361a05a0cf0", x"5ca3e9690c83729b", x"bd67d382850c7915", x"883b74a38ad1bbfa", x"afbb09794b6e5c91", x"e48ba977150ee080");
            when 24056753 => data <= (x"6efd3c4615a897f2", x"a3d50d37a192c3ce", x"9ad1c087bcde38c5", x"e6b06ff55951df10", x"6d43212d7b99f013", x"f181c1ce8cf214ff", x"42ff74a790b822f4", x"4204e108e6563353");
            when 20673527 => data <= (x"b58e5897b4cfcf92", x"3114198420b53f13", x"89847a0d2840d472", x"21ca8ead3ab34125", x"c8cc978c926b70fa", x"7e0556420191c27a", x"73c17f146cabd80c", x"ad333176b2d1dff4");
            when 15698296 => data <= (x"70f4a601c1ce96ec", x"33ab6cad00ec2f0e", x"658bb66dd585b793", x"4e4ebe2a0bbe7e27", x"0c28e4d25ee2686e", x"69e945e82fc5102e", x"fe1c659037efd075", x"15e03f9f6b7ab7bd");
            when 16395501 => data <= (x"68308dffecfbb46a", x"0aabca6e1b1ce4f3", x"2d8bfa8f76db75c0", x"04893efbcf6b6a83", x"509b160d9009ad8f", x"d94a318f20b45dce", x"260d73f8ac1bff03", x"eea3d4c7133b3f80");
            when 12508455 => data <= (x"d22b5062194d9aa1", x"1cdd508a99edf229", x"50a2e78e8da28053", x"5eb0b655a43bacc5", x"4e251fd5832f497a", x"41acbe1c6f3656dd", x"6096650e102552c4", x"2edf47ded30861ab");
            when 15638622 => data <= (x"60db9b12112f5a9a", x"3874bc93bd9b41c3", x"35011fdad6895856", x"cb3fd35e28004b3b", x"7fd032f079b25d14", x"bd5cb953125ea284", x"149aa3beda168b78", x"7e6cb9cc00e6e5ad");
            when 23579174 => data <= (x"dcbd33ab9f614c6e", x"6b99cd84be360744", x"78fc303a72f77a5a", x"51414194b82a1aa2", x"d6b9631dfdc5b2c3", x"59d10a1a5e6833d4", x"d75132e00a3c8ec9", x"7445c202334b42ba");
            when 31174616 => data <= (x"5311532af99ef515", x"3041eb83ca66cb20", x"9192f307f863a1a1", x"5aa73cef59d17ac3", x"486f08c1c1fa93ac", x"c8084a210e2a908a", x"def174e5ea53afbc", x"b04abee6174a5cc0");
            when 15556237 => data <= (x"cd81980be52931c3", x"bfe9311a93538d40", x"5376d9d67260661e", x"16bc2b44bb5a994e", x"2c2f32a5775a87b6", x"88d9ad6ec47bfeda", x"033c0e034262b947", x"18f484bac3dc1a4c");
            when 5371483 => data <= (x"e444eb9437b917cd", x"d44ca10a3a5cc838", x"befb38752f255b22", x"52cd3c4e85a00f7c", x"ab0646b3394d1519", x"bb58591124eb6f6b", x"44eb68e07885658e", x"fb81fab73f908b74");
            when 10959018 => data <= (x"b01897bd2d2323f2", x"a62b6a0e9a456c39", x"3cc03530f9cb9c15", x"8bb73d9145ef50cc", x"9b5b0e5ee8821e53", x"b229b9fa72a5463d", x"b04ed7424e08f968", x"6506e3322612c99f");
            when 21963101 => data <= (x"1c135ea9e22ddc14", x"98e2a15183f4ed3d", x"62def13a8472604f", x"137a45e7b78d895b", x"e64c1a302e2636dd", x"c42c63abe8ee94b0", x"875780023df87d0f", x"e751e0f16c225a96");
            when 33235820 => data <= (x"7b1eca8324764f13", x"c95fb6d51d2e44ad", x"a3b794b018f5389e", x"1de5a7bec0d3bd98", x"a64cd41ad3f991dd", x"0a13d5c5cbba19d5", x"d71101aa283fca4a", x"2169dfcdf81eecbe");
            when 8320875 => data <= (x"eea466a9f4474214", x"08ca8c29379327da", x"fb6b9ef78d7e568f", x"f392d59a38970d20", x"88660acea10f36ea", x"506a03c240192363", x"06a8c33b1c07e025", x"ab723bb694aca122");
            when 16430090 => data <= (x"c08fe5e72876adf5", x"6724e2bff0615974", x"bacb2c46a6d811a4", x"6930e61c6097f655", x"9fbf3dafd69c36e8", x"3e9a09052defb1dc", x"78b62f48ddf09c7e", x"9121d1acfde0df3b");
            when 25691706 => data <= (x"abfa02aed858b83f", x"cad879f34b32047d", x"37c3e9a55ed82b9b", x"1f244b96cdf71224", x"8bc734a917c6d1b8", x"d7383219064b5d2d", x"1153cb7c9f74e674", x"91988347b23a1f58");
            when 2711319 => data <= (x"2e09990b8f424997", x"ec1097f1c481e90f", x"5f83c9d52375f2a0", x"523e9c4aae8564aa", x"ac742922f0007954", x"76c5fc4d46268269", x"c1af929232cfa385", x"c551198aa883f5c6");
            when 17986024 => data <= (x"51738676b62a4d43", x"6a3c12eab9de75da", x"284d7ba576b42a72", x"0de562e24dd05197", x"8eef58e791c8c1c0", x"e212b1a54d8f0572", x"2351019c97d54ac2", x"dea7e629ebf1f24b");
            when 5822576 => data <= (x"c4338cbe93296abf", x"880f27ee6a5cf49b", x"0588706c8f681270", x"2988c52ecc6d438b", x"3359f0da111265d1", x"f54c0429039be985", x"de44bc75c35f4455", x"bca4779480ef472d");
            when 3791562 => data <= (x"e5ed21161f7d411f", x"880d2c66997ee002", x"c0cfd277eb35623e", x"45cef1cd71bdec14", x"00fb51ae36b3631f", x"756f3d7bef15ab9d", x"3d62479cddae05c9", x"97cbc477c319af07");
            when 14545296 => data <= (x"1495f1b9949778a0", x"69d330bae1204852", x"58eb69d52a1a68d4", x"eabf7d7e3251288f", x"952722dbca35bb72", x"3004848b0b1155fd", x"6013200d40c65ef7", x"124700a05128d444");
            when 13351776 => data <= (x"9c9a0c7dfad09821", x"8aabbece44652d08", x"fe1f5889ffffbcbb", x"0e535542a613a531", x"2d3d195b10ed27db", x"28166c6c5a0c9673", x"0636c0dc4332052b", x"bc8f627026cf6a85");
            when 28587155 => data <= (x"2af97e45706705c3", x"07988e67633cc728", x"ae462500e6217565", x"22810a71d5ec54a1", x"eb59cc6e0f30e61e", x"321228d4a09c7542", x"c7703611717087c0", x"8cbaba7d6844b235");
            when 27919558 => data <= (x"a40ad62076d5a636", x"9aef61f848ba7204", x"090cf051bea0e082", x"a848b4b518660aa4", x"019f41f14af21244", x"4599f74e19416a59", x"edc5107b512e1970", x"89b0abbff3f133aa");
            when 30759759 => data <= (x"30d37cd5c22c85a6", x"bdf97ffdb3f030a7", x"b8679093ed5a4b73", x"57af1af29779f7c0", x"1b89f785dae7425e", x"fd02f562da0f2982", x"5e1e76d6f5a84c6a", x"4dc7fc5f72866698");
            when 17120289 => data <= (x"3d07f19a00c2f045", x"7390a9eb0661b695", x"8cd43a89fab26a5b", x"af318629bc42d0e2", x"0c2fe5a25d495c99", x"5224d0083fe32804", x"61cf22c8a56a7872", x"3935a211b558c537");
            when 11785855 => data <= (x"8caa44feccb9ebb5", x"5e9bedbf6487e07f", x"3b91e8d9c8cc341b", x"b1a6d27e16f39e80", x"56b6bbc73680c5ac", x"2e146f4118b9e81e", x"5c211d464a58d96a", x"e01ce961076c129a");
            when 18550141 => data <= (x"c6ea2f806ddeef13", x"bda1f248d90b35f6", x"d415cc094bc45aa8", x"f9b18fe673ceeebe", x"2e224da12aa79abe", x"14ebc6f015127594", x"9d63bfd389875b04", x"c95e61e93b5e40a9");
            when 31631694 => data <= (x"f80c7d35decbd988", x"afea5799b5eccad3", x"742d3cd7a5020d4f", x"131f84aa3a56d381", x"50b314bacd94ebe4", x"d70831857e00f73a", x"2bc3ab836521c0ae", x"510a00e421af4871");
            when 33471234 => data <= (x"54c0e7fde8866ee5", x"3a7ea5508d780914", x"4c3216ea2454a700", x"e765967a48aa8d05", x"37f4d3ae96482263", x"38c00fdbf3612a0b", x"1aa6df05164890d1", x"346d8c890b24821e");
            when 6889990 => data <= (x"ed4159cc00c6b518", x"af765db967e1955d", x"be78f9d6739301e2", x"fa9b1a788d933083", x"f96bf8ccc85f8507", x"066ec0c246c69b20", x"17ca3cc630d98d4d", x"7c53bb3485a457c9");
            when 22259874 => data <= (x"12709bc927317dd2", x"50aa6df22ea694a3", x"21f62142acb43831", x"a76bc48bb9ce5006", x"93d7792d7052fc1a", x"9abb0e013b9b08f1", x"cce381c5b8ba9c5b", x"b3d2619e64191821");
            when 12852497 => data <= (x"14aba80d09db1ea8", x"6a18c7fb251f2186", x"da0669c405141c14", x"f5bf28b80b59c784", x"0b0a60deaecd3441", x"e708223ee869ceca", x"a597fbc998f9f016", x"9b484ec117d26a3a");
            when 22295428 => data <= (x"bddc7b2bb916bbd6", x"5844f08b1adb105b", x"c3dd161243870b85", x"fc20e234fbff7022", x"e1e0712e275c7a37", x"22fa5993f5607746", x"89245d467e850559", x"6447d4d61b4b7722");
            when 31498870 => data <= (x"5b563ec04f0106ca", x"3806db7af1fb330c", x"723509626cb4d19a", x"2ee0b8eb08b4ab99", x"c80f66bf73ef6e1c", x"60bd2987e9d3d922", x"f5e086479ef20b8b", x"14dadcd56764c1c6");
            when 10403637 => data <= (x"c417e967843d1ee3", x"63c9494151000712", x"e5602763bf3384b8", x"0ce5064e2d35680b", x"ab7288586d5893b4", x"4f219dea65739702", x"d92ed6f754a0e6a3", x"236cb64d75825e90");
            when 6424640 => data <= (x"200841a59bcebcdf", x"a9472f0adcba32bf", x"1a18f46e2f2b1833", x"ce0f29c8ada36d69", x"2774f656b4dc9c91", x"9a0c3b92ab879a69", x"373c56ccdbb538e5", x"ea60ce70cfb53b1a");
            when 7700401 => data <= (x"a0af917d6f1a73a6", x"4cf406d5cb5b5739", x"e2a5e0bb5ca1c0f1", x"93f16a4a2e2f6adb", x"16dfdbbd70fbccb7", x"4214a0efff4588fd", x"e98d062ea2f845ee", x"6b958fc6477053d3");
            when 6714152 => data <= (x"b9869129e14b5ad8", x"fb41a93c4d23081b", x"bbc6c4afba8a84fa", x"f6066b1f16be65a0", x"8ca4038b27763525", x"a0bcdc4ab7f6c254", x"d2c637f8b044de78", x"89bcb3664632ee13");
            when 20568780 => data <= (x"59573ad27ca57aea", x"f5fb59d3961b1c20", x"33e10367deaaf2bf", x"76dc90b687b1e637", x"c5ff59b3076914c4", x"46eddc7c80b4d2e8", x"a10d5d4eb1a59e5d", x"bcacb54be7024d06");
            when 2447958 => data <= (x"919e214a0df9b0dd", x"0fcdf0cf5e458fc7", x"068e6f9b93d4d2f0", x"e412e67cdec3afa1", x"edaeeeb521343e0e", x"dada0eebde9b046f", x"c55b65249968fd40", x"580d0cb435491711");
            when 5083930 => data <= (x"881eeaf18b331d38", x"e30547792f8efd20", x"a107915262e9a056", x"02951995e06a90fa", x"d85927c11ea9a49f", x"d741645a62129fc9", x"8d1763914d450436", x"2e4c065f688a8aaa");
            when 15880508 => data <= (x"232605e4f25786f3", x"51d45911943cc6a9", x"68b435ebf853d678", x"cb5d9a6dcc2a19d3", x"61318ba8032d9aa5", x"50dba7b0440c010b", x"f916e9b64a63d5c3", x"cefecc8acf79300d");
            when 28605511 => data <= (x"421e8d2adf8fc55f", x"4d6860a682b730f6", x"1d4012387cdd15f6", x"fff8aa3256a9a414", x"3968540b407ac7f5", x"e4548964ceef0d19", x"1ebb761726e5a2a3", x"d1ab32ea2c5996a6");
            when 21304416 => data <= (x"411d4a00d6c8f8dd", x"4efc615f99881965", x"38bd402bde971c4d", x"073f67ec1d32265c", x"6c15394a109169b7", x"2496209267d0d4f7", x"c6b360ab4568cd33", x"ce49dbfc2dfa8e29");
            when 32786190 => data <= (x"43f910a3f7698bef", x"42d10d955bdfb721", x"45e28f31af8207b0", x"60a2a9227b0619db", x"f26558d782398d26", x"475745cb0dd84d9f", x"4fe3805b0289980b", x"0b4af47f7dfad3ba");
            when 17980379 => data <= (x"102dbad58521317f", x"48d010842074d1d6", x"5f851add97db4cdf", x"dde83af59d6e4f09", x"1056a19cd4676df1", x"1128cc13fb5c19a7", x"e400b0b783923dc7", x"abc5473431e48807");
            when 13204062 => data <= (x"6dc50c9a42ef3dd9", x"3ca5bee803dd4b21", x"8d49147fc29816c5", x"39b454f8b9f853af", x"ccf5be41ec2fe171", x"c5d4313e0486c1e2", x"9440a6b8c5e03830", x"2c833de9a50926aa");
            when 13959168 => data <= (x"ec84d71c54a05759", x"f89237d0ed27bdfa", x"a22f2876de0dbef8", x"379c8c8dd2353136", x"d75227026a544a5f", x"f66db1ebcee88b3d", x"b75a0b9e4b78fb3f", x"ad2ac936a99124b6");
            when 14396040 => data <= (x"65117dec46f10e67", x"bc664c079717a650", x"86780bd3648667dd", x"1e6aeeb9e6b3e897", x"01e62932e46f4fcb", x"4ff470b72222fcd3", x"9706ac67d5f1c1de", x"da558d94b5f66e2a");
            when 17914674 => data <= (x"6790c7dd281a06e0", x"6a3ef0631eb91d44", x"2c5b896b7c94b763", x"44a308d9f0bd07a9", x"b9cf52814b97425b", x"91ea647c3db103a6", x"a99480ce8739bf3f", x"f71e1fd66685f849");
            when 16402432 => data <= (x"3ac140243870e9e8", x"e458f221c4f478fe", x"36b6d9805d890d43", x"bb1722720f117427", x"91c01f2dfe7b5bcb", x"adc4c7cd619c3462", x"56c35320028de8f0", x"ba4e6a2bdeaaaa01");
            when 12451262 => data <= (x"e3a2ee7e2a7ae55c", x"ae5234d65cf388e7", x"24f6b660e38fd64a", x"42f5af243a737da5", x"f0ed7bb5cbee92f3", x"1f4d06969473c399", x"dab9ad9d88b4dd98", x"62b4e7b80c3554f4");
            when 5121435 => data <= (x"cf2b9140724541a9", x"a062ec33da38e6a7", x"49eb5dd952a022f4", x"df740f185527b92c", x"a6e6b49ea1890a00", x"b0bc4f48b6330d61", x"6a96d6481e171c44", x"116204bb6546de60");
            when 5910704 => data <= (x"d4b68ab29e1535a6", x"bf51ff1cddf9edc2", x"320b575aeddfe5ca", x"b3daba171394f9c0", x"7caa8df4d53e6ea0", x"c4159bac0a15620c", x"57769f77c8eccb0b", x"efe8a9cabd743127");
            when 5023519 => data <= (x"83f8c99d4df0e0de", x"da2af5d794ef00fa", x"7b966e1334ce0a0d", x"bda8343adb0899a2", x"d9879c62eda6a2b9", x"640ab627c115af89", x"6566b6c696d743d6", x"1e46656b2862f4cc");
            when 9423855 => data <= (x"f7cbe46df704dfeb", x"7eedc52c8965dba0", x"8d64cd3eafc15c81", x"08cbd23548239c17", x"dfcbeb0d8894129a", x"e42d3d34e947bde8", x"58f93e717cac47e6", x"9d6f4f3174a29ee8");
            when 24514182 => data <= (x"c346c8331b80a445", x"4ce740fe48c7fc19", x"ad6a57af69783511", x"916e4814fef0edbe", x"5e00a378412d9b0d", x"b0b94494e61e2038", x"718e85b989d569de", x"5cfc45bf246fa8d8");
            when 19978849 => data <= (x"51f33722a697ee19", x"87a0493aaf77bc4f", x"772fcfc58c9d5285", x"1c6932e48b9edc00", x"80c75300ed23381c", x"f7b17200d1658490", x"e426ac9db256d727", x"b8ef9f5f985c60dc");
            when 4048324 => data <= (x"07ebe75f71d0748f", x"10716ab7e15787e2", x"57f35ebadbf25186", x"65c97206208f443f", x"f2e60ecb2457356e", x"d156687aee7216dc", x"e4da9176047db00a", x"a916faec157414c5");
            when 33249430 => data <= (x"dc15f5940a80929c", x"9c01cefe4f17a941", x"bbfcbdede3e71fbb", x"c0b3f293316ed057", x"c06870da2e6c1eb1", x"dc2c4f79408b43fe", x"bc14135a0cf82957", x"c635d242323b95fa");
            when 28352099 => data <= (x"efcbb4d29567e639", x"ebdfffa3690d98b9", x"fc5c93ea05a0a2b1", x"ff07790a01f38e55", x"d6d292396bfbe309", x"498ee007e6e5cca8", x"053163d375cea8d1", x"72fb157d7567c209");
            when 11051063 => data <= (x"9b14d3f117343a5d", x"1982fd9af339f1e6", x"31105de0f90273ca", x"a450b3ed4eccca20", x"c7303615b5a62a3d", x"e8b142e2bdfa1612", x"0e9f96b60c3fa9c5", x"e6a108bce1767370");
            when 21588960 => data <= (x"c9773b884e7d8d42", x"a71f4a1f1373399a", x"c7acd616022e5316", x"79cebad12d6f6610", x"2a6fb9124fae4429", x"5ec5499759020498", x"559a98e978017097", x"bc8a0886d7fffe36");
            when 6775414 => data <= (x"7cae9bd65080ba16", x"d28c1ad3bc79eeb3", x"291c2b57c2c6b103", x"7ee43665c0647cdb", x"9bbd149c0f590f4e", x"412c46822ce86b19", x"54ee63bf2416762d", x"a40c54f750228c5f");
            when 33028947 => data <= (x"6f243936029ab458", x"75a6c2d5c87427a9", x"c9c706363c246f28", x"0bfaa78d963b7ad2", x"1fd241a4707b96dc", x"3cc9edfef2a1c6e3", x"9098dfaa12edb346", x"794ccf37c34fd1db");
            when 29639166 => data <= (x"b7e80d4df7149b32", x"d901d3eefff6c708", x"8cddbec3ed2a0457", x"6682a11484ae2207", x"e4757b5305235c53", x"e6ed263ef1331162", x"51e6d05d596ee0ca", x"845de2ad911f07a8");
            when 16380910 => data <= (x"6fffa2b907fe5cef", x"272b273386e20f4f", x"e264426eabcc6830", x"4ed2677d64307684", x"d5c1225dad016fc2", x"d3177684ba0a0368", x"a0fcba40558a1fa3", x"3dea3a4067dab02b");
            when 22356573 => data <= (x"e5e371afb00758ee", x"cbf84d767bd43aa0", x"56fbab8f54664a22", x"be50a5e0b6a622ea", x"521c6be37f9e29ec", x"8a3af79de0c1ed86", x"21e17eadc3dab510", x"0cfae2f3709e0ac4");
            when 16746194 => data <= (x"0f50ded36d6c4c36", x"7548feb7f68769c2", x"866847f114159b7e", x"d7f3aa7a2bbaf695", x"2dbac4531b8b2a72", x"e2d5130583074719", x"ba736aac0f3c9621", x"67233417fffca471");
            when 7707559 => data <= (x"6188947a99bd40e0", x"9ff4e19b73f1b7d9", x"227e1f426589608e", x"cc10361345da524d", x"8ae984a83496d2a5", x"bf095a35e68bf12c", x"d4234a7016371486", x"313a8c888cd18d01");
            when 23514066 => data <= (x"5dc1819064fac505", x"c7929c763a21aefa", x"d4da9d44d820ef38", x"0317363ad2cdc76c", x"d4935081001925f2", x"ec354852f54bb563", x"c7c95bdce9c18341", x"ee810af49f761dd4");
            when 31082889 => data <= (x"7d4e1613b46b1267", x"6cc80315da0783b5", x"d5b16773b28cda3d", x"aad2d05b1bd7aae2", x"9a730a841efbb562", x"3a6d24a0632b4317", x"01fdca94944a1063", x"689e4a2633d91d26");
            when 13283634 => data <= (x"f09fdf7a52f4b8e2", x"5596504cd708d32d", x"28679155e5395d92", x"60e2d8c4b3a6350b", x"f8c921bf71395cc1", x"77f4ac33cc3bc376", x"3520598922d0c829", x"3a06613cc0081876");
            when 3330256 => data <= (x"5d1a5392b37be257", x"02fc1d4405c897c5", x"b26e7a58df45033a", x"0f91b9a68df70f51", x"35590847b8dab357", x"11104c4f6131f483", x"ed1546b5e89f0226", x"d9145f82fad8da15");
            when 11169695 => data <= (x"4037f3faecbae425", x"5d390dafd727e254", x"f9779105d47f0392", x"332b0367f12c1df7", x"41aaa0ab63ca4f64", x"5b1b6b51922df2ac", x"22049903be1c4243", x"cead9366f4b1b14f");
            when 14964611 => data <= (x"00752a6193067831", x"8daa552123c38012", x"33393833823e967d", x"ca6e96a067e2deec", x"b28112e2c561973d", x"3f2c46999469c08a", x"3ffef70a877c4a78", x"42fde30680004dce");
            when 7197475 => data <= (x"2907e1b3b1861911", x"96f0c49b0da0bcf6", x"96599d5e42a37100", x"b2f0a872a250d022", x"e98dcc6287e846e0", x"36721db75b9fa120", x"c694988cef5c2724", x"1d22ff8cc56fea7a");
            when 1055314 => data <= (x"c5b39987875f6f72", x"4685f94df7e99e34", x"d0d422dbdb02600a", x"3edf0cc032efca24", x"c92c60e25557dca4", x"1a6ac8caef7997a9", x"62e778fedb9a97e3", x"f6bc9d62da6ce310");
            when 21920452 => data <= (x"1e2b587782e4aeb3", x"a9ee18b0ca7b731d", x"f51a1ddfcafc998b", x"ad34d8d948d4f596", x"7c4917483f9a184a", x"026c7e2fc0a7c026", x"07031d1dfaf3854a", x"387fb6ebaec76e00");
            when 14758890 => data <= (x"b2bdb1b4e52fbc22", x"3d9fa311ae982faa", x"8c0ecb27c1de1a3a", x"92fc5e3c092bac73", x"761e3acd6894a532", x"22239e4811f395ba", x"b74e32cf8d940914", x"ee1948b46caae202");
            when 21170431 => data <= (x"cdee4fb1714340df", x"b221d266ecaf2c39", x"c3fd2aeacfda9197", x"c7e3c94f8a7a5bb8", x"6346cb32700cec01", x"883ebd4565a19d09", x"8c786e1abad098a9", x"7fcc5ff21072175f");
            when 16434370 => data <= (x"0eb097d2e4e586f8", x"e9e50450b6c7b116", x"e291dab0573a5fce", x"fad842a4edef9426", x"c8a7021dc692b7d5", x"3cc82bf0ecfff40b", x"87f903fa5dff6f84", x"45f1ab5a0cf5053a");
            when 12963791 => data <= (x"074ffe5c7ec16ce8", x"80f8c5e677172e03", x"6f315d93d313544a", x"f8c3a15acb540458", x"030d4cbdd53f88d8", x"f90eaa3c036bf9ac", x"10bee1ce8e225f20", x"b9580bda6fe42e85");
            when 21247059 => data <= (x"25f5ea264836a1a1", x"da7c3d3b35e13b7c", x"9bef22d4fd46e56f", x"50e1031d42a28e3b", x"63707160655b4505", x"4014e027a5224e64", x"f59856970c296dde", x"b68e5283923808e4");
            when 18686044 => data <= (x"74eb753d263bc208", x"1ee90015da1f64aa", x"c7eef02dfb4bee42", x"e8b7064bb0a99b3b", x"1d2ff566f15c9108", x"ee442d4198f2d545", x"3187eb70a6fd93d4", x"3ebbfb020961cb35");
            when 18331447 => data <= (x"f4488bd7707ba4ed", x"cf70812144f3d0ed", x"5981fe6fc821255f", x"6b0511e8f850b40b", x"856c80685178582a", x"584a7ddd086fe673", x"1e25bb1caa219d80", x"af55054f31b541de");
            when 3969295 => data <= (x"7feea35c2cafc94c", x"f00f7fb697819f4a", x"20476d304cfc5e4f", x"1aef72267b5acf3d", x"227ccbf54babe609", x"e7aec386ddc25989", x"86022e05bbefc03f", x"0dba15cca0de3a57");
            when 17186525 => data <= (x"bd1ef6e979594e7d", x"133312e38063d3a7", x"5a592743ac34b06a", x"846b1f104982d5de", x"ab15add54be19eab", x"518844447116e5df", x"20b7df20ac56e9da", x"53708beed186c095");
            when 29004087 => data <= (x"3e70a05e09e0f225", x"06df5ff9a3956c16", x"fe032710927aa05c", x"216e08fd9c1aa157", x"dbbf9faaa6946459", x"e8d5cc8a4c0c8465", x"c42bd6d402dab4a8", x"4fd57c0400f942e2");
            when 16589251 => data <= (x"ef8baaa9a169c17c", x"5597a2118f5725e8", x"6ed8cada0eebbf62", x"c4ec196625def855", x"88eff4276efe5eb5", x"b9a1e40ea9d87389", x"52235f74945ae5e3", x"d23b4d9ed1b08d89");
            when 28493081 => data <= (x"3cf504a784a62a21", x"f55e04a6ca8636c2", x"22b634cf1a8e713b", x"4cf91b80a9fd6aea", x"1b734c5e71fa711b", x"fbd57e4262e1bfb3", x"9bb17724382fb379", x"889b6ab81f2a3879");
            when 12811556 => data <= (x"8d7644e9aa8198e3", x"77ff960bc9fd8ffa", x"606980bff704fba0", x"f009189c60d5450a", x"f6752c13ebaf8ca2", x"d2cf9376da1c25d5", x"509c42fb102bfdda", x"0bd6c6a19c86aba1");
            when 26019229 => data <= (x"c181d83f3f8383ce", x"15d3bfc0caf2e4c7", x"8c81d89f7d40c067", x"78dbe2134599ad79", x"70a0ecaa6873a06d", x"4045149e2a797e8b", x"054d4c99b275c071", x"425aa3b3c554f89e");
            when 11559467 => data <= (x"01e033aaf11019b8", x"377b22d5cfc20ed8", x"6f7a1eb6926aa1e2", x"7aa86141f8998631", x"163d16b5a9973bb7", x"b21592424dca9ecb", x"a94c20287c67fd68", x"be00bbc8e9d2c5b3");
            when 4992773 => data <= (x"5b79f568d39c491b", x"262d22acd368a743", x"122f6bd2d1dd8bb5", x"5a6d829e89f3144f", x"ab1f5b1157599d20", x"de7f4d1acb24a03c", x"df23b076eb9fa7c0", x"9c0c1b5bbb241bee");
            when 27305968 => data <= (x"8708fdeec78a4c90", x"ddcbe450949934b4", x"32fd963340d9b25b", x"3f22c96b4aaab18a", x"755bc9d1b1105c1d", x"273ab55e66ae5a17", x"aad16d3778cc0f2e", x"204ac868d6c25233");
            when 24923341 => data <= (x"008b939505c425cf", x"aead0ce7f9e090e4", x"4e1543a74fbf87f7", x"5ed405974d9f2d8b", x"9620c94d7a4877fc", x"3ca49a01014240a4", x"47186667d1fc9a5e", x"2c3afb09151b20ff");
            when 32026050 => data <= (x"04d2808593a92f02", x"18e3cbe31b6239d8", x"f7fafbfa7a6bc233", x"628dc650a658f121", x"8aa7cc38f826ddb9", x"5b8720ce753af4a8", x"30f1f647d4fe6448", x"895a719e632fa1a8");
            when 29858801 => data <= (x"75d091c85df5ba5d", x"21171f71e8e7b8e9", x"0b358714d3dd3f6b", x"5fce93f24e47e97c", x"013be3a9f42d64d4", x"26daa48b27f2aa7f", x"97172f6f134e672d", x"273229d45ad2d296");
            when 1891775 => data <= (x"cf0258bc4297a03a", x"24dc4284a990d8d6", x"aa1fd7325c151fea", x"0df90b5e58c35f19", x"9f81ab75142fa46c", x"e871eb901abac215", x"2cdf168657e66dda", x"a5f7ed74be61e61f");
            when 10476629 => data <= (x"1719d25d839e6c13", x"8ab04f577f023bf6", x"d3ff28e5656feae8", x"c976579492761cd5", x"c60b434c4feaaec7", x"47457e059bb6ced0", x"63a2df0d39d70b24", x"fb2ee94c180c9708");
            when 28257880 => data <= (x"8eb5b64f77063593", x"7bfba41c7897502a", x"ec8b12cc1ab94d1a", x"22dfeaccfbeaaff5", x"78f55262d2353c18", x"85dd1f218995f7af", x"1bc2761c2d343a65", x"1ce53056d17ad02a");
            when 26119269 => data <= (x"0be4d276305afa8f", x"89d10aec3d833740", x"a05ae72250cad5cd", x"536b911a54820c38", x"f6e3ac7f4b0b8d9c", x"32f85f1f90c2dfb7", x"6bf7781926d28857", x"7918fb72ec4cead4");
            when 18314808 => data <= (x"dcd04f07d817d127", x"d54b41f4d6fcce89", x"ea26365a10535460", x"7f184092082d9e0f", x"d5bebc72e8748b58", x"7738271167675ab6", x"deb6a49ae171963f", x"63876fac24c0fa48");
            when 21603311 => data <= (x"5f678aeaebfa5541", x"72c9dd576d129375", x"1118e8e3b95cd252", x"d0eb877c6b575c1f", x"b2972489cbbbb4dc", x"0d97cdd99cfa70d7", x"c1f524da938e76a4", x"ad1f70fb73242dd3");
            when 32300994 => data <= (x"fc62e67c0cd064ea", x"7c42dc75462a19a8", x"b9a7e48bd9c25286", x"abdab8d981b9cac0", x"95a706d0162ee4d5", x"84104529eec3d3f4", x"56dd46e5da8e0c8a", x"9009b58fc0dfcb6a");
            when 21658091 => data <= (x"0ca08e1e650293f0", x"466a41c7e537fd70", x"c25718712ef55fcb", x"e5fb2b7186bf24f4", x"888bc7bee27e211c", x"4744fcf3a0a51546", x"aabc5d7856f882c1", x"f9b7bc99af9f633a");
            when 17397557 => data <= (x"f2b2972144fe84da", x"9870bde0b30f9a02", x"31bcdaa457c7907d", x"ed1da56d69c5fac6", x"05b706ec11e3437a", x"dbdf88187fe6d44e", x"001b9b8a7e9849ac", x"99ad602a1ee3fc4a");
            when 26869830 => data <= (x"1da46725fb96a9b8", x"9f6472220590d8f6", x"56b087fab1d466ae", x"b4681a5a9768f1d6", x"77253c717016f63d", x"b0d9199d071c6d6e", x"99c6befbe32f62ad", x"6af404eff921a6ab");
            when 5227544 => data <= (x"c45417b8a21de52f", x"fc9836b6c6e2475f", x"9e639c101532fb7c", x"9e13196cf865cc2b", x"911e7c93b0c18cc5", x"2241d26bd2e0c01c", x"be3a09cdc369a96a", x"36b63374569c211f");
            when 22027196 => data <= (x"4540de9c3360dff6", x"fa4d0d18afff9ca5", x"a6be1ae378f3b256", x"e13f0c91584c96a4", x"40654055d0865ca0", x"e51843ccab91ce04", x"e4137cc4583445cb", x"128488a16d926579");
            when 14123285 => data <= (x"e64d2ffbae93f9ae", x"f11502a6ae518566", x"1abea6a29d75982e", x"a9efc96ffa527b26", x"072eb8d8ddac6f92", x"e5ecaf2ca3abb3cb", x"fcd90ed7e1b11b86", x"a8a3251accee0aae");
            when 10257467 => data <= (x"7204dcf23aaac7de", x"aabe17478f367702", x"d801ebca538e3cab", x"74490605bd9885f1", x"9c3974d6fc160c5b", x"6c3d8341a4565549", x"d8b3e9ea0d5b0b68", x"6c15f8ed93dd3ba5");
            when 3246327 => data <= (x"03cc87d822ecb3f5", x"300d8394759305c7", x"59901e8fde763f41", x"040d61cac22a41cb", x"2fb4b5544aac41a1", x"4aa6df6d7ca24e19", x"728d861963e52df6", x"d5bababa9ffb14c5");
            when 32386429 => data <= (x"fa6b6c7fc812f51e", x"2967277273fc5be0", x"0aeacaf8ebcb8d28", x"a9dc40a51fd7b1b9", x"d31b1bd6404c6463", x"084c90df9e84418b", x"fb426c23cd62561d", x"b3de9265baceb68d");
            when 6491130 => data <= (x"754a50b6fcb164e4", x"31b2795143b71a52", x"00e868c1a8ecab15", x"062cf7aff590b638", x"be3eed79ff5526a1", x"7ff256537f27dc20", x"e8d7bd9769646036", x"7ac746eb41bac40e");
            when 18799336 => data <= (x"7dff354a7207f758", x"ae3fbddbf07e1fa3", x"abf045b5ae84826c", x"df1232286a6358ca", x"f619f0c1c74963b0", x"e114311fd0a27add", x"4a219e2edb7772a3", x"93df1ba821b44037");
            when 3408096 => data <= (x"09687a0cc55dfd7b", x"26e961972e0029be", x"d0bf216e9454a6b7", x"bdb522e3c20f24e1", x"6a5df3720e3b721c", x"4126c2b4344e7b03", x"dc2b8335f2af0f73", x"425b71950cacd2b7");
            when 31239908 => data <= (x"a98883b47f96c0e4", x"ad16bde8bd3f4b4a", x"9d0042fce0a04048", x"2a4e88c9e83f2bea", x"940621c93f4a6ebd", x"16176284688b13b6", x"56b862ba50c73e7c", x"f9efd241ca8fd38e");
            when 3963915 => data <= (x"fefb800bc1d2bb90", x"f11df0f7e84c4e00", x"598e0df684adf344", x"c5508a28a596939a", x"91540ff0e543d7f9", x"99e300aaf23d407a", x"21796b74d626ee50", x"44e0fce4c7246772");
            when 23072891 => data <= (x"764872f38ca9627f", x"bdbcdec1e5d18523", x"29af1aaa103858b6", x"6fd4b71a5566469f", x"64c36e7786cbdb73", x"5eb9805e7df73e31", x"fe2a839c445ca72a", x"c35b85983cfac875");
            when 14196777 => data <= (x"ce7d7195b86803f1", x"66cff73ba615f2b6", x"323cee38a006fa91", x"8683a97bfa0c5e21", x"40ea4c45524aee77", x"938921955e26c9fa", x"f2568b9b074331e9", x"70a8da315edabfad");
            when 32453781 => data <= (x"819685e3e690ec2b", x"3ff55a43b68647ee", x"7a7eba85509dc8c4", x"32d8e244cc1e3e1e", x"9e428a429cbfc2f0", x"27cf63714ec5e382", x"8f3ff8f343d224b1", x"ff1fa7d1aae59457");
            when 2673499 => data <= (x"da7ccbbf9efb8421", x"a326e4347740feb7", x"e8861631c3622836", x"77932400453b1be5", x"b95fcea91c1bddd6", x"ab2a3a0a359abcc0", x"edd9203612da1a11", x"216b8749bb42882b");
            when 14265232 => data <= (x"26ab543ff1e96b4b", x"31d7ad16ec404fed", x"50004c1ddc2c684a", x"3e1314f4ff8b8f87", x"36bbe8d4d49f7318", x"ce9f8365e206c71e", x"0221af61a5145002", x"2d04b276d485fc59");
            when 17636510 => data <= (x"e097f038072ded23", x"2e09b7099c48e1c7", x"def6e17d91833544", x"f4ebf692cdc9f024", x"5483c22f731d9621", x"2f7235acb4d8c3bf", x"13d95edb3cce1bca", x"8ffc07008cfc50c2");
            when 9305982 => data <= (x"cae5eccc37f8fa7d", x"f1c8392be21c5c23", x"320461a1e311db18", x"4cc9f62cb7f15411", x"f973f2e8a7d46d04", x"fc7313ffa8088119", x"021c5637da68c104", x"b19726b5d542fcae");
            when 22631175 => data <= (x"feb82c4bf6a13b07", x"f3ccd3166bbf478d", x"85dce5839c863899", x"f353648ac52a3ae2", x"7a75d634b3be1f88", x"3f69029372a8441a", x"4c8a47169759dcb8", x"b6f1fae16494684b");
            when 27986748 => data <= (x"39d56f4e2d42d27e", x"d79fbea0c5317c36", x"2e8b4e2ab4744b37", x"b8661c9adeb3afed", x"22e508a2d8065cbd", x"c2a4990469fe2775", x"63359e47a98ea20f", x"199c2b6e4eae859b");
            when 1412952 => data <= (x"b5e99de5fd6ea87e", x"4f4230fc401cbe0c", x"e47ea99326fe1178", x"a275eb4ace9a5f7b", x"dc79c2dd4da1025f", x"d11c3b56359498a6", x"338eacc50469a6eb", x"e73e71b79ed1f2dc");
            when 20419835 => data <= (x"efe2774cc5544ff9", x"264adea1db2753b0", x"832b1f96d874757f", x"c2fc9d9ce48c7d11", x"0cb8a63334c48d92", x"74990a8a69e94a04", x"b685f2cda22b9e50", x"fd9d23ecb8d89290");
            when 3940058 => data <= (x"c6da8f0292e35ef1", x"d114bce58e075915", x"77940186dc63f799", x"45891c61a724fa70", x"c7b6d59e8d2ed1bb", x"c65eebd6a0181913", x"003051ca261c472e", x"6ad15d0b9b3f9b59");
            when 25577142 => data <= (x"74f95bc4b3cee9a0", x"1bd86afa1eaad274", x"f38560ce4fa297d9", x"cb5b36adfa29d596", x"228dd17ee6f7ee82", x"c25f8ad8e13e27ef", x"f3448d97d956b1db", x"5c312a0ce27d4292");
            when 23873080 => data <= (x"5a39bf2bdf0a1170", x"57ef898a9fe3797f", x"b1e49ebdc2175003", x"6a98aea9172e5be5", x"4a53d18d9babe184", x"65090e0845bb57c3", x"ad88dd318c53ca2d", x"e96a0c84746f894b");
            when 29151473 => data <= (x"794c3d0f37c7faa3", x"28658faf36cf3f1e", x"0b4cd18cace80120", x"1cee5600042235d4", x"133fc8e4b209c655", x"5b6d24fd0f2c5d50", x"3364e0874ec6b182", x"b4ebeb3bd7628f0e");
            when 30030154 => data <= (x"0714e40363ac236b", x"9537fe8f4a72d8d2", x"35d70cd3108147c6", x"8f26398444b43a9d", x"62d20e9c74d05253", x"e248b731ce1444dc", x"291ef42450a04550", x"e8d4c61d4d078af1");
            when 13621768 => data <= (x"31eaf05c800b4ddb", x"67609c992d7217ac", x"a3e867cfd8d44004", x"6a01a101b8b83dbb", x"29ab7654594b5083", x"a9ff913d3a0e9674", x"2d0177cbbd54e52f", x"ad83f0691a3ac980");
            when 1914164 => data <= (x"64b984e53d9ab30a", x"1be7f38cd2e2127e", x"7a8684543f260cf8", x"faa0758fbf3f5a8f", x"985dfe712fea15e4", x"e70db4dffab607aa", x"2463d69e9e0ed3c7", x"c89a0c5b19758790");
            when 20828540 => data <= (x"8b538f06fc3433d1", x"9baf8b6f9a92ebd5", x"85245852cdbde722", x"de4534c3f7b33ca7", x"d9c998ba47779e89", x"10f50fe4f1ae7459", x"63e0250f673899dd", x"039b4206430dd2b6");
            when 14547597 => data <= (x"b605b4f6e638a676", x"fb5cb21ab6537828", x"f0624f2603ebce46", x"d1588045404930b0", x"aacbe7ddddf74221", x"4eb909c7bc65d48a", x"20c7e10a58079430", x"b80c627fe939a2bb");
            when 7762326 => data <= (x"a38184af972e9620", x"0e776df2199aad57", x"03709ef530a5139b", x"7618241b82cde358", x"68e0dc53c8683b64", x"6e5fa2eab5ea4075", x"6dbbc1b50a814481", x"66e569c3e34c73c1");
            when 28786358 => data <= (x"bb75fd9a75e683ef", x"88a531c038aa5081", x"3829cdf206ae3ea1", x"5273e63a62ddef24", x"e56cadd10fd99a59", x"f42137f5993880b7", x"f81655a3517cb353", x"07aae1da42b7afab");
            when 14307528 => data <= (x"f1ff48e7f8409186", x"70babdb55513d566", x"692c94e91ce674e2", x"1675a108693f1795", x"dd265fa2c10cf2b7", x"c8e5ebb51657fa9e", x"7dbe4cb46d0f4504", x"be76eb1fc135fa78");
            when 10212541 => data <= (x"13233d3756582ea8", x"f610333c9fd6bc0e", x"0aa59db0b09958cb", x"46dedbcc95e0eb7e", x"0383fa438cf401f0", x"e6c1e6f3512aab90", x"9ac6a61bb1ac7daa", x"852efa0cec6a012c");
            when 26278943 => data <= (x"b994b2d710a83e09", x"5b97dc0fbde3fb45", x"245c78e862328d1b", x"43d8cb5d388c58a6", x"b38ee3cca12ee2fd", x"41b0bbdd36613f72", x"448a2a330f495c93", x"e37f07427ca75ab2");
            when 21448169 => data <= (x"3127aebc2c8a5105", x"2797de63a9fab6ac", x"62f73773eea9f261", x"f498007f5bdb1107", x"a6d57767748846ca", x"64f99ff3f52150a5", x"2e025fb934ddf287", x"10860408c35619e4");
            when 16075206 => data <= (x"ecea126562a4be0b", x"86bfccd612fe843c", x"f1443b89a3ad77f1", x"c7f60a6a9146c2fc", x"792d5438dd3ece7b", x"53bf477ee33961e1", x"1ea5b65c2a973ab2", x"fcf543844f283b61");
            when 25211090 => data <= (x"968f643a3268aa66", x"8817e3923bd49697", x"bddeca412ad81fea", x"358a0ed68107b690", x"c6d8a74f4ccaf263", x"b07064d59ea8d0c2", x"c50379a8f7e075da", x"932dab483e9c5068");
            when 17262800 => data <= (x"2d162697239d6e57", x"25bdccec73135594", x"950f642e21903431", x"6aacbfc2105a5c2f", x"727d5524ab4b4b12", x"13f7a21fc723373b", x"3411e84ebb0a7ca5", x"58ac9e2abd6b271c");
            when 2060759 => data <= (x"71c66c9d2356f17d", x"339f17f68db61ad4", x"84c7b30aebee13b3", x"440e68b97227a136", x"6ac8ba8891fea888", x"7111224e0586d5c1", x"52ef904071bb96b1", x"dfb878821170bf75");
            when 24933902 => data <= (x"60e8d5d83c42da7e", x"791c2a15ab23761e", x"407acf0cec657e92", x"44236707acf94fe7", x"a0d8cc187c08f623", x"2cd2051beb8d4acf", x"a58c7f91e8e117fe", x"b1dc4e07b7a787d6");
            when 5688340 => data <= (x"1d8f211dce4e1658", x"055dbd7f4b7d2ded", x"c18923a19080b60d", x"32ff5006ba12df53", x"1c3654867f5007cc", x"bfbcf2817b454c5f", x"e61812e5d8e6aab8", x"5bb36f555fb21947");
            when 22331729 => data <= (x"70146eee144ac05f", x"df474a4d1e1babcd", x"f030fb0a602bbad9", x"097fc42dc951a876", x"954b663c25243e97", x"038faa55026beea9", x"7e6cb60c02a1d337", x"fb54b86a79154cc1");
            when 26149663 => data <= (x"6738793a66caf327", x"175af6df5a6d1301", x"5cfc87f6da742033", x"821fe4872a88f4f5", x"9931eefb10e289c0", x"bd6b914655b24b74", x"c288b626f7183c07", x"3fa61c5bbbec4751");
            when 30537248 => data <= (x"4b2a987496e3f700", x"0d42cc5a6d7d7c76", x"2bc219a144f64766", x"4223e16c90366929", x"8ada1b6c1e116477", x"12621bdb0693bf88", x"ca497745905454eb", x"821c1cab530e6b8c");
            when 20108444 => data <= (x"95addb179015c118", x"c111ac697f8a01e2", x"42337776fd250437", x"23cc6628b04ced72", x"43898272b4a937f8", x"36c10e45314c7e8c", x"f15b20ae2d649bca", x"5610a2983d55ffe4");
            when 23101180 => data <= (x"6ce37d90cfe1eb27", x"c19b9c5266ad9e10", x"8135210444cd389e", x"815b0a47c47b837d", x"43bb9b883be536f9", x"d282337bfd492f2a", x"09c04d4fc8c4aee5", x"7daed15eeb8e28dd");
            when 16056336 => data <= (x"db4c473afc073331", x"702d2395f0b4d34d", x"61111721a17c6f5d", x"d038a5fe76b8abc8", x"0d3feadaf5f93b6d", x"3a46f9fc295a9c2e", x"5d26ca4b187ebf5e", x"60b560ae69aa96dc");
            when 26323632 => data <= (x"4f8e496cb65498cf", x"77644505d4cdb9b0", x"e0054805408bf55b", x"3b4b41c54ab0bab5", x"e9591b3311f2f06a", x"f3543437fe48e2b2", x"f53ce9c275117bfb", x"0284e49ebde35bff");
            when 23245084 => data <= (x"d3e1d136a4fac191", x"0d589280261772a5", x"f5b90e3fa84c1f6c", x"77e00b3947ef0f90", x"726c453b437fbf6c", x"ea2ce00c1a7b853a", x"5e001cd35815a6be", x"7d726859dcdd1527");
            when 2548048 => data <= (x"f58ead4347fecb8a", x"969ae44f7b5adea4", x"a425913cbc4f513b", x"e490234915a7f25c", x"aefd44c226be2d2f", x"f29a609dafcd5d2b", x"326196f338ceb62e", x"de0114e0d181c66e");
            when 22561539 => data <= (x"674a63940341c035", x"333f6a95eaa1e439", x"7c762c9a947a185c", x"abef73e2070259da", x"ceae52648345fa76", x"f768fb2c0df0287f", x"cd3d1199f2a874de", x"845b1768ec881cee");
            when 5559756 => data <= (x"4c67402a5cb774b9", x"22bd6f6f54374e4b", x"7b1387fa84200c29", x"6a4113e7cb825235", x"8ffc7ac8c81d728a", x"f27e515ec610a261", x"e4ec6f15334b3d10", x"708b5f155bdc01e4");
            when 9823834 => data <= (x"6dd7c4c70f3be030", x"ebd06d2c47a577e7", x"d5ce364c57178629", x"334a432a75abe917", x"88e6381f6b155985", x"9e021e6dc7ecc654", x"52915728ab21d990", x"70ff334889afc460");
            when 27013826 => data <= (x"846c02c6aeb5a5ec", x"c141c20a1a59d05e", x"d3e496bed9f07d1a", x"9d1e600c0295272a", x"f2dd90165a601d30", x"918df410251fe2ae", x"8ec71a0128670997", x"6819a58b28bb1204");
            when 1587084 => data <= (x"4f282b4c67efb51f", x"120e875ece7c52ef", x"e0b619220b996b32", x"7f91b6e3ac333846", x"51504b8dda1a5d69", x"d10369794cef4b6a", x"2e854115211531eb", x"e971e999c1bfc526");
            when 15171357 => data <= (x"b91e342218979cf7", x"e5609cd0f8e6e0ec", x"d48553c34de80c92", x"a6b4c98900b64a66", x"6462f64d30a0a72e", x"6db6ea8b7f72ba3e", x"58ae6cba75fc8d36", x"7d3baac47c898a80");
            when 32753780 => data <= (x"49fe2c27ae5ccf8a", x"b586699e5769e2c4", x"2f25c779fe2f94c8", x"5bc389701c34bfca", x"716ef68c97eca119", x"bff890079c9670bc", x"a742effc8d27728a", x"1f98476e7beaab9f");
            when 27315148 => data <= (x"5bee79d21304cdda", x"da9a7be43b588837", x"fe47e72d397b141f", x"08fd4ce322a5d9cb", x"0cf42d2d834eacb7", x"3d2046c5bde7091d", x"96b2af135d8c16ab", x"948188e466359794");
            when 15561927 => data <= (x"a7392001fc26dcc0", x"309e699e4c1dcc02", x"ccc600f3ab3b0773", x"33da635a38e6e481", x"444ee731314bddab", x"04a0ead89e1ca4fb", x"fe220a3194295285", x"6eabd6ab0ffb679a");
            when 3614611 => data <= (x"732d0c91f9ef582a", x"b2f08dd46594d0fd", x"f48e80215fdd091b", x"e04f1b23cc6545e8", x"50a614abba9e7432", x"b05ea5019c99d572", x"ff4b69584a4c7d4f", x"12346dcc6a7418a0");
            when 7788566 => data <= (x"2332747dceabf797", x"a66b9f3ef554077a", x"8bd7405d5085aba8", x"adaf39d1bcc8c4a5", x"c9afef6b99eb0378", x"ec6af7ba818e2272", x"fc37c400beba19e9", x"800248022a846e46");
            when 15939366 => data <= (x"d82f494171f8761d", x"6ec36121936d4658", x"6cbe40c6b131f06e", x"636b438de2b1ae14", x"ee0e756c2beb0c67", x"1908111f1be3b8e5", x"65a9f06ae8d84689", x"7513a4f639b2cf8d");
            when 20559801 => data <= (x"920a72a34ea6c729", x"7bea4faa08207238", x"5b0dfc00f219e73b", x"e73ec3b1c1c1b218", x"4094e168acb8bb2f", x"a805f45d90ed1b0d", x"d3b1b9645ca287d7", x"f9adf1af2631ab3d");
            when 30606975 => data <= (x"1579c91ea50eb393", x"6056be123be0e280", x"f7cb28765ce742c3", x"dffe3a44af37b4a7", x"8d8c8768604995af", x"6a728a1f43d01a97", x"ff9f99f2df56f973", x"dff7722583d63caa");
            when 3750300 => data <= (x"b94852ad9c7ea302", x"023405297b6b7940", x"9b2e7d57701b5b77", x"27b32607cfe98fc7", x"ae8bc2f02dddad7b", x"e7e7e01669667593", x"dd3a42953d1ae50b", x"0b98343b382e99d4");
            when 26507647 => data <= (x"8c45d34fd170be75", x"a6a4248bb988aad3", x"b897033d96dec19d", x"ebf857d8a2adb953", x"cae146943e4c1f3b", x"fbed14b08a03f007", x"5cbc16def08f187c", x"3d747f4ab4edddda");
            when 21923172 => data <= (x"4f25cc1588f3f9be", x"a41e5fca3d1212a1", x"ed8188d716ddae59", x"0e0a63e561c96688", x"b4f7b9bf039cf211", x"89b27d779e4adebc", x"058e9823a5b56c0c", x"31e91b7d63f6ca9b");
            when 7487806 => data <= (x"bff7aa76921d143c", x"6e63318c755dff96", x"8fb186373b8285e7", x"2367270500a1dd8f", x"40adca31b86ecf87", x"de732f8f32b47b88", x"8d1fda76a6f7f897", x"bd5a22beb528fb7c");
            when 28323967 => data <= (x"b175fd1a5cce7b59", x"231112b481d77a5f", x"7b68a31f6790f09c", x"d59b1ad7e027cb78", x"ff103391642f4d6f", x"99cb78b4cd4ea23c", x"90d290853866aa97", x"5a7608b12b403ac0");
            when 3735692 => data <= (x"ade81e295c811b1d", x"233b3bcba3d34452", x"99c4a20d1cdcc708", x"e745754f56c5a2c5", x"b120c15ad96c4ae9", x"448f39cfc7df4d33", x"e871da6d85dd7ef8", x"4b292b53a1ffc835");
            when 10866696 => data <= (x"03492d852f2d7513", x"3ee5e84aa1771bad", x"e5ff4ee59da8b3a7", x"f25efc33578fbc18", x"f80b8f9bc8bf0562", x"1f9f10f98597f79b", x"c5d63f81b5402505", x"0d71c7da18b08bf9");
            when 5400964 => data <= (x"67beba5011ad457f", x"7a037077f2f167d3", x"8fca6219cf0a99ca", x"07749479a1aa8004", x"d79b01a82b8b1325", x"9d7fdbd510740694", x"6d6c23462562cd11", x"756c22aeb3b4538c");
            when 4413849 => data <= (x"2fc273621b5b2312", x"9b9fabab9356998a", x"1072d720f103fab4", x"f6395d48a6708130", x"84a5a8b613c7ac67", x"2940f158aacb500e", x"6b2ff1f91283b6ef", x"74fe89a2cf18ff74");
            when 22904948 => data <= (x"9041a93c211489c4", x"cd99be5ae04baca8", x"fd6e2311ad86d2fa", x"e1abfabbe4f47847", x"5d0bbb311bdff4a4", x"0c3fcd502875fd8f", x"fbd963045dcb5961", x"709ea6a0bc6a5950");
            when 31733856 => data <= (x"0c7caffb18cea856", x"8a50d60c0abc3419", x"baf317adc4eca2f5", x"7bd614e5fb163277", x"716a298b6277c131", x"864b749e87e843d9", x"966639fedbf1a873", x"302afbbbe53166e2");
            when 27261674 => data <= (x"6b89772b623f263f", x"db8a09e66ee28a92", x"787a18d929514ab2", x"b36e1b72abc6af16", x"575967f99b873d00", x"0b0c658f1c7ea464", x"7350b454cd131890", x"a2d9a15523654315");
            when 7393966 => data <= (x"1fccd214bd121996", x"4c33eaeaba5a3402", x"315438d83a6ea371", x"1d01b64e2f350f68", x"1439d129302e91a5", x"c240ba84899e1513", x"37bbeac0c0258ad2", x"3b166d43d46785ba");
            when 24120562 => data <= (x"1b0347dcfbc7ce0f", x"7ef95c7ad4daa3a8", x"3ac614e1bdaeef44", x"e9b719c151a074f6", x"3aa2557df7b4999d", x"c0f832af1925dc83", x"67a45a00945afccd", x"d202996ffecadb80");
            when 16724303 => data <= (x"890f5d2ac21cbc04", x"84f678b78eed8726", x"3d4c8900f2dde973", x"3245f8a0d424559d", x"1a3dc76082c1600e", x"c752ba2f0680353d", x"104fe48456d51387", x"9c8ca45605ddced6");
            when 21170086 => data <= (x"b9ba63c693bfeac8", x"b1b5ec45be49ad79", x"85668b2fd4fd01d4", x"7784c137c53f95de", x"ebb5b233232f0d6d", x"a80bb991968e1513", x"a13b7c805cbabafa", x"85b27632d8c45c86");
            when 1810485 => data <= (x"9c495579d98bf7c4", x"ad8ee5fa15fd6336", x"cc6d4fb803863570", x"d11926893490056e", x"cd13c5348e7a39a2", x"9e90291166c21414", x"ff78dc8329fc31a6", x"0c607140ecbee1d8");
            when 6034559 => data <= (x"0cf80b726592364b", x"8cd8af974b2701d7", x"d7d6cc545ff64133", x"b7b84b5c095a78b5", x"bdeb2aa5e692a43e", x"351d276443c12153", x"835d96ddc27204c9", x"cb379867a9354c24");
            when 28317569 => data <= (x"98cd42e205c761a1", x"1a51974679352cf6", x"d3eff557277008a3", x"af641590e80ed8d7", x"8b9606147ea5dbe4", x"097e391a7d1c130b", x"ee0cbb67199d8459", x"a0fc894a2e978411");
            when 362407 => data <= (x"9ba306a4d7e76e13", x"59162307ee6d2341", x"521ee25e4ffca78f", x"2cce1b8404e6fca6", x"a10c3195e9bb84fa", x"3f9c44b19b8ba9a2", x"0191dcdb575c5642", x"4aeebef108903fd5");
            when 21429521 => data <= (x"dfd9e58d86c5bab0", x"20c28d296b62357a", x"317af37aabe5e13b", x"365686c66d110598", x"63a651f6aa5a14e4", x"36727ce0ed236f5d", x"84ec3d1436a931b8", x"5bdfcb3cd0bf2c80");
            when 25273823 => data <= (x"c97133f7d1800597", x"de830fda9fe6c597", x"7768f7812dd33ab1", x"c638afc56fa39872", x"3ce02d9df7b52ea5", x"cab5d98d69a56efa", x"4a4db4d7e2ff5921", x"695309f4da9fdf0b");
            when 33294130 => data <= (x"5649db711cc9feab", x"ae00356b50f877be", x"5facaf947b71178f", x"ca5c38f0d1e5276f", x"e82023b92796d434", x"3dea18c430cfac3e", x"9941b0e9e2a98d9b", x"321e0ee9d8e625f6");
            when 24372796 => data <= (x"9cfae330f7b15843", x"7f0cb9f33dda1261", x"b700ec3f65871274", x"59de5a841ab08faa", x"08f6e5386ff81548", x"6cb7f29fe81d5eed", x"29c0893c3377a9f8", x"92d62821707f0653");
            when 33822342 => data <= (x"cc79db21a002f533", x"e4cb6a88c5b6fc27", x"802bc4a46ed6ce8a", x"4d2ce1fd1009e0c4", x"9f25f062bb5d45f5", x"022787a9a376561f", x"b6173f0df2349d44", x"9246bd39d0c64dc5");
            when 26410135 => data <= (x"e4006017d3b2827b", x"31553156996e7836", x"0741acb4ce3ee36b", x"908ee361f80af5ec", x"d9d687ee9eb8f68e", x"f28a1b9f122eba04", x"a82aa071b2428b99", x"32cb8fda96195233");
            when 6960710 => data <= (x"d2169435b8da7b0f", x"9417b9044635f050", x"bea703e2cc392898", x"1318bc3b2dcb5455", x"2d55c8cdcb3c055d", x"76dc798b76da60e0", x"bacbfc6a8de9c9c9", x"0bb1dccd964068e1");
            when 29682983 => data <= (x"66b5e3c7a0207f1f", x"0a0dae2ef7cbff46", x"463b466e1391450a", x"f985b5fd66cc4821", x"2350d4d5fd6c61a7", x"7c3565a0592c3d01", x"4d65a90891019848", x"f2f5459c55b99043");
            when 19541103 => data <= (x"0bfb88d2a2a92466", x"c6134b48fa298a31", x"820c6d1a0775611c", x"60e25ec49f3eb419", x"54fb16e53113a37e", x"76764eb05936160c", x"87d07e71e6cbe5d2", x"526c2f907435cca5");
            when 13347120 => data <= (x"a73bd7b4ab38fdc9", x"aacf4e17d201da95", x"535a3e8367331e0d", x"ece7b4f3478e015f", x"418caf9525872dbb", x"4164544a2bc2a2eb", x"5eb55e0e71a2dc3e", x"a0e345d1c125965e");
            when 12364560 => data <= (x"68978f79a034e953", x"38b82df8647d2997", x"b46c25fc89a5e8b0", x"5fd6d7a0a7d5783f", x"aca1aabc29242a67", x"042a3faed1906406", x"eb0f45800b6d3067", x"1b613e4a324081d8");
            when 12564465 => data <= (x"ede1aa5a463c2a7a", x"494305e067dfcb2b", x"f801ccc57c7e623c", x"0643c48492de8ed3", x"a33a967f80816047", x"96e82d9d16c41290", x"111f0b75aa09eec7", x"1bb98833b86581b3");
            when 32291025 => data <= (x"cb7859368a350ea1", x"80262c6cdeacabaa", x"2421cb78e9d84b28", x"815687023401cefb", x"0425f6d04b5945b4", x"3a926dc3d9270909", x"c6dadd01c2b9ad29", x"fd467b6403422553");
            when 29646167 => data <= (x"e0996bd873640175", x"9285b5304d0565af", x"9f5775f8a672bb83", x"a4b7ffba0955e907", x"999dd1b0f2285b67", x"08e372785fd03941", x"19e8825ed9f21e92", x"48e01a372c20ff89");
            when 25456289 => data <= (x"98f73d505003fe21", x"1fa1a6cfd02b6d5c", x"022e8a87a282f482", x"d4139aac8145041f", x"63610da9e9dc565f", x"f5bc206212de7d51", x"f329ae5342744a2d", x"12d0d0800a9e6fb6");
            when 21317072 => data <= (x"42db20f8713ed398", x"78cee96b9fa884c8", x"ac33211a7ef9e7f2", x"7d5b18a8606a00d7", x"7294b0d8dc18e21d", x"a34da573054bd9c1", x"a9007f30205f36c7", x"fa51f476ae5d4a8e");
            when 11361450 => data <= (x"c29138f23d06026e", x"1373f0bd3e3bf392", x"d7920af7d784f379", x"84560dcfc314ae4e", x"6ecdef977d690d81", x"16b4d4487921005f", x"6e6ef4c295c53fba", x"8e76134ff19a6765");
            when 955371 => data <= (x"d5563a87d8631a19", x"c415a3776700ae1e", x"d4fc83b43a2b87fb", x"d83bc63cef996d61", x"d0e5c3d298fd9480", x"19a691e1dc9546b1", x"6659481e49d1859c", x"10c0c044a0cac2c2");
            when 4018863 => data <= (x"369fb3f58a30e27d", x"614173344daed64c", x"fbe0d5b5f8afec01", x"7d546c646ce5fa2a", x"4212f8ebd390c47e", x"913562402cb69895", x"f6dd434b7f106834", x"0cb9db541a3a715d");
            when 4096270 => data <= (x"fd729eadfde95f0c", x"39b824c4dc4b6ba6", x"10c8d9f1751bbf95", x"82e066f45ac35803", x"161226a5abf41d28", x"75d7775973669fc4", x"093956acfaba94ea", x"7b2157aa3dd57ec9");
            when 3565517 => data <= (x"0de201b44406b6f1", x"c30f25d186ab575c", x"bb0282cf7ee45965", x"e0b227c2abc80e5c", x"5d9f13f20a2efa12", x"e9707d657b6e5c0d", x"fc0f8658d4d15c63", x"3082b34c7e5c1272");
            when 15904666 => data <= (x"07ac6f60591ca525", x"f353625944b5c6ce", x"d37f57908ffb9da0", x"7683b460cc52991b", x"a6216131c001fbae", x"a14cc5c6f09b25a8", x"718eb275608a635b", x"04cc903988537861");
            when 19629400 => data <= (x"430dd12429f72eef", x"c329d9c70c94c538", x"2443585155b3b09a", x"ba20d8df2fffebdc", x"db81a28827c68c35", x"62256b341f2dfb99", x"8ee49fd59dd16ea3", x"9f211c2828f567ad");
            when 19450012 => data <= (x"c033c4f8f39942fa", x"92d86f1993c8e513", x"be41aa7c69f7a9e9", x"524a4f5c5ed2597c", x"32f4afb205f33c53", x"0a3e0ed03b204622", x"80a322ee231d083e", x"754fa673b4c47aff");
            when 18317565 => data <= (x"de691cfba503e09c", x"590019b02e50ed3d", x"30b10a99af4194ed", x"23d13e4581888220", x"247c6cbf014d8047", x"b726aaa003c6f89e", x"3c6ffc8e0a91c974", x"a3d4baa3f1a971bc");
            when 17560873 => data <= (x"5c01146e12055272", x"ec70664858dbe748", x"9bc788a96f36d80a", x"9030ea6694d413b5", x"18bb16f45b2baf81", x"25890f9a5688ebbb", x"cf529fe981c3f135", x"b59c64a6f1ed6949");
            when 6544503 => data <= (x"a4aff42988aacd56", x"b54b37434f949904", x"e836741ba2110b21", x"1ed5f4dac14d9d9a", x"39d72af9793f3444", x"a0729a2b104b8abe", x"392eb2ba8f81f83c", x"6c2cf2fc6db2e293");
            when 21952110 => data <= (x"91471238ee10ffc2", x"6a25eda304f7622a", x"84936cb989f89a5f", x"7e58f2c03ecb1dc9", x"2b2344de3d9ed94a", x"fd707f2f17968752", x"49be0cdc50aa5b3f", x"b43abfe912f7bb50");
            when 15789700 => data <= (x"ff600394af89aa31", x"f51c1ef8b42a6bea", x"6f33ff765ed9831a", x"2c80d8729ca68c55", x"2a9ec320921d3b95", x"15b3b24993feb9e8", x"6fcb1b7fa61b66ed", x"63d909e7c3401ac5");
            when 6115984 => data <= (x"e079740870ab3880", x"c515264339a0049b", x"8a6c851045dd429f", x"850a5c42e6d55c64", x"4ddd693eb262718e", x"a038bce18dc06205", x"9a120bb60ffece7e", x"e14e208647b184e6");
            when 14660357 => data <= (x"49bf9e7151661192", x"ad42baa116afb70e", x"5179ef3866ef664e", x"e90961be347e5f02", x"8d08ebff6f6ab0ad", x"09e077d0a53608e5", x"91f54a22860bf7fa", x"ef29a587409f3607");
            when 25314809 => data <= (x"bc8391d59bb275f9", x"2dcce3b3b4fda6ad", x"25f8396d023fc3ce", x"08b4dd743a809796", x"2b1663e9728ad0d5", x"acb8097c48f4f933", x"403aa4d082dbd309", x"c32ff907deee50b4");
            when 31147155 => data <= (x"26ad6e97b146b7d8", x"a0b5e419a7aa9fae", x"fc5893e7439a0f59", x"502422d11419b136", x"df08be0fad2a0221", x"363d9c0dd0518f37", x"e096fd4de71bf330", x"a32a4cc171306a14");
            when 20367009 => data <= (x"62b38e104d236b57", x"ad2f58f989b2c8d0", x"7063844a6dfd208d", x"1e90376578a5059b", x"23d3f96dd36f8a3b", x"c8634b6ae79699b6", x"bbcb2d8150a28733", x"a3143d4be186e6a3");
            when 6976772 => data <= (x"24618f1da99fa9dc", x"7a6f21a66d15ec5b", x"de0d543cd9e2c6f5", x"9b268ebfbd4ca2e1", x"47e81d58b4a77261", x"c03d9d203fd2d557", x"52ba177cb7461347", x"a6a330298b0136b9");
            when 33385881 => data <= (x"4c3f90fd83df9cbe", x"054046a8cd5325fa", x"aefc01c8110125ce", x"cdff57cf93ea499b", x"d1463337c89f139f", x"3ba02635456bb94d", x"ab516d30928b413c", x"4c054464b65d2745");
            when 3936282 => data <= (x"417a2b9e84184cc7", x"9fbfa8e6a84fc64a", x"197380a48d8ba11d", x"5034f76a7f9632da", x"411a779305d3d781", x"208fa31164418b0d", x"e331f10558956f6f", x"00fb356fdfdeda8f");
            when 22316248 => data <= (x"fcd2a3f688881c70", x"4bc4a36316b7d61b", x"84d2aa20edddf4c9", x"5535a906fc66ffb0", x"6e8626adc5a482dc", x"49de3b1b27d698bf", x"20c60f4067e5efaf", x"119f98c1ff1e968a");
            when 9476248 => data <= (x"36fefe29df01fe0e", x"13f5f28f76778342", x"2feb5b4acab36387", x"b4d07d5e99111ccb", x"7b5c543fa47dadcb", x"601d9883e423ae4b", x"dd1cc62c27ca3403", x"fdf9ece7380f6503");
            when 9927047 => data <= (x"fb0ef4e0b99a3125", x"8363265608a738ee", x"d146a311c6dbf588", x"11247872857dc889", x"ca2d4214c3b2133f", x"43f96a66afca4c47", x"37db4e7d0bcee61d", x"28cc2f27e5de972c");
            when 28691738 => data <= (x"fa9cd909f87695d5", x"90bc628387b7abcf", x"9fcea5ab61c47bf9", x"4f72daf153e905df", x"1cbd1a6e794355d5", x"0561dad94b5e399e", x"678a96bd56d65255", x"cd9ee7b85038a84f");
            when 30478384 => data <= (x"ce37c83dcba1573d", x"e127f3a65694f140", x"75dcc07b8a75160d", x"00b0b4227c28751d", x"61c05e634f86b8ed", x"e44270e47213c358", x"284087649d76bac8", x"97a184c0c1c47d72");
            when 23773290 => data <= (x"b2e55aa25a75ca05", x"44750d86f1e31cff", x"bfdd5c710dccfcde", x"ede25f63c752c286", x"9ad5a5c84557b634", x"fcd7fa281a09de7e", x"641c20c0c5346e01", x"de9d9f1f56676592");
            when 18153090 => data <= (x"8b6e888eaf2c457c", x"c7536405a4e26aee", x"fd514c692afbbf95", x"071602605998bb74", x"b2d4b16605a3fbe9", x"d60b6bdde551f573", x"2c88f3d54c3bc510", x"54661040d3d6e538");
            when 1598591 => data <= (x"612e35d4a3e7edc8", x"83eef7781c69049d", x"28436c0d537cef08", x"7f386ba05c09920a", x"772adb685415b667", x"f7942d9574295460", x"c2976db3aed61e7f", x"7d8629ab234e8fb8");
            when 9737420 => data <= (x"405bb63229196340", x"49e00e02cb8b3f8d", x"9a1feb0007cfa815", x"9ce3800eca3eef79", x"1eea92fd167f0498", x"1bbdd554946052a0", x"cd3cd1a3ae11f01e", x"2a7b377b671c0615");
            when 17848152 => data <= (x"760fde979491c33e", x"d3b5ae60cdd621db", x"0a37b87107e27f7f", x"67b7796b0cccab56", x"df9dac5123033dc2", x"1b07d31c9d8f79d6", x"b00ad8344fbc906d", x"97fe3e6eb4c60a10");
            when 33007315 => data <= (x"abfc9dc790eb8485", x"a8433b65486b06cb", x"40d1aa10de17a5db", x"30b47f9e51648058", x"8fdedb1d0634053f", x"8e8999e90b71b3c2", x"dca0e67db0a20cba", x"73ec0cdb452c7e2d");
            when 33385124 => data <= (x"5bcfd0c9abf0eccb", x"fc9f8bb2a7c89f16", x"cbd8fb078e34f3eb", x"ff72560a066d9f83", x"f32074a394751611", x"543c3696e4f22020", x"13cb0938df5b435a", x"49ac608391cc7ca2");
            when 12678793 => data <= (x"de0e9a5b5e3a815f", x"d1461526afec00f4", x"c6ebc36a092544b1", x"63db1c8e3c1225f0", x"957abc17f22c24d4", x"4a43df8eec3febc8", x"e867b30bc9a2ed9a", x"3418b235ea57d6dd");
            when 7653911 => data <= (x"64aa17a00dc74e56", x"c2c3353a6ca72a45", x"d593f1930afed8ae", x"0df4d62a07d5446e", x"0ee0b457a2302e3e", x"b46631ad435d5246", x"a35fe56490079912", x"737e9859e0644a2d");
            when 33566071 => data <= (x"a4435adeaea6b844", x"31937453fe0ad113", x"be3f41a5c0121804", x"8766271b2bb8dff7", x"7b96f1084c84f42b", x"6b57fbdb30dacfa8", x"38c9da6a2f48ff31", x"0d2865e0c024c43d");
            when 12732447 => data <= (x"08fab2e287b9bf52", x"61d767b58de2f54a", x"462dad8f696c3c91", x"da4405c4887e37d0", x"814c678d8a0ace0f", x"e50b6dd5896a8e4e", x"6482640d3e8a5707", x"284fbc107900b23a");
            when 15575154 => data <= (x"ad49aad6e8029ec3", x"7c70d96d4d63f414", x"8935a76f0f144f48", x"350856fd3242b154", x"717982390f7e1261", x"ec34e0c88d29a7b2", x"1b950ca719a05eea", x"0a479a595537e327");
            when 3023809 => data <= (x"93cd7712247c6f27", x"3895f2753d730bfd", x"e5a3020f8e976dc1", x"fd4f4ef12b1eb1a7", x"9f091468fe71e320", x"65cffce36b52555b", x"dcfec6f955ecea7d", x"e3ce51f921dda3d4");
            when 17967145 => data <= (x"44a52d420d5eea93", x"fb867034e6847d8e", x"e6aaac9fadcd83d8", x"8f31270e121693ad", x"c2ef34fa530e75f9", x"4211a675172da903", x"46afa7a0af7919c7", x"73ea69b98446aa45");
            when 27766406 => data <= (x"bc2fe16989ab19a6", x"8fd78e4ee94566d7", x"94a599173d945379", x"01694043bf8d8905", x"57f77dd85c53c5b2", x"efac059e1415a4c7", x"159a885fc0673523", x"e45a3e660b49e9fb");
            when 20388835 => data <= (x"7a895af4f21bea3c", x"678dd508662b0287", x"39b3045d55f9aba0", x"32f608797508d24a", x"13864157141f26f2", x"e238427671b50276", x"6f1e24c7eae06b74", x"59f9bd01ecfdc9be");
            when 31792250 => data <= (x"1a3b167027334b38", x"2f9597fa27c0b030", x"232faac75d81007f", x"a1a8efc8452754c1", x"332881f54e9dc8c9", x"4ac37467d2b6a777", x"c61a4520cc70a129", x"2c8c42e103e3125a");
            when 24605584 => data <= (x"f8b86828dd1b24c1", x"2c7a1094dbcbb6e1", x"8a1ef518a5818ec3", x"ee00acff1f4b0c37", x"116e71179b0fbc12", x"79256b5770030511", x"576a8e30641ad4ec", x"54153c1d0fed79d9");
            when 14781042 => data <= (x"afb01c3009324638", x"6f6493d1c5b932be", x"8804d8889462cd3b", x"785ed3ce2184a767", x"54acfe9ef390c935", x"edcc9c8dbd7ac410", x"98010918e15a5fa2", x"20c28909d8bcea05");
            when 5673391 => data <= (x"948bc2f995fe63cf", x"3e4422ff4271d0c2", x"21acf275a907ac82", x"b754645f3296a1a9", x"f6c85e8dfeb0b4e9", x"7fed7ae636fcfd1b", x"0213ca7d435f3e78", x"0f39f4ed3c23210a");
            when 9573197 => data <= (x"29d4519b26f8bdcf", x"065d615e53e011e7", x"eb91dbe347041cbb", x"83b06480871badc0", x"a2223a17c1edb951", x"94e72112da7ef910", x"77f5369a61260605", x"df9c08fe465d991a");
            when 356315 => data <= (x"97d4147f10f0a00a", x"f781b151ca59f3b5", x"a3d705979d27883b", x"a91283e9986c4b94", x"83c072c02b25bd94", x"78c34fc0390b7d25", x"f2bf480eeb74424b", x"a9e65f37a9cb6b9e");
            when 17669147 => data <= (x"96b9a0e8a4a3e180", x"adc668895afc94d4", x"7f1206a1a95805a6", x"0185681e3633d1f0", x"8772cf6a11553c48", x"c5ee55875471b197", x"733f51a0f069a713", x"2cd3db2a91adaf01");
            when 4634320 => data <= (x"cf268cbf8859851d", x"58df9fcecac83038", x"a2da99a2d16afe39", x"f2c397d06bb76690", x"f0a0b41f002a209b", x"7d9fec0df5b63edb", x"3b5e5d187f927215", x"55963f4ef0d52bd5");
            when 30582740 => data <= (x"80f6757f1566c414", x"1f27378aff635e22", x"34ecd503fde2e837", x"215410b1af5092c6", x"627e2c8c7dd97bd9", x"fbe45249516827f5", x"a257f7d7687f2549", x"7bf93374c000e650");
            when 1216665 => data <= (x"d812159bea84c3a3", x"8f91b528bdcc6227", x"39b93fac1e25fc42", x"88ccf0c845780e0a", x"7989e8b48af3f5b7", x"54415cc1396f62d1", x"4edb6174394f65fd", x"e98a9018d0510925");
            when 3070901 => data <= (x"ba2ccde19c20cf5b", x"63ddc3d9511683c3", x"5a7249ce39576481", x"3b5b54806497f7f1", x"1bf69a0b81cda937", x"099e774f4f837cd6", x"fd5beb4738bf26eb", x"9cc686b12d0bb145");
            when 22610432 => data <= (x"e2bf8e9e8a9cac9f", x"1cbcbf793699a0d7", x"d91e2700cd0a4254", x"58a405721d831a98", x"39ed62e386df80d9", x"882dc0f0fe139673", x"834fbc5cbf038df5", x"4d9395705f9d3481");
            when 5774895 => data <= (x"f34edd4c3d74fcd3", x"f69c2ab0cefef4f5", x"640910d72360b7ea", x"674be36ae4f8c9f2", x"5cdff6d8068bba74", x"9a27a52308498ba2", x"27a77727823653e5", x"2efcbbe68e457fbf");
            when 6921714 => data <= (x"d04d4cb7736772f7", x"5298cd3aa17c9780", x"b872c2d234808a83", x"0f71a4ffd9b23d1f", x"f9029d8615a2ec62", x"29b66359bf3d12d5", x"3dbece5ce3b1a284", x"7bc55dde3bf89f1d");
            when 11428663 => data <= (x"e37cba324f4ce84d", x"0490bb6643974927", x"fc559013e35abc5f", x"ab7e156fbea925d5", x"637189052535c334", x"c87b023b570eb5ef", x"e1a32bd368799bcf", x"bd5838df355bed04");
            when 33401459 => data <= (x"261a7a87f63da94f", x"268946752ea75b0e", x"74ed386f4e8fc26c", x"241a96cc3a69cedd", x"072691c08d4c5333", x"ae1b3c673fe39810", x"dd16c129100b8c76", x"e956f36833dfa562");
            when 7492306 => data <= (x"fa0958116e7b82b0", x"66842002d2f9c550", x"1e8b46aa2526015c", x"4cb2a6de07eafa3b", x"07ad4da189501de7", x"de4081d5eff44940", x"3642445077ac1757", x"8070e2e3623966b0");
            when 33287941 => data <= (x"ecacc9709fe33d18", x"4f591c20ad1d512a", x"458f0a85508aa0f2", x"f777fe3d6aa20ed7", x"5de4b1ea2269b6de", x"5532865db84bf00e", x"c9bb99988cb6154b", x"6ec6abe22fe16370");
            when 33665495 => data <= (x"e732d6f0f26a9a14", x"d28d68558581915d", x"d734d6bf7eae6814", x"b83bb9eeff0e1238", x"478a425fde991def", x"a4725ddedc593d42", x"6eef5ca77a69f41b", x"42288bed94f76a2f");
            when 5404404 => data <= (x"82c299f304b378d4", x"3802990d78b7abb3", x"4c68bc6ce56d8933", x"e6c94348078d365f", x"6140cbe27b51a5ec", x"818d95a1d289217c", x"f70d712649bcb714", x"83fce7ba44c76a27");
            when 29293258 => data <= (x"6500cc0328e749aa", x"7c2c1130bb05b1c2", x"c0d369fd20f18753", x"31c75e3161443b36", x"a529a5cf37d277c9", x"fd1bf3de087f0d18", x"cb3a6e5dbb7da062", x"8cea92b8d278fe7c");
            when 8331105 => data <= (x"2b6a3d4e6652a09e", x"975c3fb877031818", x"c47c4bc7cace0c30", x"a5e5f2e32dd31941", x"b88ac7e01e1fbaf2", x"70526d1b634d73de", x"789504529ea7ed54", x"11ea6f9baaa037a5");
            when 5641515 => data <= (x"a904232b15e18a50", x"a34ec2277b847359", x"27c9db64549a04f6", x"cd7f23b540852b34", x"771c7092b18890b0", x"ffb8548461eb0bc8", x"534d67c8b9513144", x"e5d75de2768761a5");
            when 5739676 => data <= (x"3bcad7ddcab4455d", x"caf104eac03f8c5c", x"33a8a1396bb2817d", x"81dc116a4584daa7", x"b3468935f5603a7f", x"da544d1d14d3978d", x"340d2e26c4435ff9", x"0b896fa95cfe4c02");
            when 21567915 => data <= (x"e99fd8160cb28c95", x"db2247f7b14bc57c", x"56b4843d0a9ae9d0", x"6c930ca33715e1c5", x"aed95c08841fce7b", x"386df1c6b680305a", x"d4de0522fd2b71c5", x"7f1f1d6836b13917");
            when 27562280 => data <= (x"8d3f866ce449758d", x"5d43ff05e0ac38e1", x"90015e2ba6bfaa30", x"84f8aca338b65fa7", x"016a58ae84d1385d", x"8f6cfaa8f42e4c7b", x"ff6927ff52c87f95", x"d21234ae9e6c4dc3");
            when 25695328 => data <= (x"8bf7da4958aa2765", x"f3b4a6553aa9aa0c", x"c23e9187ab8b293a", x"9ca488617bd5b367", x"083f6394193aa55d", x"005fc32d9b9bcafb", x"2066f44cec047d5d", x"f9c9263e97bf0b1d");
            when 20028392 => data <= (x"b41b3bbdd2b5ad08", x"67452c3bbac99a61", x"a7a6dc2a28e4dc47", x"f4c386e3f3e9a249", x"55884cc6ea9bdc45", x"3a820ce6dff409b9", x"bdf8fbd59a2b03db", x"2479a410ef823291");
            when 10315061 => data <= (x"a0f5f4e85c10ab22", x"d051bfaef79c933f", x"1ad176c4288fe1a7", x"76dbbfe461bb33d6", x"c839bac7238be1f6", x"5ab5365f04c4455f", x"660de3e89dfcb8bf", x"2aabb5b9f14c5996");
            when 33225376 => data <= (x"2a103171e3b30a0a", x"d8a4fdffe62d3a8e", x"0c71cccd426d3060", x"00a69489933d737c", x"d925875b057a55da", x"60341bbaa95cb273", x"98f397aba49bb308", x"13b3194f0dd6ee46");
            when 22429701 => data <= (x"6ee2666a4c6db969", x"07132b464c98dfe4", x"451c2b41bffecd54", x"79a95179b3a78e93", x"293bd2286dce3b89", x"dde3ca268d20cf8a", x"3db92a6d87edc937", x"921841e866739073");
            when 27797394 => data <= (x"6dfe0e15f6f928db", x"99f7b5e3310ae61a", x"5aec2bc8cc6c4ad1", x"65d9a62217f05855", x"80b45078db0b5fae", x"c790b220190637c6", x"e1674ceefd6a511c", x"16f1ec15a0b9f77b");
            when 18965054 => data <= (x"9cbaba395bd8fc7a", x"a6606d0107fb72ae", x"a04b7aec8cac9043", x"de09f03208c08bfb", x"acc84e8707335c5e", x"4f6518deaf131149", x"2081455d479e6b53", x"c779fd4bab61f84c");
            when 15611891 => data <= (x"b5b8a9970231a55c", x"792ad97c70a72aed", x"b55eac7f5ab84852", x"e332028c8e8fccb2", x"0faeb82c42f36e66", x"95f3f4da2b876ad4", x"202e017df73aa0ce", x"5dca37ab48517919");
            when 8402993 => data <= (x"cee752d4f26a31d3", x"20fffaae0804996b", x"dc3281b946f6aadb", x"b8ba9ef50913a16f", x"8669510d67ae87f8", x"c99baa0a5c8f352b", x"995be34a71bf57bd", x"2325e37e6afcf414");
            when 23746816 => data <= (x"89849f24108da9a7", x"f2e5cd552826bb56", x"56144420a3fae3a4", x"03cfd17953d3cd51", x"5e5d11699c41cf2d", x"a31f591714ddf6e5", x"492c97e816430630", x"f538df00faca0e60");
            when 9224382 => data <= (x"4ef8f55644e8385b", x"f4c5218bdec3b684", x"98ab88acf86047db", x"7656c811f11e0b15", x"e759b91cfee8b32d", x"46470f527b33e291", x"cfdcbb62cf93c872", x"f54458b2e855b1ac");
            when 9364651 => data <= (x"a71852a05f71ceb9", x"a319bb35935ee5af", x"c3a0b615b6441010", x"49ec72aa5069055d", x"d38a177c868bcc6d", x"e2ed4fc63e0b6e34", x"ddcca2972e4226f8", x"a508bca1b5930036");
            when 7293524 => data <= (x"a4f4df6677bf87b1", x"9cda0b24c32ca257", x"dcba167e854e1925", x"a736dffd47052e51", x"0635e1e298561ba2", x"f8ec804838c75f8a", x"a5433083f9c27177", x"c0db004544bffdbd");
            when 20646840 => data <= (x"02430dcbfe2afcf0", x"c9b13257cd3d0527", x"874de510e3c895c4", x"eeb9049c53d7ca1e", x"3ed483dc35f35c7b", x"663bfa0e28895e18", x"e2576fe492705eaf", x"27963258e5157988");
            when 30483727 => data <= (x"0b3cfa563ddc637a", x"2bcb111f20d47003", x"3371322597055afc", x"3d48837fc01ab856", x"f1f34208d9e650b4", x"e47aea7f2d8d8443", x"ee4ff432f2a504f9", x"7690eb500442c028");
            when 5591934 => data <= (x"4a7c3d0862c9fb88", x"f52726b7b9f1ddf1", x"6490826d6737ceb6", x"02d8fff524ece3eb", x"2958d5e1634ad49f", x"72092d68cc5c7b7c", x"f0465939d9dabeef", x"20723171778d104b");
            when 9711248 => data <= (x"2d6d71e747530ade", x"ca565b6506ab0408", x"39a46c2ef244f87e", x"d795c9bc27553246", x"b65d8d9a19ffdf74", x"a4f420694ae0ef8a", x"e6eee5daa1a2c09e", x"cd894faeeea20ee9");
            when 3289901 => data <= (x"9db1b3697de084eb", x"669c91c839549396", x"341cf825997f0a97", x"82bfe557614043d9", x"b968d802a55bb4ec", x"4f89b902577f1577", x"7456ec06fea45f12", x"000a1746f5939dfa");
            when 24142153 => data <= (x"e20e046f1f147ff2", x"f962989f4a098032", x"95a68633cbc8fe24", x"6c88279ad384477b", x"93c7cdf43cc7b69a", x"c3512bd3f07aa3a4", x"d553aeea1caf675c", x"16e094fac7876053");
            when 10739615 => data <= (x"06e7374c05080741", x"28226885654c52a4", x"3424140871248206", x"3c6040062a81364d", x"b45531e8b2a0d6a1", x"b99f487b8d4d8185", x"467c6d207a258cef", x"08d74d3133612523");
            when 1313491 => data <= (x"3782ba5aa0ea2060", x"d08977dd8c2510e3", x"f1bd971e30ba2d1b", x"1c628c1e9e1ba7e2", x"d162a0dc91183a38", x"f32ee92f384f2d51", x"f72bfad5260204d8", x"54d4445c018cea75");
            when 12481436 => data <= (x"5a15b335fcc33e2d", x"8ca54ba43d72733c", x"ae9d136623fdf8ce", x"192ba91c2df8f6fd", x"14b27770d98ccc96", x"8a8cc483e7091f52", x"fe634d8831fbbd10", x"0ac29778936cc27f");
            when 15551029 => data <= (x"9fde1c675c8d3e6e", x"2b5b578fa15efdf7", x"fd3c9de99c4c2352", x"9fbfedae287fc35b", x"ec9950b3633463b2", x"6aa9c28c4d5e2694", x"9694b654f0185685", x"255937bcc46f556d");
            when 33372977 => data <= (x"e38a53321eb2dbd0", x"a40c561e54ac6ed5", x"a7ec3bda4c6639f8", x"265e6524ff40b635", x"cfd9637b1bad4a6f", x"3cf7a92b9ea9ec1f", x"bfb0cdf9c481c1df", x"74598feafea8bf52");
            when 26534390 => data <= (x"62601c7e3c87656e", x"3abe8b40831fceb6", x"17b350f02a715d10", x"9ac9e6a07ef6561b", x"cba1c4d6b89e4aa2", x"272066219a0394de", x"85c3a024581f7d17", x"c4a0b3c5e740d436");
            when 27928873 => data <= (x"63d4cdb4522fb984", x"0022cf8dbeae2060", x"4713bc19adf2aabc", x"56f0f5326c43101d", x"3b3e848d01813761", x"c037c40f450a73e3", x"015ee6b2f5d640d5", x"ada9fa6ccc2ca44e");
            when 7402467 => data <= (x"f166807dcc254c83", x"d2bf145661bbae98", x"03c768c4b802ea2c", x"b55b62e1c92506c4", x"c8d97a64fc365c53", x"31ecc9ead21eb35c", x"7d526d14c2175d92", x"6eacf1fdef379b14");
            when 22584758 => data <= (x"92c021c01886006a", x"0bb976427313027c", x"182f778a75c9a9b2", x"d594aa54f1c13497", x"f950fc463df4f45b", x"e7718adb1ae4765f", x"c24ae47a464eea46", x"9ae4cc3af7351d0a");
            when 11831290 => data <= (x"3fa80aab5246ed76", x"11e87078ca65d604", x"6b448b5dfd4a022b", x"791e0c5cda60d048", x"60261a085ffda22a", x"d2f57e174649a48a", x"e72d980eb8002217", x"3f242eff03fcea91");
            when 22694237 => data <= (x"d2453be070a13c66", x"a064111247d45f0c", x"58111e22e81286a2", x"b6dc3e126079f1c5", x"525b36289b385dc9", x"95e5cee2d78a4577", x"2ab302a0e62c8737", x"e8dd121a020307c8");
            when 11421487 => data <= (x"a771e079354228fc", x"0f8777a88e5bf913", x"9d948276ec8f6ec9", x"416159fec2fc05d0", x"6433d87580ddf22c", x"b1adc0882e0da841", x"dbc0730bf32deb9a", x"d434a4636c167797");
            when 2119675 => data <= (x"c3e44873a2bf1082", x"70dc5b313c1e3599", x"7e863203f73d482b", x"648ca2c76e5991dc", x"8e2a254b68c00c4b", x"3ba42ee6bebdca12", x"52f87637363bf879", x"e53600ff786cfc6c");
            when 31629783 => data <= (x"e8c540b3604066d3", x"cb59d1e2d47aaef2", x"f9b12faa5c39a0f9", x"f04e44f8462942cb", x"33a8a4a3c81f32e6", x"af094e740ba4b85a", x"7682d8ea12d547fc", x"41bbf996deba6e3b");
            when 14638112 => data <= (x"f867e7f0aa86e778", x"41518050aa59cf88", x"16049a6ce3ef0c8b", x"d68ecb7e11d773d1", x"953c42ba8c2f029e", x"c39ee9809bbc5a92", x"9545146ca1cc8ad6", x"550174bd3328dace");
            when 30292120 => data <= (x"d869a88fb66c2f11", x"e48bed1f0dcb01be", x"abcd60c2d6217b46", x"c8eda2ed2dd601b4", x"3f9de0babe694f41", x"6b98bb1655cab4c5", x"b3fffe57226fff87", x"afd38241b7d8d248");
            when 33556214 => data <= (x"b3eddc8a3d5e7ef9", x"4a0d2e9c222ea1a3", x"2eba5dbf75e3951a", x"a4fbbfda5281e1c5", x"5040692e7f8314ed", x"510d68498f9c81e5", x"d0754031c0bf4c97", x"51dc62c1169acd77");
            when 2999447 => data <= (x"c8620a98e817c2e2", x"a8e4d0a50f1fc893", x"45d8ada9bb122796", x"88bd9b2de0a06d9e", x"86cd885089ba58c2", x"a09958298bbd3d90", x"675d8eb7f74277e6", x"861254f65254a8dc");
            when 14149228 => data <= (x"89d8244ce0d4f87e", x"af35fde393a06346", x"9e32a0c7d4d9ef6e", x"28353f1eec6c7a5e", x"c6286e9509362e7f", x"fbec15f422288bb9", x"bc826adb00d47c34", x"309028835c5cbf6b");
            when 4724950 => data <= (x"303ba784dbd1295a", x"cc8988896f19544b", x"71c0c734d16d5ef1", x"e8c425dc29240341", x"2adf2cbd112e1432", x"f79b2fa2ef7cb88f", x"da3c86efb8125ac3", x"3ca70cc0bf27b822");
            when 10032684 => data <= (x"b48d5d269c1cf5f5", x"e94fb9c3943210da", x"0a8b467f7f1c210e", x"666b6a4e2c9ff71c", x"39f9a52477d171a8", x"fc26bbfc3420c5e0", x"355f2e39961bde75", x"8d437f2750a27d07");
            when 23646218 => data <= (x"1ddce11593095659", x"721741df604e032c", x"8561310eb94daf48", x"f4957a0a5ea3f941", x"4282610aa796cac9", x"05d2f75fc57aa86f", x"394bbf4be0f6b34b", x"07f2de43dbff7471");
            when 8993449 => data <= (x"56dbc5d3f4dea8ca", x"0204ae52d0c9d364", x"9985edda11882abe", x"2d9a1fed79c4df07", x"9ea5caff9a39db6d", x"bc43f97f0d539c98", x"5ca277b9a100f3a6", x"d4adf74378b97d69");
            when 28817465 => data <= (x"505de7708840caa9", x"23dbae3680746b56", x"9be8d4e25627c8b0", x"2663cd64be9ac1ef", x"2cc25be119e0eb43", x"df2a0fca0ea284cd", x"c10eb383ddb9be6d", x"e4a452fc09382df0");
            when 18319193 => data <= (x"60a10941ebc21e2a", x"ca4f556e1735ab34", x"7cd27a690f35e601", x"ff501106a70fdbf1", x"ce01aaf415a4653d", x"47e98133018a043f", x"85acca9d88b77b55", x"5cdf66d4f66f78ab");
            when 32442325 => data <= (x"7ef005c1bc35028d", x"a485f30501014dbd", x"c9a5f93168b2a171", x"39e96449e68cb657", x"ca3f52709b8f7748", x"2dd635b1f1cf6114", x"cd1931d056fc888e", x"9addfeaee0787073");
            when 32080613 => data <= (x"4e43dee17d86ff4b", x"bc4d286be4219db7", x"e64b3d078c4be729", x"fbabb34fcc7cef29", x"bb06a1beb5e6ef03", x"a897aefdf5eeca3c", x"7e034aae74c9f482", x"991be48a7967d4ef");
            when 13146145 => data <= (x"717c29dc1bb4e720", x"2782e47cd8348074", x"733f1d66d85146af", x"7d28b10073ececdc", x"2168ea379fd3e035", x"a83635cc57e67bb0", x"7e703c7518ce9ea6", x"c8d04c819b683f0d");
            when 24751137 => data <= (x"d3fe6d4bd016efa7", x"bf7e22acc9cd7558", x"81c2023c5675fd5a", x"1bccc93cc6515e65", x"505ae2d7639cf327", x"8d0a4dfe5012923d", x"9d7245b514debd8e", x"1b22d592e031b419");
            when 32699457 => data <= (x"3249fb8b048737f9", x"cec251d7df6e9420", x"341d9ff51ac68eba", x"989f4f0426361fb7", x"5fb669c0bb135fc6", x"5d2c7bc063ac0138", x"5fad13d1d9b93b0b", x"868beb5512e7191a");
            when 18014276 => data <= (x"7aff41f7749f9908", x"e7ca6d60d80f13d9", x"1136df4403604a03", x"abbed503368c6014", x"08ad01cc9f4cc94a", x"c27a75e7e9c74bba", x"4fd1b2fb90164ad1", x"c62ce960453034db");
            when 12731768 => data <= (x"a8c0dd6f00221f04", x"54bc966bde08fd0f", x"1a3bc92848ce7de3", x"0bea516be84fbb09", x"12a20dd95b21a16b", x"88a6de1b1ad731d7", x"ae206147c94d9e5e", x"7fa7f7072678d46a");
            when 1833137 => data <= (x"92964607bdb746ab", x"66941deab1cc642b", x"5d3e1a81843e1542", x"60de66cbafecac14", x"614a30b63d81b61c", x"25919ada01321c62", x"b449badc449361b9", x"1705091285f55d9d");
            when 17062205 => data <= (x"047a2882b4b3d55e", x"2570a6eb0be7c129", x"41620a56bd93d344", x"c94a6d2a48905492", x"308668a1a5e98030", x"01498db5eeac8e0f", x"7fd647dc3cfe2d88", x"f879ad2393c4e71d");
            when 1736043 => data <= (x"d1ed555ccd919cc1", x"23a135416bfde427", x"6d66a89e711b4209", x"93454c9243104124", x"16e59d93f0d55ba7", x"cc30d54fb0ad0bd6", x"634a9262a511985f", x"e289c08dd9aa55f6");
            when 31228681 => data <= (x"f56bd59a382fe0fa", x"792e944dc5ead6dc", x"73dbf4d566849b08", x"bd958c677785e478", x"c8b8d899b6b183f1", x"e6a556ea24199183", x"b7a4c3acae19b76e", x"530ea2cd3fbda04c");
            when 23231368 => data <= (x"f6809bd626e0035c", x"ba5da8e312971012", x"4658016a57acee01", x"d173daa5c3d3486c", x"f05533ff11fd4601", x"0ea0a034fffd85cd", x"c9316d523f7ed2f1", x"158cdd45a5f52468");
            when 24584106 => data <= (x"8c988cfbffe48a50", x"b62a003f597bb403", x"db623d43441002d0", x"86a2e00b2edfdb9c", x"a218d8f2dfb35e84", x"5d02578e15c4aa1e", x"e25869b014dfdadd", x"9660c1fcbd57d078");
            when 33214404 => data <= (x"f6dc5865b2180dd1", x"dddb89dd6cf053e0", x"78d817403ffaf631", x"004bbd77f30df528", x"24e2b8950ab6eec2", x"0e8b5cc65f4bc52d", x"20c1952a6039ddc3", x"f0ea5dd6f4959470");
            when 14201436 => data <= (x"2ea13aea2cbbf42e", x"e7856ab650db03f1", x"2a36871c41b6fa11", x"ff2f865809c89c18", x"4627d5ba99c60418", x"33015bbe302a3bdf", x"370b80e4a1a06f53", x"1c906b624ee2bb69");
            when 28183213 => data <= (x"7200ef7ee6feb554", x"da387cc66f021a52", x"a5863e6eb8a599d3", x"b37cdac6c631385c", x"0b69d13da332161f", x"74a0c960596431a7", x"7c5f853e463538cd", x"7903c69aea82f8c0");
            when 17806881 => data <= (x"bf36b764fa58fe01", x"e577d0194a46ec1e", x"59369140cf703fa3", x"ef339aba67c929b5", x"dd32d1f5c2378dda", x"49d4db4c6dc8b6cf", x"04b9196455a2b63a", x"04d0b1d03297f1a2");
            when 21750385 => data <= (x"e94b8f8510ecc113", x"9c4a47530e16a635", x"fc831a5e81e5fddd", x"c2d4a77cd712e660", x"0e70e9c383f1c20a", x"5bbbcb94b336958d", x"6ed067d8d751fc36", x"9cd73cc8c23956ef");
            when 18762731 => data <= (x"3fc5fd0b322ab9f1", x"6ddf10f19a8559ab", x"b12ad686b6a1705a", x"0efc4cc543fbe1e0", x"134f0cddb49cf54b", x"ed5c25e48322fcd9", x"918c53ac88ae18b5", x"785ab8082fef8ccb");
            when 10918793 => data <= (x"abc86ab5c4ca54b1", x"b101df55ca17f4aa", x"2e4954b30fe94452", x"60e922bd1d270aed", x"caff681c20be2dee", x"3382bdf597dfb5ae", x"f0dfa388185cb3c0", x"e9600f8f24fb3c26");
            when 853227 => data <= (x"3e943f6b9467ced0", x"b1eaf4e865db4165", x"4f5a1d86c4855cfc", x"e239a5fd309bd75c", x"86870f3f7c3a913a", x"4607c4d40f7ece8e", x"b0aefe59ed6ca47b", x"17504a6d33bdf779");
            when 30931954 => data <= (x"28170d6116f879ed", x"c1f2867e55274655", x"93a4bb050cabef20", x"1a69233d94243cc8", x"5965580008e0f4a7", x"4ce8d2a9b09c6a2d", x"ae75ac2a02a209cc", x"dd6841488d480ff2");
            when 33037769 => data <= (x"78ca74fb8cc77428", x"6442823a86dd28b4", x"ff591732fa9e859a", x"c65adcdc006b568c", x"94cafedfc9811c1c", x"7c3a9e829f6c5bf5", x"50fa8d3320763da2", x"855ecb64bc6ce988");
            when 7266138 => data <= (x"30a0d9f61f0b57ac", x"eebeda3e45426f91", x"0cc291826628d71c", x"500cfa74018c35d5", x"e944a15d0883521a", x"c0de89106813bece", x"266582dcb8f66d38", x"9073ddaaa660cd7d");
            when 23261456 => data <= (x"8bab4bd574d012c5", x"c13ac557bd0fca11", x"48d6cb5a2b31f51c", x"230b123bfea9836f", x"ac762fba3351a81c", x"fa08b0e1fab15f3a", x"291c050f826d0c2f", x"5a3d8dad914fbb53");
            when 27061733 => data <= (x"d2ddcf4a66cda7d2", x"f6ff822d3e42f7ac", x"6620dbec5ca9e433", x"891196f821399dba", x"203bbcb3a98ceaaf", x"84fd69c85d334351", x"0a686a52932cf83d", x"d915dfbbf147319d");
            when 6971876 => data <= (x"0844caaf5bfba29b", x"ee3408098956fdda", x"8959161aa95eee1d", x"7efaac3600af26bb", x"c52a0099c3e0a392", x"268c52ae164ea6c5", x"6c4c907a7f2926e7", x"28e450d35b9b292c");
            when 11678635 => data <= (x"18a01d0de5e7b691", x"496913bd8ddfb598", x"814bc70ab0cec155", x"b566fabbd758f9b9", x"c492b40b3e85c3ec", x"efc4a63b41a19fa4", x"d9366e30633ece0a", x"ac63c1a59bc6fa9d");
            when 25177565 => data <= (x"407eb658a8a586e5", x"7f3f6df1c5348650", x"0007bf12ee448b7f", x"b0408e3dd17a429a", x"256795b659294b7a", x"e7da471b6bd9bcc5", x"1f937a0e72b0afd5", x"059a2eeb4a3521c0");
            when 16035547 => data <= (x"2eb355400e1d78bf", x"e7e94c32a5010c91", x"20adcd6efc679312", x"abe030fb3e62e345", x"3ba506b006ddb50d", x"8051ba8d17ea2900", x"b42d8995c1b16faa", x"9f84f9167da3978c");
            when 20712525 => data <= (x"ee1e5e782a7e59f5", x"ceef85bd5064dd54", x"dc69efa0867c9303", x"0e4c1249c4af1250", x"f60f293f5b75c145", x"ba4fdc5f1fb0094c", x"5a74f938fe3e25ba", x"47f30eb1d2dad759");
            when 31069362 => data <= (x"7f06f67731e92c73", x"32b09c576ca04151", x"89a025f933e16c32", x"221bfae15fee8c2f", x"864f4c8966734049", x"faaff9008d15dea5", x"3018804c1eba8c08", x"d6a1c3d14cf77997");
            when 31490419 => data <= (x"ad95b4c399c95940", x"cdedebe8ae10e579", x"6e86fe00d1caeeda", x"b2c1db3dd5d5abba", x"8069abd90dd9951c", x"292d3161e47b4810", x"5e10893528ffa5d4", x"f23e49929bd6f800");
            when 21637529 => data <= (x"36f29d7e50b621d0", x"583b6bad4c5ff206", x"5f74a22abc55bf0e", x"26a3222e299ee95c", x"0ece206211e7699f", x"9b67f939dfb65487", x"fd61ffa9ba05cfcb", x"0c52bd2f883e735d");
            when 3821893 => data <= (x"0795d07176420d18", x"6b6e3b99e52ccf8d", x"20d0991b06e41148", x"fe9d02279acbef29", x"d371d273b83b9a55", x"5a8a23573707f0bf", x"7265c8ce5ec8c4ec", x"7162ea628a52c57d");
            when 20156895 => data <= (x"54f931d08e3df8eb", x"1d909ffa4f8377f1", x"bf60bcc2f703c562", x"9f76c849b6192d02", x"f787f9eb3c1bb415", x"ab146ddec5de309a", x"58625444bcea4ffd", x"88fc7b03a2344659");
            when 32995440 => data <= (x"6ab33237650e82b9", x"112e521498d8c49c", x"3b634213267a77f5", x"65e812cc859391a5", x"142f9f4f7e119cb3", x"25cb13b63dc4909f", x"58902c058ed59ce6", x"a7f5097685db96d1");
            when 20325981 => data <= (x"5db410ea3bd39270", x"e0b1b6f55ffee7c4", x"35aa94ac9f8c21b8", x"3291ec23c15f896e", x"c7e7f352078ceaaa", x"1901b95545f85e8a", x"24af1f8a289e87e6", x"e72ba2a7225f1ca8");
            when 528633 => data <= (x"4297f2000ad4d757", x"71d0ff3915d9e3cd", x"5c77b0e9e2e83116", x"4d0156ac2b7ffbbd", x"19650af2b601ee22", x"7ef538a33828e646", x"7d804a2861c576fc", x"ade8c8ccf49a07d6");
            when 27391283 => data <= (x"1b2e784fe10f3a6a", x"3609c4493d5aca08", x"1449d8ae5dea87cb", x"e6e00f982f49dc55", x"80e0f819f3699ced", x"0847d9821e16e96f", x"3cd2359a01f534de", x"8cea665e8e43cd5e");
            when 29270643 => data <= (x"11241d8cc4959790", x"c5336f5f657ecb2e", x"98e6aa0225432751", x"24fc7d4b07af286f", x"9008a606e5dcd5a3", x"28a18d7573c374ce", x"7c2c3bfd0a455424", x"cc4585c2abe24fc4");
            when 16252158 => data <= (x"be35c605e7499d63", x"a236f56a0a352c22", x"ddfd9d9ce5f09d50", x"3ab12bb62ecfad4e", x"1e3feb40e7561cf7", x"d411cc50d9b90878", x"53e52321b9256da1", x"7809f42e173f1bc1");
            when 7503570 => data <= (x"0c1a365bfe3b30f2", x"2a22bb5e0f6354e4", x"3b0d2731e23ab9e0", x"551e61af4542a8e1", x"00534e88e780d210", x"39ec60d92c98df5f", x"df43249a900731a6", x"56041053884c28b1");
            when 13234299 => data <= (x"968fd44c5fececbc", x"8ecee72f218679ca", x"fdc85734eed20031", x"255385aa630f25d8", x"04d7c540597ef90d", x"068caa9038eb8063", x"4be43e17a81b18ba", x"145ec5e51985ca9f");
            when 27976553 => data <= (x"92120aaa603f39b3", x"6e6beca509f9a51d", x"ac8af6ccf0485a56", x"f8691d0aaa9d64a6", x"690913ed4760ec3e", x"aeed5f2fd3cf5096", x"183cf0b24ddcbe6e", x"e08379b6ec17f61d");
            when 8048441 => data <= (x"43c9f08a5f9a2e4d", x"903af86f3308665e", x"5ee61223e867975c", x"e7aa13af17d10039", x"90d6f27fb84347a6", x"5a630231fc56ef49", x"a54a483630f0f168", x"205e02a355111bcb");
            when 8178377 => data <= (x"eafe64654ed867b9", x"c56feb122c59e881", x"00090c0a3fde2a4c", x"9da1bcc0503356a2", x"8c75d461ba97b637", x"ce207af26a74bbfc", x"d3bede1ee50d5478", x"3cf672939b2e7a87");
            when 17719880 => data <= (x"91c322c29679506e", x"db8bce3104c2c90f", x"2402184c587c0343", x"c5c901c9c67160d6", x"ab80f6db256c8640", x"a44ad0bef5f01665", x"517599cc51d060f5", x"8700487106d9576a");
            when 18340285 => data <= (x"4e2921d2a8c580ed", x"108003d815d0d7d2", x"e7a270c86d0872c1", x"377e59b928db9806", x"1b6f90875211ff78", x"28536acf54d33cba", x"5d6d8a4ea8af8463", x"06afa94b0a2e2839");
            when 19547008 => data <= (x"e7f7f9486e1e5073", x"76e9a998f6e40eda", x"7c12bd7196ae5ce3", x"ba39ea86b9033b28", x"8f085800f710ed4d", x"e2cd9615773e6bd4", x"8787fbc421320862", x"83b2038ae1098bf2");
            when 31339331 => data <= (x"96e8d7d85610a3aa", x"d00ba06b654a8172", x"96a93e1875dd4a82", x"88850edd24bd80c5", x"80479cfb682216b3", x"286e7a77eb4437b3", x"3c23770df68fdcce", x"e6d32ac68b1d0dad");
            when 28045265 => data <= (x"b7bfb50c2aa2cf5a", x"026ada80b5a28d9e", x"40375c8ddcf12092", x"cefc34759d6a1511", x"f6b799cee99333a2", x"09e97d5dba0754f8", x"dc219148cf3fa85c", x"e6ecb8989982475d");
            when 7087257 => data <= (x"20c53257c5875c8a", x"f006845446d0f421", x"eaa830e432343c68", x"59647202d0b01675", x"ff24d4b59e804992", x"48b45b4f312669b0", x"ea252470a26db5f5", x"e62192bcf1e0649e");
            when 30396159 => data <= (x"73496b737baea93c", x"2088f0d088bbdc89", x"b94da759a5c52f1e", x"92809d9205c49646", x"3a5b29cfdd126d84", x"3eaae0e4770c9274", x"5ab8ed37c6f5408e", x"af74689933a61d38");
            when 11196846 => data <= (x"c39d45ada1568eb9", x"8b740fac483a879a", x"bf3f5b10bb344854", x"b7dadb78d693ca40", x"c627724f63e5be44", x"ca6cafb0cbf6f2a8", x"d246cb90492d51b1", x"25e965fda04656c1");
            when 15613910 => data <= (x"e85db5472b24eb1f", x"b4cd6596809f8a20", x"e4e8ff0e3a818ad1", x"8a49768077243ea8", x"b1ed24bf5c81573e", x"4d8723404cd30dc7", x"af5ecc81b0fb86dd", x"b4ed9a2f78372c87");
            when 26577227 => data <= (x"51162d25fafa8a24", x"9c4caca1ce063227", x"cf6f894b76726645", x"3227fc1eb43cdc85", x"625af8459031a4e9", x"6e71e932a7da46e4", x"48ddd7b90ce0803e", x"ae49c8d7ba04e464");
            when 6863881 => data <= (x"6372461ba0ffe32e", x"3f4faf72a0569d34", x"095877bdb67abb0b", x"ccf244355b993b61", x"77971af6d62e9793", x"cc443d916ace046e", x"7d37c37c864e5965", x"4b497d4bfdd0c2ed");
            when 32582634 => data <= (x"42578cfc21089c58", x"28327eaaac812c11", x"b4eed1bba09c1287", x"ccb7e1fa215aface", x"2288cee65eaa2aec", x"b8017afac8d0f411", x"dffce0a5d0c86665", x"0bff929c87578b6c");
            when 21602832 => data <= (x"3e84d9f59024806f", x"7b30e8e38ce348c0", x"e78c365989a3dc30", x"ab6432969f09bfa1", x"0064c43fe2e2199b", x"c91754807a850169", x"deab78db4c35440d", x"3279f34242f3f1ad");
            when 17700933 => data <= (x"f31f7baf014e1e57", x"6b556caae3efe0b5", x"cae8d0bbf37b4843", x"65828ce70774266b", x"87690c6f63eaa90c", x"7763dd610e5d228b", x"92fc2e1490830bfa", x"dc3025f42c694145");
            when 29742192 => data <= (x"ab17a889a66d6409", x"62289e863947e231", x"3ea7be9437180b71", x"1f5bfe0c056558c2", x"97d964ec3041155f", x"39d415056172ed53", x"3301abf7551d82d3", x"68633119f7ea23ab");
            when 15836196 => data <= (x"3860db11cc7fe60e", x"a64f717a358640a9", x"0255ed81cf43c7ef", x"8b14504f8b1d7c6b", x"4b4cd41d8fc0bbbf", x"055fc6d700c5820d", x"65ac073b6c40e091", x"b09e9b4f9e6c2df2");
            when 23975761 => data <= (x"d18c89e17faf13b7", x"bd5954c6c143bc17", x"82d05b5d75b76ae7", x"4e9fc0dc96d4742e", x"9bbedb1c848d9bf3", x"5adc4e3bf0556407", x"08913e5da5127462", x"6fcd69bca3df2f8f");
            when 28870812 => data <= (x"8fc416b6aa482a2a", x"0dae50b4b1d30ca2", x"4cdfcb2413d54731", x"f593f8e50a78435e", x"7c8a8373f93ef7fe", x"d26df4e42b660ccf", x"83e9779b77c8d265", x"5e271fa5fd76efaa");
            when 1937051 => data <= (x"c898d1d2c0dc1bfa", x"bb7895be88596656", x"8a15caa1f11227c0", x"47edfed1c04591ea", x"2bf74f877beca8c5", x"09ca7af617a472fa", x"9cfc87296668a6a3", x"7effecae2d6ff220");
            when 6236276 => data <= (x"177022ddad6bc4b3", x"8f28adfea7ae5029", x"1c7680305a88f8ad", x"2e45da01b3fba878", x"a7cbb1aa40e9d575", x"cf1f1d649aed7e88", x"ff12525213451ef1", x"593681458ac98754");
            when 27765004 => data <= (x"d92fd17e72d67b0b", x"ac61a5818217124c", x"367e522b37a6bae9", x"82a46446a013cd20", x"6c44e414611bf9be", x"8d37eb5180e18ff7", x"f9125d6d3878dc5c", x"10556e9de701feb7");
            when 17559468 => data <= (x"049222e753ae0ff8", x"5ca28d5dddf50d92", x"a19747f38c24ba5d", x"24cf7e207aa6be2a", x"61afdaac9a51c5c6", x"44a677442c806725", x"0c8f0ccb0a67eb1e", x"a678aa6a38e70b49");
            when 14543948 => data <= (x"2d88ee05dfaf1dd9", x"72e0574cca5a3a09", x"c64e7b0a9fe56adc", x"f676a0c14b3a238b", x"67df8d63361b4f53", x"f6876dadc2cf28a1", x"f737d8b6430e8cd4", x"9045a07db9616c36");
            when 3592794 => data <= (x"8c96d6433dc17190", x"d0727ccf048919bb", x"1a6ac7ddb2864dbf", x"f078792dc05634d5", x"bf5c9ce54fcf04bf", x"d549e3279e514c49", x"3bd92c7d89f0b52c", x"df17c42022c4ceec");
            when 24647067 => data <= (x"b8260df364457d91", x"259acf9635be855a", x"e3f2799de3edeca1", x"ab6c4aecbae4aff8", x"377aee30e2d0bd8d", x"8c7abcf9d8295c31", x"1e8ab2d37f18abc1", x"aeb7d18a5872cf92");
            when 9694772 => data <= (x"b665b8abf457b6ff", x"ee84724836e49132", x"536167c8d3c823a1", x"f308338898a58320", x"dccc0eab1b16f7f4", x"2a9e1b69188613c0", x"73a371964f648a17", x"32133776d33553e4");
            when 4066548 => data <= (x"f0b6f33de847bd4f", x"51dcbd284c78b539", x"61af12a159138c16", x"97125d963a9dfe39", x"8bcad8e80270463c", x"28f432308097260a", x"090a08a574a8e0b9", x"90a35e23ed62ea32");
            when 9469271 => data <= (x"0de2bcc38d9b8e9c", x"ac128cc237252221", x"984a9f1e0099240b", x"6ecced57ede5f223", x"63689457b9d2997a", x"56576bb97e2d420e", x"638f52627a9f2bee", x"ae3a3bf3ebb1a057");
            when 15779040 => data <= (x"2b8edeff1dd2c560", x"4452b2762abaa72c", x"2be5305a6f23ea83", x"0c2f4311a99a07ae", x"7731427f4822f2d1", x"22f7d0d8857f81ae", x"a191b9f2de6cf762", x"623cd8dd20ec9470");
            when 27487581 => data <= (x"2ab630f703eaa054", x"0fb5ccf837eb1e15", x"873725af5244e110", x"8679548e0ebe9f1d", x"d984b0051ec05af7", x"c6e3c46632bcbaf9", x"58dcacd36c330e75", x"bcf00e6fd41e94b4");
            when 16752565 => data <= (x"62950ccb6cb1bdbd", x"e149b8f2449384a5", x"1561640970936f73", x"7553600f94a44df3", x"0bcca0f76c738539", x"128b00d408737258", x"58a64f082d0bc589", x"af1e21d8bab56566");
            when 3371419 => data <= (x"788b4b85060d7406", x"3ce7418a98688aa4", x"7816030cba21512c", x"f67e3eedb8736c38", x"43c2274cf419f020", x"c93b1162c3c8bdbb", x"3a350052762f6097", x"32302d7f212f3081");
            when 19690171 => data <= (x"2f5772ccd295e0f6", x"265535ac970cd347", x"73b04b12276e2a51", x"45082ebbc01df251", x"4de4ca0091ff0162", x"2ed2ff98ce6e656d", x"36d7084a32ed6e9c", x"1cf73ccb37600268");
            when 4887305 => data <= (x"ef721eef0ee32d9f", x"693536f49b095936", x"52ba616fe85c4891", x"2ae04da5fa9f4133", x"20ca5551c7b78b77", x"f857820e57424186", x"e92bc513ace2b6d4", x"5d871cdf26cfd92d");
            when 989889 => data <= (x"8cf7be39b62ce347", x"3c38e700642e8207", x"7dfa2dc003d01488", x"bf92220b63777b0a", x"887846b8222457ff", x"5160902b2a3b54f5", x"6533c04ed78d371e", x"15c177c30f0676fe");
            when 21750242 => data <= (x"eb2ce85aa77d1186", x"cd269c4c2c4c86e9", x"b3e1641a2b9d9fd2", x"1a06cc7ae54fb214", x"3840baeeb86c08c0", x"47da7ef2bc1ba846", x"b9f0c16e32516ccd", x"96e204ec6d847b47");
            when 10462518 => data <= (x"832aa3c429008958", x"49de253bc549b637", x"4bc04730a0c472c5", x"4af4d3a828fdf1b1", x"72c3679042f8959c", x"4dc7adc4b760a6ce", x"415abd9ed01e5ea9", x"1ba1b3737f0afd57");
            when 31817889 => data <= (x"9429bf833284d9f8", x"eca245665c4b311d", x"b093e5f3c66d2223", x"1a357d425c6d224c", x"a307803b99068c41", x"dfe81d99bacb0935", x"dabf12baf537b181", x"c4f5c43442c1b09b");
            when 2816967 => data <= (x"0effb1358110c997", x"923c17d58e400539", x"40450f073930f3e0", x"d0731ef1139cd0e2", x"fdff2636d5cb1192", x"61da1036c9e4d6dd", x"3f0e235a398d535d", x"6181778010360627");
            when 11649432 => data <= (x"51b52519ae50daa6", x"00f79a5ed95094be", x"633994d4e683a011", x"14a1dc10a77c33d1", x"450c40137aec7df2", x"1ad863cc1028af2e", x"c36e459aa562a52c", x"8fb26eb43f445924");
            when 12369061 => data <= (x"c0d8e0331f317daf", x"ded4764051b3795e", x"fbeed15f7312989c", x"b00438ca7a02b4c6", x"5b1ddf747e55faa7", x"946ea8d9f9b148d3", x"bdff91352ec7559f", x"e4daa35426261d64");
            when 5804258 => data <= (x"7e79e6f26b4f25ef", x"fce39def7ebff7bf", x"c8af68fda53f966a", x"d48883cadb719857", x"721064a49958157a", x"40256c7e69e1dc42", x"2dd4fa81e16cae60", x"ce6740139242ccb7");
            when 6673080 => data <= (x"72f3e654bb492276", x"ec3d0e7765e71326", x"06e500dfb0b07708", x"eaa906d14a3a48f1", x"aae075682ec06e9e", x"a208bbc70a5f943e", x"d9f304876a92d743", x"09c6584573f0b525");
            when 11881935 => data <= (x"21a07d32e8193fe2", x"b2a3e775f6a33bb3", x"0559168c4e78d05a", x"82deb53ae67b733c", x"8f5b0ae345789d7a", x"84fb81a88af205e4", x"43f70d4dd07f8511", x"aad18fb120c9667b");
            when 22012570 => data <= (x"cf8f6bf9b3b87e80", x"49f0067c98e74598", x"72f453be4c377d18", x"60595e64c9c27d89", x"a35b602c6493fae6", x"934ab409c0490b88", x"e7f6ac7c280e33c2", x"84277c479a6961e0");
            when 30273480 => data <= (x"3bc42059bd984c46", x"11c889a66c7a2696", x"61593b8a65139ba7", x"f51702fe7f7473e9", x"3bcefcaf5a519fbc", x"1f2d468bb4e2cc81", x"e9de7ec3ad071742", x"1edf34db15e65d19");
            when 5395395 => data <= (x"354ea1b63c014542", x"cbe13da248fa35ca", x"9213c4a388f76bd2", x"49282ee4f3dae6b5", x"8e65daabc419af48", x"1673e7d8ef0e4490", x"ba47f91ad1e00e56", x"d560c52ae0c72db6");
            when 21861947 => data <= (x"afbb5e8208737fcf", x"c4dee2b1f35bf3d5", x"b0aed2767720c624", x"7fbf434c53f92e94", x"e58aac4ce9969d52", x"6152e9e380ea59bc", x"d753eb2782cca3b2", x"8a193425d19fb281");
            when 26914817 => data <= (x"32267ccfd045fdd5", x"0aa9efc3c5984a3f", x"e055fbb768a7673c", x"03cb3658675bfedc", x"16480f7ca9660a33", x"6affa40047a8a68a", x"355a8d0af722683d", x"e7b8cb6b0e290900");
            when 14314029 => data <= (x"e2bbf551016b1c4a", x"7316675e5282da01", x"825a40aeecc60081", x"1c72132681bbdfa6", x"9ce54b84a07e60b7", x"e4725701c267a721", x"57790d1f6640c673", x"8916a5ee46f6f6fa");
            when 13817512 => data <= (x"8c00c24cf61264e4", x"250c3f8ff45e91a9", x"cc80c4f662a7fb8a", x"4179a0049342edda", x"38a85f350ededdab", x"5f6e9dfc6f88b465", x"86dc560a5c49c0ae", x"0c19bc2a157197f1");
            when 27451656 => data <= (x"9cc540ce22da14ad", x"bde9180d95ddc6b0", x"9c5e75be053c0b94", x"fa5043eda339ea18", x"ecda906f68af4371", x"bf7c52dcbeced759", x"57569d5891495973", x"42071b333853ade8");
            when 6558256 => data <= (x"973a96a0a0a60875", x"2d9f400cfae49cab", x"0f7fcede68936ece", x"9db2845807f32441", x"4408f8b28d831947", x"34617965f7ec635c", x"940740f5b6b990a8", x"4597ab810928a01c");
            when 1855692 => data <= (x"cca8f9f7cb6bd98d", x"55d7ff18fb4c4643", x"75e3cca819768104", x"bc4101c662f27b98", x"258b82b8ce90cf50", x"ad490a987119d935", x"28c8ea6cca3e8ff8", x"64e28cb1d887f3b0");
            when 14638205 => data <= (x"fbdb9bb9d08ca60f", x"2e23a1b428aa906e", x"741bb6e51f1f71c1", x"b8b6a7d704f0dfdf", x"81c091f57a947d20", x"1f8320c86cd6324c", x"dc57b8ac447395e0", x"9ee5b14a225d0d12");
            when 9179039 => data <= (x"1824ccc8697761c5", x"ab5aa3d807e938ac", x"00906e2f384dd557", x"6cc302681c77413a", x"da87ae905d09367c", x"bf1bdb852d8963cb", x"c7bcb8a98e36c5e8", x"e238d79c49a6aae5");
            when 32059287 => data <= (x"ba7c4e681361142c", x"38630cc725c3bee4", x"8e3ce0eaf3314078", x"05d7b9370f814675", x"20568d6584361710", x"95df927c14d8b235", x"cd44a261f7e60eca", x"9c43878e5f7979f4");
            when 14885447 => data <= (x"58d52bfe967e70d0", x"1d524ca7c93bffe9", x"067478714435bea3", x"f5b6b2c2b72bfe6d", x"321c9397103fe3f1", x"29295a89cb12c4cc", x"c8ab6d66fa324eb0", x"ac640253997399f9");
            when 22407140 => data <= (x"b8623da8e070fd57", x"342de4ffdb2b6122", x"2ca380f112ed3408", x"9dffa719ef7ae2b0", x"36223c82eb829404", x"d78a6ad03a232819", x"869a4432585d8d09", x"868ea10d4a2997bd");
            when 29995206 => data <= (x"f1aac21ecb4ce35d", x"58554c87472e9d36", x"e905d54dd3743a84", x"0649574830e3fb86", x"04eb5126dc972694", x"4b77a6dde12810f5", x"cc820b5356603789", x"9d8ded96c7fbbdf9");
            when 25713504 => data <= (x"1b3bc003339f706d", x"18d149e21911329c", x"9b385d3c2ad32686", x"7122b160c33de741", x"10c97c8a2b62402a", x"ca4b119784bbc78c", x"6aaf70c0447da7e5", x"3691ac52b00120d1");
            when 22412462 => data <= (x"3698be8874245b37", x"84d8f53cc83890f8", x"c5b769bb2509cd64", x"ea5438b2c2d19e2f", x"4ebc57fd73457f93", x"fefd07fd8c791bcf", x"cc9f5ec61ed98c35", x"5d333d3079dbf3ce");
            when 30508948 => data <= (x"ff926bfd1babb242", x"4231e6dcd05a73b1", x"4e59c171829657e3", x"15c70fecdce4a959", x"339c0193b4187e85", x"4a661e541202d64e", x"7f471d2da8da5343", x"2f3d017c60a02ac9");
            when 17242049 => data <= (x"8d5fa0c5ccb500f7", x"41992cafa5d459ef", x"7099e32a3e1baa3c", x"f98b5c3654f82421", x"bfabd4b8f12151a1", x"1f7fbfe7afa23b50", x"81a68e9b12aedb07", x"8d3eca1a6d2137a6");
            when 22038914 => data <= (x"6ae821df48b4db94", x"8ace284c299b28bf", x"5ef5525ff7ed2a7e", x"60079b6703c86479", x"bc67353b1a18774a", x"2b621cdfbf66b216", x"7853170abda577f8", x"ec0690c6110e9a04");
            when 12508884 => data <= (x"7fd6202d9480cb28", x"9ebd781bd2dc3dd2", x"a30ce18a51d09680", x"1664ed926642d0cf", x"078059deef2a5802", x"b0149a51eb0d1b50", x"fb2ffd89fa2015c3", x"a403ff292593baba");
            when 4391134 => data <= (x"e18aa2fd5101edaa", x"e1e419174edd7073", x"7d36806c4d5e531e", x"d02eee29b20bd3f7", x"b293e507a6b1dc6f", x"dc306b683f4262ab", x"3b74e11b84ad8e86", x"7e8df949938e8820");
            when 7623143 => data <= (x"3925c059673356a2", x"df8b6dd5351a96c2", x"b600a59901b764ec", x"94c567032620998c", x"af9192cbe63098e8", x"120722795f666b8c", x"3a2ed9843cb50a1f", x"6d1479c33caed54b");
            when 27999044 => data <= (x"3ee053cb6d6a27e7", x"7de3cad3b6bc6b13", x"26d84c37b9ea77c6", x"23edf54038305bf0", x"70d95930abefd925", x"3f85dad6f547cbaa", x"f6112f8b71110d5f", x"6ed8fbadbfec9cc1");
            when 1171114 => data <= (x"eaa83a6296af63c9", x"2c8acfef6a3ecded", x"ab458434d812f3d0", x"e2cf1538950513a4", x"af2bb592472bc529", x"f6f5914cbd121e42", x"2e25fe828b5f3021", x"945bafe0fd7ea32f");
            when 21208133 => data <= (x"51668e9c2d8f18d2", x"41f08c16e5e390a6", x"ec11ed77d70a6042", x"173af1a3d3880158", x"dbccee5dee916c08", x"c2df8e0880807462", x"d49f4700e28a7081", x"0c8ee7d739e97fb4");
            when 13856901 => data <= (x"16ed84773ab9b2d9", x"94a947d77c51d8e5", x"9511dd639b723f3d", x"fc344aca24305af9", x"19b50995698549e2", x"8ae933020972c262", x"d4d85d8425d6b225", x"3b37d4c880f21a99");
            when 20213001 => data <= (x"64f392aede6e1bfd", x"d29a781329537d91", x"7964d5c13ae75235", x"f947d8b146e58eda", x"7f5da6ed2e48af7b", x"eb4c12d17489d0d6", x"aed5231982e33479", x"a55c03618eb107b5");
            when 32824624 => data <= (x"132bd64cba8854f9", x"469a3c78a586e9fc", x"1beeaac70d9eb2d6", x"977a61f54473895d", x"18c6f5c8aec74c86", x"68eeea930e57b6fa", x"9942f2cb1a2a40db", x"01e5cf4e3782b394");
            when 10070155 => data <= (x"7de81a298ef9ee86", x"064dcbcb64f5129c", x"b986cc0c4dd6e7f5", x"d1e18a9c7af12d26", x"41d8b9c9e8a4a9b2", x"7ba0989caa34bcf1", x"e6e4004ebfd3609f", x"3ab973b451559e95");
            when 13689597 => data <= (x"3b93c64039599fc7", x"691d8d08b2735a60", x"88ef11a5f1459426", x"d31c0d5253490402", x"60cbcda9215746d8", x"f5d231c55cda163d", x"56844733dca54187", x"32e3fb81b8503e57");
            when 32035279 => data <= (x"16975ca97c1a5a2d", x"72fe248e263e7ed6", x"af148582a9e6ccdf", x"35d9d7785e2fda77", x"1d563008a657650f", x"19fb0251e7e44949", x"a41f074589d45394", x"86cf385583fc97c8");
            when 10134947 => data <= (x"3ccd3d8a3b561e5f", x"938d8e090f581b39", x"878ec43a5d4b219b", x"67a2b92c4588a3d8", x"5519ef73b90fbd91", x"e84ae886f2742c0e", x"a2ca847c8bcb785b", x"70e4c65c5c9ac7a2");
            when 18110056 => data <= (x"fe5f348aee4b8766", x"cccbb1f8aa7a0462", x"2c7730502bd98b26", x"40bb3795d949ff3a", x"46bdb1ec55f4191d", x"f687b10af5dc944c", x"c3bb3e9271f79134", x"d8dc097ec060c1a1");
            when 13823649 => data <= (x"55357fa1ba2c34cb", x"eb0b9d5653447ab0", x"0dbea1497266a54e", x"f2a29263682264b1", x"3d643da7dcacfe08", x"e5009d8e5cf1a562", x"5330bd15d49405a2", x"9ac83b70576dc6ec");
            when 5107013 => data <= (x"800b6709383e69e2", x"4cb123a97398aa23", x"7bccf4d592b5b94a", x"b021c5626529d172", x"3179ebd1b4cd2328", x"70871e73ff2526ad", x"fd51026dd85063d7", x"979f818b11732e2c");
            when 21034529 => data <= (x"58c5a2f533f9854e", x"a7c5730ec6e66ce4", x"0ee2dc14afc80f89", x"31eafca747b5d597", x"2a934f2eb132b211", x"ab05985f359a2780", x"df7a89fb8ba3ce4d", x"badacca938cca07b");
            when 28107096 => data <= (x"27bbcb10bc55166e", x"3b49856e824f624c", x"8bca36b887b15a7a", x"84e9a728b8cb9532", x"d0936f9bdb76f1e9", x"842faa8b64a8a0e6", x"21f12cdc0874a5d4", x"09f7a436bf6d60d3");
            when 15471800 => data <= (x"9a5a6e5b57375f3f", x"5dbbe38a6501ce12", x"d9ef3229a1a853dc", x"724f2f44bde69579", x"97b37bca88e814cf", x"9288362b5e64efc4", x"12e426dc88b8f234", x"cbbe3e46ef1777c9");
            when 25321852 => data <= (x"353f4e023313fa5c", x"3456e8fe24cd68cf", x"4e84a367e52c344a", x"a9051db8faa0094f", x"31c4ce5cc94df401", x"dd22b335df25ef53", x"a8cac7583e611aec", x"9ab947092519d79a");
            when 18312720 => data <= (x"3e8f2349de1bf985", x"d5d74dd7c5ee6894", x"e35d588711573c27", x"dcab555c81ea1680", x"625e5c28471f542d", x"758e3d51f597a406", x"65c7f0df3c5b7264", x"07f004597b73f7b6");
            when 7469019 => data <= (x"b553730206ae096b", x"49dcc197caf06c90", x"8a03d90b58e09958", x"93b70c95d30a7ce2", x"9d654136cd01ff55", x"d1910d491177d950", x"cfd17c2cf55e3116", x"d3b50d329d741cb7");
            when 21781041 => data <= (x"95d5e977b1d747f1", x"6040e05cb2700e9f", x"2a342c143b582e20", x"a9c69d2a6451443d", x"577eea5672eb706f", x"03abd76a121c2f1e", x"6e303fa445585e16", x"92a5800d3b1404bd");
            when 2420431 => data <= (x"3db2e16614c55e07", x"b4b3cc1763118787", x"6bb29df9d89170fa", x"cc10649630ca1d48", x"5e2543309b3ccf43", x"2e30c010728e26ce", x"250c3a90d9757e3c", x"a122d6a1de8dc948");
            when 12721101 => data <= (x"67726931b6946976", x"cc9475eb6d5168c5", x"3b672c620ea16f3f", x"39e9e998131c66fb", x"64c0926d1f07ef28", x"74a00a6ad854ff7d", x"4df9482be99cbe58", x"2b5c50bab947acb9");
            when 31411959 => data <= (x"c62ad6a0a34ff1a6", x"ca6fa3b62ba897e8", x"320887bab42260b0", x"f671f767ee583741", x"987f120fb1766b63", x"ad9371709189a37b", x"832ae71b009953e3", x"f86bb0ccfbdc35ba");
            when 15004764 => data <= (x"51145f49616f457b", x"3e3dac8b301efb3a", x"7c75e2117ee90059", x"221a7d9a1690f5a6", x"d211d334c3d7c338", x"1533c59c7765206a", x"dfbb545e2ee55965", x"dc6a44755527bdf6");
            when 20305029 => data <= (x"9e7353bd585a8507", x"633b58c17d758394", x"c7eccc788351d6f6", x"79ff4ae72264589c", x"ad1bf694b2c48387", x"a149bd71f484b538", x"3dced40b6677c40a", x"8bc35eb2b4872213");
            when 810259 => data <= (x"0e6f51b918ea130f", x"ebf29e4e71b6b835", x"4f7862618f610f06", x"0985408dae3132f1", x"23368bd1919f2d16", x"f2b366028c55a5af", x"55989de0d417fb0e", x"cda5837b7971a73d");
            when 25420851 => data <= (x"c31977483d531e03", x"79602d95ebc55687", x"365acb5eaeba12c8", x"a2c645a8f680cbd7", x"adc65ec223f1b7c9", x"9acbcb7d6e38b77f", x"c771815428cc5e89", x"084a87e1a995fcad");
            when 11063825 => data <= (x"bdd7ce760828df24", x"59d05a565c463c5e", x"3f987b8235a412d5", x"24b1e35ed3eac7c7", x"360a7a419ebdcad6", x"4b9beb815dac03fb", x"fd9c789e51ef9f55", x"b34ee161b45db611");
            when 11527994 => data <= (x"3d0e3b6e0d889036", x"dcca331eee653aa1", x"e24d014a27ff3d11", x"230b58d348d41fa0", x"fea45091da83923d", x"495494a5b676c911", x"649d30c6d9ef0037", x"c231c1b106a71e84");
            when 14358860 => data <= (x"0f8b7e90f780930b", x"5884d99e8cdb9b85", x"a339d9e5ba9a36e4", x"cae205f0d84bde19", x"a786ccb211ff9f17", x"de2109ffcef56cb5", x"aca1908206b975f3", x"855a69f3dc62fe1b");
            when 30614203 => data <= (x"e06acc15070c20cc", x"f011d4bf5c76a0fd", x"1f03c1fede19db1f", x"d46a86b4cda9f6fb", x"4a3259861d91897d", x"3ca2da3bdab1a952", x"7b25488859f1e627", x"8d1df90079830640");
            when 29134850 => data <= (x"92aa6a4a10687323", x"f75feecc87432370", x"0d37dad3e9eabf88", x"18fab69a3e089f72", x"fc200d67658608bb", x"9dd394c687a1b887", x"cffe638114a749be", x"a9cd7f4ccdbd159a");
            when 31279455 => data <= (x"fbeb21d84d004f82", x"2f33eab74caa0ed0", x"320957447aab0850", x"279fb5f9d2900725", x"1a4ba45c00a21f37", x"dd8b20581ae7426c", x"66d769ccd8f836b4", x"0e89928dc36b0e3b");
            when 27222820 => data <= (x"625c1f0d4137999e", x"39ba49b7de72be38", x"8a1f99551bd3d97d", x"40b6c905eed88f78", x"dfed5a2b1be31d8c", x"870502f11e40fec3", x"fa1d429ebd37b682", x"40d4d905565c2769");
            when 5569950 => data <= (x"763aeee310949461", x"68fe31b28bf71628", x"7fe4aea02f08c589", x"3bfc4b28a72bb4ff", x"4d67c4754bc5d518", x"6ad21ba4515dce9a", x"d91115a095b0428f", x"81d7743865107106");
            when 7988847 => data <= (x"3c71174da075f76f", x"695acc606a7f2578", x"6ee68504df46a091", x"4baa39e8a7aaaece", x"9057f84ec26faeba", x"e53c968ef0a2f58b", x"d6aeaba26f3069d6", x"56bea686a7d619e2");
            when 7406773 => data <= (x"0d2ed02c8a1b4ea0", x"633b8c44ef8a3d35", x"dd261902129697f0", x"9a7785b45c5640ad", x"0cab60c7d8f819ac", x"e4146758a9d6b7b1", x"4675286c72ce942d", x"08ec3845e5c14958");
            when 16043218 => data <= (x"19c38e763be01e14", x"cedae9b603bf18e1", x"4ab5522d5c9a512e", x"8380d41055c59a47", x"925cc96320da5ec6", x"9e88deb97cec78f4", x"b0ac8d74bb4f8ff8", x"5c59c2bbddf40ef9");
            when 14617654 => data <= (x"ce5782db65996c2e", x"5addc65cf96e3e2a", x"97fc3f1db742d357", x"0fa58a2f9d692d39", x"a079f91c40c5674a", x"0c20aa38c6320cc0", x"3e9829623d938280", x"21d2efbc8ded10a5");
            when 5324826 => data <= (x"8bc7307b4327ca6f", x"d3fea78444ca1569", x"833599e41fb4ba11", x"5075a137f477c15b", x"b3310bb2e3a00de4", x"a0c68fab7bb35043", x"050d9c65c02ca9c3", x"ce19caa2930eb3f4");
            when 28514952 => data <= (x"ea45359b2d4be33a", x"4a887dcffe3fd462", x"1bf457c4fc093696", x"6f415f6ddb182199", x"6d5d1a657d86b622", x"1598a03c3c43779e", x"3117bfff4e95db7d", x"9d1eb75e420af54b");
            when 28063718 => data <= (x"8c4bdd73bf6d0d77", x"c4f6189b1e14a33f", x"b3408b6ea7b55cbc", x"4e24aea3270ae93c", x"83c00b2f90f9b569", x"f286f3fc2f2dbf00", x"8dd09a80e05b6f12", x"241e884eca5bc9f1");
            when 28025244 => data <= (x"38d226928f1ca899", x"72a6156c0cf7dbeb", x"017cb32605b544e6", x"50ea95e8526f6eba", x"a9ac2d96f099f687", x"a72ea4ada3ca2839", x"355f1e7bf89119d3", x"5f2f53562337950d");
            when 8640136 => data <= (x"3a50507d28f5cbcf", x"069af72a229e37a5", x"96bae45ce407fca8", x"01b5cad81917d904", x"e23d1a4f43f08621", x"778a6b13b752e536", x"875b8a976e9b79df", x"c0b63c3199708416");
            when 16191448 => data <= (x"3f1b82e30e226654", x"d535b7bf09d4c82e", x"121a3afb51261c8a", x"be1734fbefb0d789", x"5704fd04f99637d9", x"ead26334b28c6ae0", x"8749475b031f6470", x"776507100c59b5a6");
            when 18998426 => data <= (x"a5cdce2d698d9518", x"e2c31e32a1d3790a", x"b1aa17b2c26c44d0", x"e43efdf6d6ffccde", x"fbf292fc129fcd87", x"bb0536dd0b978c85", x"25cd5eec12ecc894", x"6d66b8bd8be1a043");
            when 26605580 => data <= (x"4e8b8c99b3c1821c", x"667a10255a255c7a", x"9147db81e060eb14", x"9450b744d88bc170", x"2a7c165228a4e265", x"250a368d84fbc366", x"51fe6ee72d5f2534", x"47de2aa2da411619");
            when 16298633 => data <= (x"f31f046d069fe3dc", x"7fcbf91db7f0a6a1", x"205e6428a898dc38", x"23c289df2f10e739", x"43dbb786f5577277", x"ccc123df2eea82e6", x"514f7c52d336e482", x"3c962fc6f55d9e28");
            when 14802579 => data <= (x"245435825d688c58", x"0f2329844f332b79", x"79b29363e6437a47", x"f4f6b7bf147d21f9", x"4208f19b1a25b4ce", x"07ab1d816d02c7d6", x"4324d41b56218934", x"a698c41a8c3c9f1f");
            when 19423376 => data <= (x"bd65c81d5d6e5c0f", x"683a2dd8bfc17323", x"864f5cbe5e6777c6", x"cb2074c905f470ef", x"2f7977ac83f4d590", x"133100717cabb701", x"6ea6cba997a6e4fa", x"4cd859416500c04a");
            when 12719565 => data <= (x"abf34dacd8fec2ac", x"5d42d62819124a3c", x"49d13942af9aa614", x"04e8e5a388629c3f", x"a940cb072b8e7748", x"7614182eecb7331a", x"b78a3f112661c00e", x"2f905ee45a9a684b");
            when 29862595 => data <= (x"a730e11835607f61", x"34eae31a7a85968f", x"fbe2c7a9513aff0a", x"c78f47891f874455", x"21bd41428d93602f", x"b7c76b67c81ca3b9", x"7e2e720e6eb6c0f6", x"b4b736f2fd4c3bae");
            when 11635949 => data <= (x"04274898478a9262", x"ba62274ee8fd1ac3", x"8cceb398c3297d0d", x"89ac60ea1a4e72df", x"69cb0cbe443e3418", x"30c489da30979355", x"d9e88c93521f2fae", x"390f22be4f34c591");
            when 29047857 => data <= (x"c27eeacc9196c990", x"947946a70ab47870", x"8cb6a7df5b48c7fb", x"15eaed03d746b0e1", x"88f2cb6add28d9bb", x"080654e60ee64bc1", x"abecde2c83bb1186", x"53f41f45fabcb1b4");
            when 776909 => data <= (x"11167d7c868137ae", x"742dffc65f6f1fe2", x"dc08cf03b306d2b8", x"f45f6e1cd69da349", x"87dc9521273e7301", x"d1bdc15b637ee249", x"40bc12ef0e48f9e9", x"ac75741a802f33a7");
            when 16171831 => data <= (x"70bc40a75741286d", x"9040d0ea8aced0ad", x"8dc84950e4a840d8", x"7c2411ea979a4722", x"47cd7fad3fe43e12", x"08a45722802b67e6", x"b2510d0a143a950a", x"08f6833cfef59e27");
            when 25001935 => data <= (x"7d6c64fbc9bf36a5", x"e696f8ee37bb8699", x"1ba5abca7e4283b4", x"ca93d3df63fa4897", x"10a54b6998339e99", x"f4103ef86ba7ec13", x"348c101d630975a3", x"8b3514470f286068");
            when 16046148 => data <= (x"7c40fd4116e74f45", x"50617e522c32393a", x"71c2772205f2602a", x"bf8477c5c3e5a51f", x"edacefd82b976b77", x"2d6aaaeea9345b85", x"7d71e07d47060bb4", x"074f6cfc36f4ddb6");
            when 2989363 => data <= (x"cf2780d8819c40e8", x"9e8ba70cbd6c1825", x"cc488ddabdcecdea", x"27d1d5a857263230", x"b3af646b9695c92f", x"0f4088f03c349782", x"cda01a14846dc0cc", x"99ca42d0c8735adf");
            when 20032226 => data <= (x"ff8ee35fc50d6760", x"eac64f702f08f5d7", x"3fe96e60f45aa4fe", x"25010fe6a4a9a12f", x"1ac151381a06351d", x"64b86b34ce730494", x"d03302dd7ce3c130", x"fd457b4236df35e3");
            when 27126872 => data <= (x"f4d4e9d65d42792a", x"fa39615375114544", x"656c2d736a662f23", x"8705e9b920eeee5c", x"41f548eabcd9cb6a", x"3b7f8bca2a169609", x"01de4329c6b1d6c2", x"e32981612ed7ff8c");
            when 24044324 => data <= (x"4d6e585ccc2de73d", x"a6799e7c8cae84aa", x"d07ee3898f7cba8e", x"7a2849741b6b2e85", x"3278fa28a446709e", x"bfc1d7a27680a8ad", x"94292956ecd4167c", x"aec2a266de4deff0");
            when 26074205 => data <= (x"f87af049f897807f", x"837c1ff49a8f9920", x"8727309c6048d853", x"b390eb85b857bf50", x"cd732729609d35c5", x"22e6506bb2507569", x"19e7d919436f4933", x"6eeac2bdfad8362a");
            when 13760096 => data <= (x"eac103542c785159", x"d4122291a755e4e7", x"e859f5c3cc51d90a", x"5dd4fd7aeb7ac793", x"a09e9fe23eb5a9d1", x"9b59a243001cb7be", x"f335654c999b9e5b", x"5ec2e30d19a5880c");
            when 18806813 => data <= (x"60f3dcc8969785ea", x"b74ec8b28ba9416f", x"2527075df1f5b07f", x"cce51881b99b848e", x"f5700f07c08030b6", x"05b3cf9a29134846", x"0b90627ef64cbf7b", x"b261c37ba4419b4a");
            when 23730755 => data <= (x"c5210c65beae4d8c", x"750f9cbc66a007c9", x"ea8a16f2f5031789", x"793d80e613b7e86a", x"3c3ea8522d88cc58", x"93862c04d516832f", x"89c2edfee1ec4546", x"90d933a7b757c858");
            when 31493895 => data <= (x"75e831a63405e9e4", x"6e3d10c3080baeb0", x"3455bba9477aa887", x"52167333e27c51a0", x"ab2c65dd73e61460", x"bcace0c86fb06382", x"3fed4fc75aa27b6e", x"8a55b7bdbeb82a10");
            when 2348683 => data <= (x"45d30bbc935fe1de", x"975008534d930ef0", x"96d3e1957f8a3c9b", x"7bb63de5428c3406", x"47deff14c2c69ef2", x"2c0f856e5ea28716", x"4575015ec5526b8d", x"00e9de71a9772e17");
            when 3344913 => data <= (x"e472348178a0aa0d", x"d276f3a89efef64f", x"208832f3ee523e05", x"cf7800a5d0d0d163", x"b48ca885dd7fa04c", x"e34c07570b8f5f36", x"37336e8aef7ade8a", x"7ce4dd43346b90cb");
            when 7564731 => data <= (x"e1dce874ab4ffa9b", x"7cfddbb1a9c55d0c", x"fa0c4701a4cd41ca", x"dc19571ab4b3bd00", x"ef5f3ce095b5badb", x"faa9c8f657fdb214", x"7310f691ffb10d50", x"09f4dc74638e1b37");
            when 7219553 => data <= (x"0961a892b68e8f93", x"a63a9752e3dee9e6", x"a40047374dc15b3e", x"a9adb9193fcfbbf1", x"d2545dbee754b295", x"3d1696a2573c9cd2", x"79edfda8e5e8d6ce", x"33d81579cb013b37");
            when 6288865 => data <= (x"8a693d281233d0ea", x"4e2e3c81bb5900e6", x"27e6bf603330d8a5", x"9f7934f27eb002e5", x"8b8e3718e11c09fd", x"3cdc0ab1e2ac38a9", x"a766e87980b1c430", x"4fe7beaa7154dc6e");
            when 23230612 => data <= (x"9d257e9634aeb4cf", x"9952afa08c0ec111", x"2a0d05fe6a7ecdf6", x"96017266db31cb7f", x"c020aa09131fe652", x"daa684f6f95cb8ad", x"0bd75c9bf572cc51", x"fafb7dc31b8ff74a");
            when 3173253 => data <= (x"b03f1cf6dc718afa", x"a546f79225190fa0", x"9200bcf77bfb9262", x"12bfdff16a5bd26c", x"8f4ce6a20769a672", x"1443052d6c8307bb", x"b4c03bb86b7f3ae0", x"351bc159fdc0011e");
            when 2791347 => data <= (x"cc703fbf922af722", x"9fc0223a4815a357", x"6856aa60656ffefe", x"f28eb78fd98e05db", x"2b1fd8a39e5498dd", x"1152291472a23a1c", x"4d099e8e22633c8b", x"02b813eac61a6ec6");
            when 26338052 => data <= (x"3cfa341eb184e603", x"8bf3196d5b119057", x"7a27c511047d342e", x"8dffdeba7f60d2a0", x"cadcd015aeb1d3c2", x"9a67d8148c79484c", x"2690869414f96f13", x"4c67c9d9f8bf05d2");
            when 32198390 => data <= (x"f042d5ed2ceadccc", x"ac7e69b4c3a6f3ef", x"7c40e3fbf96ca332", x"0adf7d183aaf4a94", x"21a4e44755236383", x"a4d53bedc598cea4", x"843fa567c6e530eb", x"73835f14008c1f27");
            when 8135672 => data <= (x"b5d0c04e264efe64", x"67ce5de504752abd", x"c02d7fea3c9431bc", x"d722b22bc7a2e084", x"ce12515dd6902486", x"9846b2de3f7cce53", x"6a92d9d05b1be24d", x"a106b36549b6cfd5");
            when 3271612 => data <= (x"1d808dad42442468", x"5427ef936d66178c", x"d27ec3930510970c", x"a9b21e55af12dce1", x"1fb3b1d680ba3f3f", x"79d0ca5cd45668ea", x"272709e13b84ec6c", x"cc9bb7bce18ccc08");
            when 21314914 => data <= (x"dbd3b9196617c6f8", x"06fbd8a7563cf6e2", x"d692808744a66ffc", x"7a2c3eeabacb0a18", x"f60aa78b330357d8", x"88dfbe476b1736e2", x"513dbe936ae6cb97", x"e0674fce2428d019");
            when 3859464 => data <= (x"403f8aacfb86c808", x"078f7446d6d55538", x"f03f3e0eaa16c98e", x"412fdf0dabc36bdf", x"ce731edf2709ed97", x"b824acc671fcf0dd", x"12b56ba7ef97022f", x"b8f90a48989a5e8a");
            when 19766264 => data <= (x"682651c85547df4f", x"6a25a3524c45f633", x"7914391c2533ebea", x"e64f0d658fc3306c", x"ffb43025b5a3637e", x"c82c312737140a30", x"c0837b14abbd53f6", x"8b39acb9d5eccebf");
            when 8588798 => data <= (x"6e6ea755dec98381", x"d50994cb4b3128c7", x"4c539310f19200ee", x"c6148e9294daecb6", x"125d0723ed96af14", x"22b9e5ec4b765df9", x"973b418aeab98463", x"8746a14acf973a25");
            when 19733623 => data <= (x"8df895391c00a53e", x"eb37e651a624e1e9", x"79b036b2e3ffefed", x"cd04042f397873f4", x"69dfee2252ae666e", x"2552329473e63f6c", x"ff3481a864f0092f", x"8eccd004b1cdadd6");
            when 26016827 => data <= (x"34281d067fcdb8c1", x"fb161624168ac5f4", x"9a0e22a1d58b103f", x"32d5d2070cc34f1e", x"4c732c37202f6e08", x"3c364a952be0c804", x"f723f14ebd427923", x"73fb9e2fa6b27b67");
            when 21964569 => data <= (x"f823bb1374d8a822", x"1c31c310ecbf9bee", x"b2c19562c0a1366f", x"aaa3c5fd69978a89", x"c0cee09c9806cb8f", x"f41f2aca58a363a1", x"ff43da19920ccb03", x"d8ce70d9f4994723");
            when 16673818 => data <= (x"ed8172c6ae957bc0", x"67148e0dd2872c1c", x"19b6e761e0fb2ab4", x"fe3470f786959d17", x"d71d90c482d8940a", x"ee41a5f01ae43f67", x"ca860a347fae6ced", x"dbe00ddfa3640d6f");
            when 33780928 => data <= (x"58252bff926e58df", x"c867f38fec63dad5", x"561ee2b243ec9af1", x"3bde450449b481ca", x"476130a5c38621a1", x"08482e7667fd0aa9", x"920d74ffc4c1d75f", x"571cf3bca998ef10");
            when 26445066 => data <= (x"de3a0d65570cdb72", x"919f23d2d9042197", x"b6bf2737b3c76ef3", x"4acbaeeb6ad9829c", x"0049f54e03924cb3", x"d3111e6d1c1ba4f0", x"ef3255b842d856d3", x"861468df331b9dbb");
            when 18822779 => data <= (x"28778038b5a150f8", x"10a8eaacd455188f", x"520a91319cad6287", x"41aa98008c3d5dbb", x"a17ac2203d557aa6", x"2435b2d8035e7c0c", x"738bcb017190d4d1", x"770806c2a24c3454");
            when 10813526 => data <= (x"070f7520c99b0b80", x"81dca6368fd48c2a", x"2d8a09ab83babf22", x"d019e24bce8f30ae", x"3c966f1a87cbb901", x"dd2ac17edda4df15", x"f4dcb938bdce8f63", x"e6603c3899b8f121");
            when 24777647 => data <= (x"7f1ebc5955d79d81", x"7bd72ae2e9f295ce", x"d5be5e2fd637f8cd", x"084133e5ac6127a7", x"5523e035467fc3c0", x"918a98ddc9fac12c", x"d9d3b419a7c2e88d", x"027fd7dbc0d5d82c");
            when 4600014 => data <= (x"c5d5998c5a809719", x"38f26b0ede033bd7", x"7f51fe92c87a87de", x"644a93f884c2446e", x"c544880f180f4450", x"8db5a3dfcfb9b751", x"3f52fa6e50efbc63", x"65eb153b39df9c27");
            when 28163017 => data <= (x"4bf35236a350145e", x"590141d0d4a93576", x"becccfcaeca0594a", x"5e196746d81434cf", x"6294da37cec5219d", x"bf4d9e4b72e0f303", x"dd072d439dff6c45", x"a4010058d51cc688");
            when 4916410 => data <= (x"a7f293670b090a8d", x"5df64c64eb2d4ff9", x"00c13db804140a3c", x"57a84f9567c4a4a4", x"e89306c356d0e261", x"f5c49e5c8ece55cd", x"131bb91037b60a2b", x"43ec9ea71a106c17");
            when 17787888 => data <= (x"a5cea6df86e1bc99", x"954226093e52e88e", x"b5e5b8e63f92bebf", x"ec26548ffbe99151", x"b4a5a5a356a7d64b", x"067e089903a566f3", x"3ff676fbb32868a8", x"5f3a97495b0bd99f");
            when 8556039 => data <= (x"e8d9cb3a35b8d6ca", x"609830b6e93beb4e", x"f31db3a7cb5db07f", x"25f28e0ea847325f", x"68d5146972d515cb", x"d96fc0647c543863", x"5f3d466e738e00e5", x"024bf4b9da2454b2");
            when 3596664 => data <= (x"a9f740d3392dcc45", x"3422e40ff8205444", x"3d11b996ff9647c8", x"28ed1169dea59e3a", x"a0ad86b4b11f7600", x"62df36a32360f18b", x"b9b1df9e57f3796a", x"9b54f80368b2d862");
            when 9499595 => data <= (x"658f3c1cee7c78c8", x"175c1225d781ed24", x"cffbc3e881df2553", x"89ddceaac2b3f891", x"041dc3236385f3dc", x"d80c356c2ae5c2b2", x"4aa1c67ca8ffba52", x"15fa46ad9f1d745a");
            when 9762497 => data <= (x"c7677b457db5412c", x"15d6751f7060f3fc", x"cb1503947aede3ad", x"7bded3f4ebbad759", x"d15108531442a14a", x"e55800ed9ed279f6", x"d967e829eae6e66f", x"dc3424db3c8e5293");
            when 11327001 => data <= (x"c5593868266ca791", x"3cc13a044d904eb0", x"7d784875c56aeced", x"31c930fbe8d81e19", x"ef73ddb4f5857610", x"66a181c84ee7042b", x"da3b3513e10d98ae", x"bb07faefba7fa440");
            when 31718298 => data <= (x"e2308b8dee4e2d9d", x"ac89bb71f9f0658e", x"05ceb100f13bc395", x"1d9d5d0ff73bccf7", x"0c79ba36bc4549a6", x"e4b04b4dcd7dc4ac", x"480d176b420206e3", x"60cca1a67008c78c");
            when 30960145 => data <= (x"ff8d3cf67b624621", x"b14446467f541982", x"c629c0fa55abe2fa", x"c6024a49af84ddb7", x"dcbcdd44263c6036", x"c5e3aa1e68261de8", x"4a1d2102b5f4d668", x"6a98d103fda3c4ed");
            when 1428539 => data <= (x"3dd2e18e994d685b", x"371984adc25c5e06", x"2bd47763059c5bd9", x"89613d629f17a7d6", x"c648e223af9c511c", x"0bfeef77d19a6c09", x"b065f33e0421cc2c", x"871ac230f6d8c513");
            when 19107239 => data <= (x"fc1064dab5bfbe37", x"951b1e48338cba31", x"0561013006d78bf6", x"1ca180c7daaa381e", x"508a6ae991e1451a", x"3a88f74ac9d48d31", x"0f6286a4fe01e1e7", x"406c8545035de0be");
            when 31336584 => data <= (x"ac677bed4a790fd2", x"f41a494092ccc1f1", x"a9e551e5ede2df45", x"95ede48a69fd55b0", x"b4043e917e159ce1", x"9168d6975b65104e", x"4c61b6775737400b", x"2856277b93239ad8");
            when 23054010 => data <= (x"a23f1a4e332728be", x"03edc98f54792d47", x"871c42fdc9ede0b1", x"2846c93ac29d53a4", x"c5032a1782950fb8", x"f8c27ec0e301bc97", x"631ee9d9c6c66a0e", x"cfca0cd8c8e8795f");
            when 32390294 => data <= (x"c30179020c48e6c9", x"6e52f2ec19441531", x"fd7164adc21e2617", x"265970afb0ce04f3", x"bad9d74ada1c51d4", x"ed373cbac124898e", x"e1108af535df330a", x"f1ff6537170c7c59");
            when 25592767 => data <= (x"64fbecc214284f5f", x"be65ec1941bdef81", x"5a7e2563906752f1", x"275bc547333f7658", x"292cba6ea0267249", x"c2f43ba76f7e37d8", x"99d9ce0a28eb98d9", x"bb0141fd14e0c9e4");
            when 17585003 => data <= (x"2a42a34de22fd04f", x"6cba086128d4f6c5", x"932878c0499725f8", x"5af132fe957c6699", x"ab5ae6543ca2f5a8", x"73250c4cb34dee44", x"001f9c1d4bcd3a0f", x"101a0b330267584a");
            when 26398676 => data <= (x"afdc4ab97fb14c95", x"8204bb6214c07374", x"6c1bb07585f50195", x"d2073650f459a4a4", x"22ec0d297f1b6c5d", x"afb5153a796f2769", x"1e96a390f95b5e42", x"63db1ee907e3aebf");
            when 584787 => data <= (x"9eb9a0d2fba78fc8", x"e6604effba3f1e27", x"2a5e3284433ac88d", x"d23002430d3b6ff4", x"92dd3b1ad6004dd5", x"590319b2c80a7f70", x"6eb1c8fd78541cf3", x"755ecaf1b3daf2a7");
            when 30308252 => data <= (x"0f4ea984a5534903", x"401c3419d229b7f2", x"fbe56c12cec127e5", x"051f8a4f0b08e4ed", x"7be667e6212130c1", x"6392150f4abd26f8", x"e5b5a48e66fcc9a4", x"b34099dedbef2c0a");
            when 10854632 => data <= (x"189b7c9560ce9db1", x"8fb920a37270d2d5", x"d0a0481a8362ed24", x"28a35699d7741bbf", x"3027bb9840538e8f", x"4a316c1fd5c62a6a", x"b0be1eef1c6c41e8", x"4640cdcbf36c8def");
            when 10549619 => data <= (x"7f2a3f5eb0bab14c", x"64215b5658d3c23c", x"d6749b6d484eba5e", x"634db8e019af7b00", x"70cd2ad9945096fa", x"9a524a0f5c1a99ad", x"d577464e66099633", x"3cfda326261d5a6e");
            when 18143173 => data <= (x"a2b8e4d97bdb7a6d", x"ceee3c0ded9814f7", x"504476270de39101", x"7c7db90f13e1b410", x"f0f1f7ba8da2037f", x"ebfc36adcf8b8c31", x"ccb485b7eb99e5ac", x"484261573ef70548");
            when 32676460 => data <= (x"41c95b847e15ce85", x"3b0632f588791142", x"b66af7d002b48d41", x"b853921d7ec2989c", x"ef9c369cd1788410", x"7984c55f8f2c5249", x"60cdedd8aa192578", x"b9dcad70f8d835c7");
            when 24750188 => data <= (x"0924bd5555549227", x"61bd8ca1a94009f6", x"3c2066eab71daf9a", x"9fb999b74042c79e", x"95e6cd6fc67485ff", x"625ebf2899903644", x"8bd091a3124eb546", x"eadd12ec8b64a3ff");
            when 23143531 => data <= (x"5bffc5d2dca7930f", x"d89c2a9acd683439", x"a336621ca6add970", x"f84baa94f8dc868e", x"a600a345d3a5a92a", x"11c0c1c02d88fd0a", x"d574f081251b9b9a", x"a70a9f781efde9ab");
            when 2555966 => data <= (x"1b62bb8b44a934cb", x"a77c5c258748e1e3", x"bc922ca8bb9b0a6b", x"ab2f1b6576196235", x"11c01f37484333ea", x"10cf9ec78882a299", x"c6a50bbbd552dcba", x"be4f6ce02c2f67ce");
            when 23803844 => data <= (x"fb8af9738df7dfd2", x"53e016d0a1131d2c", x"db1536f585bd79ea", x"2131b47f3a57b8b4", x"e29ebd543e9fec2d", x"63cc2689b91f8d62", x"87b6ea5e1df50c6e", x"cd4583ed489d65d6");
            when 4312807 => data <= (x"d6a26c4c16f20825", x"3e32b16b1188721b", x"0bae142ba2c09fc1", x"d898c94822df17f8", x"0bff1bc16c7695a3", x"77fc219defd8c824", x"77d31740da01f4d9", x"a1ab992a6007c2f0");
            when 12857460 => data <= (x"83e9e7d3bc81cdbe", x"2529234343e91e5a", x"da0af7691a552fda", x"8b472d23331c5615", x"b8fe86d1b74d3879", x"528904e1f699fc4b", x"39906a8a52cffc2a", x"9f4842685307fde2");
            when 16174653 => data <= (x"133e194508817909", x"95cd69f6b5c36ab9", x"9cf1307aa088af0c", x"f747db029bda44a1", x"d0c4680aaa9b53e5", x"3f9a93430be3cd88", x"3853be1d3080cbcc", x"51f56204c59e8c67");
            when 10428304 => data <= (x"2f501b33badaa76e", x"bd59133d648d38c3", x"b4dba7fbbf12b456", x"47d87d1bc942fd2f", x"63caaff59619a0d5", x"3f75454d1a980fcf", x"db49c5d8ee41009e", x"2491f8a558399a5c");
            when 25741852 => data <= (x"bfcd002159029795", x"517dcd9a68b0c8db", x"991af1ba9080fe0f", x"5bf25fd268eff692", x"004437b7e7533a2d", x"a1c0772b8f1b77ea", x"e5a501a2a4201fd1", x"21e07e515b2a24c1");
            when 4511073 => data <= (x"b1cf1c1842ad8c27", x"1d78f0b4016c8333", x"5636c319f490361b", x"02e9efdde4ae10ab", x"e0d7e0f32311a7a2", x"0aa2d3dfae584741", x"89b07214d1857518", x"1d0de38ffcce178f");
            when 15550551 => data <= (x"1b93ceb78819ba36", x"deecbed5db979566", x"f9c0db03ab93c21e", x"649500fccb6169c4", x"aab9865454622a42", x"206d81ad90cdcba8", x"2ebbc46c3642c955", x"cce2964b40b6f673");
            when 12688886 => data <= (x"a6991c6cf627bd2e", x"09dcfcb60e2a488d", x"850bfacb6db39d05", x"65d576e05376505e", x"f31f2cff1ff73a6e", x"056ca04c52a6188d", x"9aa4ef3fd86d86b0", x"64ce668568f42c2d");
            when 22339516 => data <= (x"74931b62655a8692", x"103b24dad9751e53", x"461768e75ac475cd", x"c821c5666427f4dc", x"dbff8154be91173b", x"badf54fa5600a47e", x"f9abc451cd27818e", x"4f7863bcbe5b2011");
            when 17137128 => data <= (x"a158bb3f147a2f88", x"94414330bfdd86fd", x"ad7f91a634707216", x"ca9735c09c103850", x"230f7e951263476f", x"a09f26bc3fedd3a1", x"b5d1039d3eee0041", x"9a6354f850515cd0");
            when 29375571 => data <= (x"13114531913a5e00", x"da1bb74f8b89bcfd", x"e1d7e3679a25c1b1", x"ff6cde2bb0b4db87", x"c496525867053997", x"d73ee65fc42209e8", x"2258604775eaf13b", x"ea192489ff9a06c8");
            when 6098238 => data <= (x"334cf40a8117f120", x"afe69da21d4deaa4", x"a4421dea6d81194f", x"d1811aadf7c005c5", x"1f447f6ee4ee9870", x"6049ebf1b68e6ee5", x"be965a727d489e00", x"6046f94c4b61b43b");
            when 21525283 => data <= (x"6a9a76726ffc056f", x"42eb8b10d1b58f86", x"5421df7bd6cda886", x"353bf560da92ef03", x"afcf07af08394cc4", x"f1b2737287a8ef3b", x"4817df207f594239", x"129ae04af4d92bb6");
            when 21879231 => data <= (x"c4237fcb9e735e1d", x"c1caa5d093dbc088", x"699a645f8fcff51b", x"87b42655aa1ff1eb", x"374e344ccb400653", x"ca8bd74371e46a82", x"67d4361f9513cef0", x"e090fab3c37682f5");
            when 9125503 => data <= (x"177f617cc1b3e232", x"704244c607748ec7", x"0a2c3e79e5740892", x"b7ba3849722c8f5f", x"6d1e1e3fc9382824", x"9413aed0c0a301e5", x"1be90b87ac209f46", x"fac911751d9f1246");
            when 6491088 => data <= (x"82a763e98c51e936", x"96ba0ba00214fa80", x"9ba22e202e986dc8", x"a0080b07c71d4c44", x"e01143cdc3c2b627", x"df2daf95c84cfdc2", x"a99a9414e1eb6b9d", x"ba9df80e8367dc52");
            when 11691472 => data <= (x"d8a51b8db6249fa9", x"4584e5100a5313f1", x"b75af3826d9382d3", x"7b473e0d6720d681", x"d6ee917a1354a732", x"ce46fbbd9472e3c2", x"fc0a3e7c3ef17cfd", x"168b68a96cf7c6b3");
            when 10191116 => data <= (x"f1065efe2302961c", x"38a05c869259aa82", x"8cf4f052b2bc9eb5", x"255ebdecc6204e54", x"150c3ffe1dbeee8b", x"d601f97fe6de41f7", x"96917572837ffd05", x"2fae9d4abad9e59d");
            when 20099905 => data <= (x"a511a5e13f9f3cde", x"7adb1cc048cf7e5d", x"f4f8b9dc7d7cdc79", x"f234bff58f0a2d04", x"03aca468ce326fcb", x"190a0a84445426c3", x"55e4563233a767ab", x"606387347af7ac18");
            when 25130293 => data <= (x"52a9e62a14fd6a64", x"8307d9651f9b8b77", x"34d4f69955d22392", x"b02ede6393d22390", x"6a5272fc53462b10", x"d7a6f8692206a3fd", x"728f0aad3e9f7ec7", x"d87bbdcc8fbb914c");
            when 24669700 => data <= (x"0939e6697f88d089", x"cff7911d9ce48647", x"21a42cf5189bd14b", x"22491618b3f27792", x"fdc6eae22aea2a09", x"a5ea794ab4b05e1c", x"1cb91f9cb5fe4b5d", x"243107d9dd17049d");
            when 12203949 => data <= (x"3dbaf5513cc2b419", x"cfa65fb51ae1cc16", x"424981b14bf6c23f", x"c396fa52a404d835", x"21ea3697b7425d05", x"0ca1cd1611693e64", x"0fb500fcf4ff9be7", x"f937a2b217ecb5aa");
            when 24878521 => data <= (x"5be964858b08c4ed", x"fa45ff1a94bbd374", x"016c99fb3c9923f9", x"5933507d30cb6341", x"003fc5658d5d99c2", x"b946192074a8bda7", x"a323d5e4ea54b265", x"95fa7f361f6b4350");
            when 31517215 => data <= (x"df0e5a34cb9c1e5b", x"408c8f31161cf9f5", x"5fcf6abe44543e6c", x"2f9a4daf968d83d6", x"332416555aa44185", x"07a2519d47729425", x"b7c0496e8480957d", x"99a32ecf9bedd813");
            when 17559845 => data <= (x"e581045f10183d93", x"7eaaa0cf7e91cf56", x"c341872b58d16eca", x"0bdbf2df1d39afd3", x"dccf3bb3a2753394", x"1568e69e5c8e46fc", x"4c706ca06e83b96e", x"df2a03da033a7a06");
            when 19698386 => data <= (x"61f7ce4c466997d8", x"9e14db5273edba24", x"899adb2eaad1e8b8", x"03126df723ccc2dc", x"d8b3b6befd934286", x"1ac41dd32b01c3a2", x"bec6bf2a5427b902", x"226f507185efe7ea");
            when 21613016 => data <= (x"33244e0a90acf678", x"207fa30470c9c309", x"a8a9df9ed08560f7", x"d0094d8ff3fcbbd2", x"948fa8d9c70b97da", x"c300c03725982761", x"03acd57411d0a469", x"419deaa790ebe878");
            when 15653024 => data <= (x"ed2fc099391d9865", x"8a638d8c07a6a947", x"dd3bda5724899be4", x"3487b0641dfe9b66", x"93b8f1e1d9965279", x"1c4963e79b9dc440", x"c504d7ccc06d6f64", x"e298961f30f6348d");
            when 10543306 => data <= (x"1c52c62d1d4dd82c", x"415f4ada314aa57e", x"a502efbaaf0ee133", x"5f51c1120d7a7b38", x"12d78934840031ae", x"dc73aad37ffa4d52", x"8c86d96b8e8f7380", x"8b857ac324b296db");
            when 1593560 => data <= (x"c05f3fe7103ce738", x"06d8bb97693d83c4", x"f83f960c347ea989", x"d4568505c1d03e7f", x"734bc169ae5b596f", x"11b059678a200dd5", x"c8334a51d1fc455e", x"956faeb4e77b7fbb");
            when 28957473 => data <= (x"87d66b2a8c72c3f2", x"132b4d4353259666", x"10070756fab70758", x"26fd9c87b1b912f6", x"afacc50172bcbb2f", x"2220ec6ca17ec980", x"68f888f12e4cd10d", x"da78455adcebb243");
            when 31759509 => data <= (x"3841c276b688925d", x"d386404f9a2f1bb2", x"60f6e25270b94326", x"530cd5a54cb70a38", x"332003ebe1a9cc14", x"856255898bea8439", x"4d9d753ed5cd34a6", x"d2e2092d87b4eac4");
            when 25300759 => data <= (x"524c0493d98cdc88", x"ad1519759a3b5c82", x"b4d71b7d5ff93bc5", x"29ae8421c4411314", x"e31442563e48bd96", x"d0c18b09501f1404", x"afc0f2f8b3a3cc4d", x"8d0687f54d811c4c");
            when 17380156 => data <= (x"9c7bec3c0b3964bb", x"dada333e745d2297", x"6ddbafaaec41faa8", x"bfb9b87884aef075", x"af92768996dbaee1", x"f52efa761fb14d1f", x"e45ec0574cf85677", x"3828839e5f10a552");
            when 15661752 => data <= (x"1dd8158016de3225", x"fbbd7bbf2b349ee3", x"7c8b830a318fb84d", x"1a283456286ba0bd", x"187f25ba9e5d2a85", x"d0c46b07e06b2df4", x"5c97f9f6761f3fd0", x"0bb78ef4153398bc");
            when 28826733 => data <= (x"03064fadd1d2eb96", x"13b5cc3365418c65", x"b53fd7f2ff31430c", x"1c9c4b4716222245", x"38e8f7f83c039716", x"29fd6cef36185965", x"6d295d9584ebe890", x"a1b38fd024ce12aa");
            when 2639147 => data <= (x"5f6f9815c02dc8d1", x"2b31f4618125bf87", x"a6704891b0677770", x"4eced096be94e780", x"860d1723dc48163f", x"b624a5b679cbdca4", x"d1625bf35ef17769", x"32365c46a765d114");
            when 14445287 => data <= (x"c54f8e765489d7a6", x"f423e0eb15f1e180", x"6c30950e1ef3f24e", x"f5651367865c8519", x"ff82b803ab07f861", x"9ee36a6af82791fc", x"ef054fc0c2d1cd88", x"718fb57e35a4704e");
            when 13350492 => data <= (x"74abe241b9d9aa37", x"69da0a3a193c573e", x"6cd6c863f038eb4b", x"a8f42c7629980518", x"9729a5cd72cd47e1", x"6d46271a1e55d4fc", x"d8e1c9347f8cf662", x"554dc9b963c578fb");
            when 25741609 => data <= (x"448caa058590b7cb", x"fca4406aff363708", x"097e0e220fbd61fe", x"6fd2a05be8175315", x"c1567dc9823ced7a", x"edb7cb6ad77d73f5", x"ac0a60d287b36275", x"499136dd5104d0cd");
            when 889458 => data <= (x"c811e6e78840e8bf", x"d8b43ef962ca52d4", x"5d65222382cedcd8", x"6c0262e26ad9d345", x"3c64cd846294a4a9", x"0c8c24a6e9f7cf21", x"5f7d05aed953b2e2", x"d022e615f3fe7920");
            when 18664560 => data <= (x"5226e982b1fc94bf", x"7b8b4f84fbd70bb2", x"6669fdcf0a9fe1b2", x"849124fb1ad554ea", x"662e0f17598f5abe", x"ed306e5da59c743b", x"47ced000ce9319c6", x"c703aa1ce1c4acbf");
            when 6752343 => data <= (x"1208ff39afb9604e", x"458c7be327419742", x"1296de83ccf8ab85", x"f1e3d42ee1605ed5", x"5217646b4f886257", x"83d97fc50c8e199b", x"605168fefe6ea2fa", x"0a496bc7a08cef1d");
            when 28391970 => data <= (x"4ec8105ba4f9affd", x"f6510eefdd88e454", x"03791b62927c5d10", x"0776d4a150ff497c", x"dddde3257ad26d48", x"983bd6a862cfe619", x"bcc9ea6b9e077360", x"3a903156ed6aee91");
            when 13137830 => data <= (x"6ee43938f13b9f5b", x"d43bf49d876fa891", x"886163b6b5b0d705", x"91d3b17ebbe863cd", x"cfa595d7b5b2a014", x"f08b91fd70e6dac2", x"f65ba7c99bbd54da", x"0ab5a65f70236e73");
            when 3330489 => data <= (x"2e3dce584bc5513c", x"4938c1a479c1cc76", x"7caf6ac4a7805d04", x"49093b65bec995c6", x"932f813d74fc83cd", x"69c9fe3dd53eb7b7", x"2f3492f107cd37aa", x"102c83a7317e2785");
            when 30851015 => data <= (x"5a623c36fa55baad", x"ab8f9bf084612cf1", x"62b91df74603ddb2", x"910dca5c072b63fa", x"e2e71aeb3155d6a9", x"2d27b1a9e8949895", x"c3f7d45555de83c1", x"63fe6f070fe5b3f9");
            when 22006520 => data <= (x"4a0e8c4d6349c726", x"99015bf5518e1e0b", x"3947187566436f89", x"666e0e5fb1bea6bf", x"33c5105625fe9264", x"ba80199dedb2ad81", x"6a61404a45565e16", x"3c67d3dddaccaef1");
            when 32069177 => data <= (x"809670abec276b5c", x"2615b6b9e81c1659", x"8cc837f312844581", x"f364033f7f313de5", x"f818050c1b976ef2", x"211b0dce2c7bcd7c", x"e24d69a6339d481c", x"41f03f6db2894f3e");
            when 9345967 => data <= (x"a6ea742ca6cd5402", x"e2d5ec2bf7fc2bd0", x"9703e3e7a8af5d90", x"3ccb16bf7838fb64", x"6441a8ea6556a9ee", x"49f6170b9cdaab4c", x"8c54bea1154ba3b9", x"4db9f4e3343013d8");
            when 7997622 => data <= (x"6f42f061ad6fe2f2", x"557bc2bed3020c6b", x"73b219d5203c6b84", x"ceba892d912ca335", x"fb90748a95b242f8", x"ad4c5906a2f84b28", x"372a013c8b5c271f", x"3236738d113b4efe");
            when 15085576 => data <= (x"b6761f0e3e3f04b0", x"a7feb591a15e116c", x"81dfda76a8a2dd50", x"a40ba6288f628ce5", x"e842b0c050c137c6", x"e8cd834b1a8064e9", x"2b9a4151c4de884b", x"52205cd2d9966684");
            when 14447628 => data <= (x"623529cf4390bb08", x"76566910ab00381b", x"10053aa31164fca2", x"3da94a8b8349ac4b", x"02f4d9fc5a993392", x"29bd28dc097bcf59", x"11417df49c8514a2", x"01dd7016f83270fe");
            when 30939168 => data <= (x"73c3e05e9fcaeca8", x"8b71731e37d6351f", x"44c1ccd9bb1b96f9", x"9f72696573f37432", x"3dca6f03be48863c", x"99233ab903835be2", x"6f972acf518995ce", x"fdf57a5e959494a7");
            when 33731257 => data <= (x"48545802c82c2fdb", x"09ee1b6b3c5f8b07", x"883d144c7af0845b", x"1289916ad98bedde", x"3cea994a9262ca70", x"f109f4034243fdf5", x"d1fc12c39931b857", x"dd897846ff85edc9");
            when 3366285 => data <= (x"361e322d984454f1", x"99a11e57ae544ea2", x"ba1e8810f549964b", x"470fa55bee61112a", x"d0028955de96b1c7", x"c163a92791ef2725", x"14d04d7fc06ad47a", x"3985fe789f18fdcd");
            when 18969745 => data <= (x"70795ee70adcc177", x"b461799062bd0390", x"97051555de00ee30", x"63406368c6eb51b2", x"787c2f2044e60ca5", x"89115649e9a56992", x"44c71dd2a32cc0e7", x"1e195d14147c7dda");
            when 16398628 => data <= (x"a27eee5590542c37", x"e8f0ea2a29561ce6", x"4194a9d7856044d7", x"dec613354d31ca13", x"e1394935b39bbef7", x"1f5ac576e019ebe7", x"0fdbd5fcda70e909", x"2020c9c027af7208");
            when 25849163 => data <= (x"4c012fa817182d7b", x"346200de8faee010", x"d4c3fdd96da5e9d3", x"43c5684ba05a076b", x"530143f9e57c6e41", x"bd2b5fa32b186c62", x"855ef9b99e086914", x"e8a6cc3eb2f31c97");
            when 28638859 => data <= (x"47fbd0560b47a9dd", x"8d01318400b1ffe8", x"349daae08b6d5c0e", x"9243aa59dd96e026", x"e419ad90953a9428", x"0de437aa6f053334", x"4c894287bef6f709", x"6ace50499ea9ffff");
            when 14169236 => data <= (x"d3b297e2898674c3", x"91f13c941039df73", x"0fbe9cbec1705ae1", x"077433649d5d0c1f", x"d1c19780db9e402b", x"8da5cc55919056f4", x"0473c9ffb38ab58b", x"ae8f52f912edad00");
            when 14019328 => data <= (x"3c5c1f40ecc60308", x"2c873b937a72e2c0", x"d2da2b7c45873f62", x"cacdad136027d231", x"0743b27722eedf66", x"f3ee849913efb460", x"649a715997c41b23", x"97579dc65a5a6757");
            when 2769549 => data <= (x"f6b061c642fb8ad5", x"220298e8bf657c8a", x"a1d57fd9f13fabd7", x"66f9bfd12e201029", x"2135a11f4ec81250", x"86990ee17cca3c1c", x"d4ec773a00a501d0", x"ffafcec4da78ea57");
            when 8666319 => data <= (x"53bbb715ff441fa8", x"ce6b377203793911", x"fbffee3ee9102b0d", x"a59cac5e8d87f322", x"f8f18a363029c7f6", x"201bc771f6d87e04", x"744b902b3e7660b4", x"261efebd59cc3523");
            when 30017901 => data <= (x"bf5e932b9ea79a45", x"2986d47e00af5384", x"f91ac501ffaba6ff", x"02553baf1060324c", x"c98f27f22e842f13", x"c53cc1d9cfc6f819", x"4fa44f2ed494208d", x"0299356751009d9f");
            when 16427669 => data <= (x"a0e1d6642f91c4db", x"6a75b25a62fe620f", x"793bbc28d757b956", x"346147aea66cd5ca", x"da5b7556dfe2e8c4", x"475d9d29b31a3497", x"862591b9d2ddbfd0", x"66291e013de1afff");
            when 26416409 => data <= (x"bccf955f0716bdb6", x"f52b792c706da484", x"bf2a106b12d77b9a", x"b2a440dce85ea65d", x"bf3ca6f403ceb34a", x"1f12d2026752f7d7", x"faca133ef0e08324", x"60d4f94ce2472fe1");
            when 23652210 => data <= (x"8c542d7b79e0e7d7", x"41f60d7cdd411f7c", x"7c03e3bb36463a51", x"079ba12cedf68729", x"ac3ec2eed8e07a29", x"057cef519f067ab9", x"6e099e43b36c3048", x"e96fc2a081ceb648");
            when 20838888 => data <= (x"dd101dde4b4570f8", x"d1bea5a7efe52a30", x"3d4a2529a2c1fc92", x"416d49cfb052930b", x"2de4c26bf74f8069", x"306c8fb5e595c738", x"76c887a3254093c7", x"5356268369d843db");
            when 24777285 => data <= (x"d4fe4a7abe50ef2b", x"6aec287e3eec1b18", x"5d683f0fb0ae45bb", x"ba006421b70faabc", x"058a750cb61df4c5", x"ba31ccf55e09b440", x"5cbb6d4c9801fb15", x"4046cbd68ecaf5cc");
            when 27204869 => data <= (x"e3e764598a45532e", x"1ffc6d99984fa1a4", x"1d0bed16308924d0", x"c7ef6625bd15cc9b", x"9576795c6d014e2f", x"f19b7a0f9597693b", x"207087e3965def72", x"d03370cead37f7f2");
            when 25554608 => data <= (x"57d9f47fa335230a", x"aff016105ecd007d", x"64c14e20987f325a", x"ae8b59cbeaf1af2f", x"e41042b7e2f06524", x"d29e980a40116092", x"c753bab275812e95", x"858d513d04715c14");
            when 22759136 => data <= (x"0a775cbfbe9ce322", x"faab08e77002bcbd", x"6fb683bd1d00d5b9", x"522c4ac098db3dd1", x"d6bd32247f2214a5", x"a556798adf062c30", x"832c846c8eed15dc", x"3133477292cbd21c");
            when 29835821 => data <= (x"0a42bd28ace5fdd5", x"6979350b1d4cabc6", x"5c2ff9f09abb1bf8", x"4bb3720d2e829a4d", x"adb0fb82be63478f", x"0ded6037cb65e5c4", x"64facffc06f9a4ad", x"78b686a23e1295f1");
            when 33198032 => data <= (x"f7b7ae66b6e7fb18", x"da4506079210b17e", x"e3e82bd164326f3b", x"ec0cb2c37a83615c", x"1ac552dbc3560450", x"402c50e655b0be92", x"612374d410b08129", x"99afc267ad7ad6d5");
            when 18632988 => data <= (x"81ed80a0e0a772a6", x"e74aa3b67933cc18", x"3e1132f4eba2780b", x"d444cf67bc1f1a0d", x"715291ca8fabbb12", x"fd3e7894747c0638", x"53e4660546c90806", x"b7040fe3ed01f9b0");
            when 14620891 => data <= (x"d2757cd4cc66747f", x"2237d68daef52709", x"aff104d49e8d831e", x"5b6ce1187b15bdfc", x"b99cc66c12a9d698", x"5ac8fd740fb6f3e7", x"ffe56a71784dfb7c", x"608d73f617e80571");
            when 24207942 => data <= (x"6d2a80ac3660b763", x"8446f6d7375e7ddb", x"8577b9f814fcdb5b", x"d47aad622072fabe", x"2b742b75cba94b50", x"68d10f50cc88778c", x"43a86cf022b59337", x"b83db077dd6ce6a0");
            when 5460842 => data <= (x"15f53f00c8638faa", x"955a0b7f75837965", x"28f2780aebe1f778", x"b49d7199239f89c1", x"8724286ce8591c79", x"20b71c23ff889420", x"15bb7e7bc2ffae23", x"139cc7c1bc1093eb");
            when 13345761 => data <= (x"a82ce42f06f821bf", x"48ad78f5a8d1a9d0", x"48720acba56d96ec", x"ca5ce701b3547ecb", x"6e48f00a5d101a89", x"3ee6a4e4aaf4f649", x"c77ea049bbb6ef21", x"4bf9b1dbb3650068");
            when 31545616 => data <= (x"6be916c77cf9d338", x"1ee6bf0287251791", x"3f7ef1c2424690bd", x"b1206d9476a39802", x"79f906cd183b2e64", x"5fb417055ff26761", x"28279e46a423117c", x"925df73475a72cc5");
            when 12396715 => data <= (x"63663efd0b95293d", x"086476841caa1484", x"eca3f389ec31e321", x"299a3e86a3a9bde4", x"4c51172616afb84c", x"f730f6b2c564deff", x"380cbc4223e1f068", x"d03ee03db11bed71");
            when 27696652 => data <= (x"314078cdf3a9a34e", x"6bb58beea3a57235", x"3879c08f46c460ca", x"fe6f88fd1882b749", x"fdddc6571e1a04c2", x"e8d2e185fbeabf3f", x"898cb1a8a2142ac9", x"b6fd96fece16c52f");
            when 25029322 => data <= (x"000195c59662fb6b", x"8ae0d000a6f3bb14", x"10a87c1801d44cbb", x"074a3e6751a5b5a4", x"6c8ef1ce01ece7e5", x"5615c41cc217b077", x"44e29de290bc4e14", x"9356f609b2c1bf44");
            when 10804190 => data <= (x"54d6382e6bbda15f", x"ab7fbf6e79f6f3dd", x"966f96441ed24d17", x"fe197d736f110caa", x"0735a97ed4031d1a", x"77366d4499c994a6", x"18d9f61bf238f3ce", x"4cf91a619cd9accb");
            when 5176071 => data <= (x"acba1f442f600233", x"6d0549efe982d188", x"b283130de125deaa", x"37a8320252cda5fa", x"771131268a11a8f8", x"99334199c7f676b2", x"86edf48f289acf06", x"49e05ddbbb79f3ae");
            when 709119 => data <= (x"2b4658584beb4122", x"94a5652fa434295f", x"14da8227dd30d27a", x"d409d81df600e0d3", x"be823047a5e3900d", x"31717622e42a25d9", x"3454cb3546a456c5", x"a1feac67b7248acc");
            when 23890879 => data <= (x"acb48a9466ef14c2", x"068cdfacb5860799", x"d180b00c4d372c09", x"d2bf8ffa52faf30a", x"7b1a15a1903f9043", x"5025b505b787cd2e", x"58b265fce71e8fa3", x"a02d8bb045618cd9");
            when 32099585 => data <= (x"a7ade7e1a17c4f1c", x"b0e6f3978aeb8082", x"153ef181886dddf0", x"6f620cff0f90c6ad", x"d5dcb3674281270f", x"8b139f710806e04e", x"f794c6e57071836a", x"ff9b3d861bd51def");
            when 24846573 => data <= (x"20498e3bed75e126", x"eff5689600f4d072", x"c704d841aad88e26", x"4ceeab4a44eb9921", x"66fd86983285ca5a", x"c161cd9c473c4eaf", x"8c06205e295d77ee", x"954f13a3d8b9e1ab");
            when 3583658 => data <= (x"b96a0e3fe4cdeff2", x"9d61c6af8ad6c745", x"9f4c0c4c684eb4b7", x"6bdb33ddd7b42f05", x"4ca1fbd1478214f6", x"e1302af59cde7ac9", x"554b3d134f289de7", x"1ac3e177af60d268");
            when 2335908 => data <= (x"4afeb6042acbf42c", x"9e72a5fb6b283aa3", x"7f651bb9e2a6fc1b", x"37b95553d553ca37", x"67bbbefa0a209738", x"d68a0c6eb91fea21", x"0c40e863dc9d2a90", x"9abe05736a1b4114");
            when 33264264 => data <= (x"0992e8b2c6627f31", x"edfa50eebb3024a7", x"32b50b24ff7d73a7", x"738179b0d7bff4cb", x"6080f8ca1dd798ff", x"11e03020afe7eea1", x"a711e0b5c26896e2", x"6099d5721c291574");
            when 21864727 => data <= (x"2178fa001be9e46c", x"ea8da151057b6655", x"40e118f92a07790d", x"bb612dbf3351b500", x"15de6fdbb6a7ba49", x"22a49aa639c7254c", x"832a9c9d8becb298", x"bd6905e12c05fd1d");
            when 26815826 => data <= (x"5eb28aea90fff7a3", x"ab9054c244d7204a", x"f0837ed92dea5c7a", x"72abc9715cf58b5d", x"d0c3f4621056a864", x"3b6444ff4b483aaf", x"b11f3fd346490e4c", x"c6ca5f6dcc791e16");
            when 7918231 => data <= (x"a8c262b26135dc64", x"b414634e509020d0", x"4da23e3cb5a083db", x"644926d761818317", x"6260e895a5aa9203", x"19cd284ee79a322c", x"c6a182d55f8235a8", x"32dcae3594b124c8");
            when 31062691 => data <= (x"0017e2cbed6f0406", x"25cb664db9107f93", x"1d52996335abe282", x"994a33159bc415f9", x"a0c86155250a7c46", x"f404c4c4109276ee", x"ffd7fef79ec156e7", x"fbb9fe9072cb2baa");
            when 20417059 => data <= (x"a6ffd3d4d2fc1cad", x"ec4a9893ff167bcc", x"b841652fffe3bca8", x"24321a4d9e5f7bde", x"9bfd158bd92e7104", x"c7a7bac9776daf0e", x"5598045e8d93bc4f", x"171be5391ffe5ccf");
            when 18740269 => data <= (x"bfbec5b37ba6430b", x"2a5569adb9798d67", x"d79fd27e62baa043", x"3897b8c19972ba69", x"709e6d0902b4497b", x"6b16eda10e8fe298", x"017fca7b2f6e65e1", x"9b613280cb11fad9");
            when 17608110 => data <= (x"c95ec4ed8d661ff4", x"00ea28a22c92a5f6", x"d15d4d12d421046c", x"ed3538f11c614736", x"20292f1f16046c8c", x"6102a67f23a87c88", x"a6b11d77d303957e", x"525954c0a256c342");
            when 1178184 => data <= (x"90edb30acca14cfe", x"1ee338606eaef7d6", x"6d236413cb1965e2", x"95aec77f74650301", x"303f60cf9b71fcdf", x"4ec372cfd4c23cb6", x"d2b48b00814d3626", x"0b62e4225bf16b8c");
            when 18471102 => data <= (x"1b3b6749a26104e1", x"4a5238c1b6bc623b", x"b6ebfc081c0c5ef3", x"0e4ab32438619733", x"0fdb6ec25609a12d", x"4ea99759f2adfb97", x"ec02a39824e0e05b", x"da1a1ca8ce99d90a");
            when 22391400 => data <= (x"9cb13fc9a4479ce3", x"0862a302329edeed", x"abf5dd31a193977a", x"482b25eee50feef1", x"ab65edf6f5763e95", x"83ee2ba88086ad97", x"8d0840db832203d8", x"d7a420c08f5c1d00");
            when 28664674 => data <= (x"5f68999b9adb228f", x"c6f5ddad81f4e049", x"51ef3e8a7a8edda1", x"390cd269c8711960", x"15b03b6a3e3c85d3", x"4dfdab65521efbe4", x"e0c534de1b761f4f", x"f1168434fb6fb64d");
            when 4216226 => data <= (x"a6210f0e146fcafe", x"8f4e86ec6e5ae139", x"c3922d08a3d202b0", x"9e5f772644bf1a5a", x"26fc73b6d33914d7", x"10519f9585fc9131", x"8447146991565a3c", x"f3b3bc2c4fa720ad");
            when 33377042 => data <= (x"6210461fd7f4cc7b", x"6b8534f3bd7dbb04", x"3776bc611c66bfa2", x"d21c96f7020a59cf", x"5e507b303f5c3e62", x"69568bc479d66a0c", x"081c0c46cb1dc158", x"adb9c84c2d987d55");
            when 19193241 => data <= (x"9dcbda14f8a07af7", x"301993806f7fee4a", x"74355b2d864ae445", x"96cc6d5db25cc667", x"dd7aabb58ee4c256", x"34ea20255030e760", x"5cb02e788593b2a5", x"e5df242814ed24c9");
            when 21390612 => data <= (x"72f6b8f60eeceafe", x"5fc3b9e3fe3a619b", x"b39e2849d3190d34", x"b639cdef76d2020d", x"ba5e3d9f085c5f02", x"ea1642a4cff0f20c", x"336a94d3a4541693", x"e5495caa8ec3c9b7");
            when 19846323 => data <= (x"07413df4aeb8b099", x"28ee7b8ce0134782", x"7753a9b6a513926d", x"c7c3dfd2f24d033a", x"5ae26160b4b49305", x"ea1424dbd72a2504", x"d96fc2f1ddb5377d", x"e0562a2efe8a1aa6");
            when 30592877 => data <= (x"f97bbfd5c092dd6a", x"7c834fbec30bd624", x"df65801c3cae62f9", x"860aac13e69da917", x"9c5a621d7ad88934", x"6bde80b3551bb1e9", x"e614b99cbbca3553", x"c45642ff4625485a");
            when 14132415 => data <= (x"69680eca8254e1a9", x"664a3ab97e6210eb", x"233aa9e019b92f6c", x"87cbf7e7db53cc27", x"ab2f4db6ba0e9266", x"6f21e3d6fe7ae0ff", x"ec9d8d75afda2269", x"5125a9230973fc50");
            when 30957391 => data <= (x"3585b59bfd61fcf0", x"7bc96284ebd9750e", x"745fa22a1944a8cf", x"41bc1a3276c7afdb", x"4dfdec8437751c72", x"1d26c8038f62dc93", x"4cf8153ffbe208c1", x"606a520538ed4e5e");
            when 2232602 => data <= (x"939653a050299b96", x"e28026c54676c144", x"05c60bceabe3bc85", x"8b7e13740e219869", x"0025fc11fe3cc493", x"25789a5100bdd2e4", x"0b7028ff4540df37", x"680fc64ab8cf9cf2");
            when 31818892 => data <= (x"31302db3e0af4c3d", x"71c332f0fc494162", x"35397e7dcaf84c85", x"6a0618cfc95a7c19", x"370854381cc92484", x"978fc947e48d4011", x"044a7a6adbe53169", x"526f5da6472625d3");
            when 1408152 => data <= (x"6aad740ecc27c4f6", x"4d1f5811af21a606", x"c4e38657b3512f49", x"c0203cacbde5e3cd", x"f71a8d22cd0d0266", x"44bee9c1294f2a8a", x"564c481decb79d8a", x"3e94f05c87e6d5e6");
            when 16346737 => data <= (x"711c4a79e6fd6d2f", x"2f327a53a91c5a11", x"4fea1272b21bd394", x"0e5e61ed439885a8", x"91b51a245426aeb2", x"fe93b53162931e54", x"c6fef4de578512f8", x"41b9bbd9144f7fcd");
            when 9336938 => data <= (x"ff292b54f8a24321", x"231426aaff9e5b34", x"1d01a98ca35c4e72", x"eb6d814a5e791887", x"04567505be246021", x"bdb9562d3cf12fa8", x"d3b04bc8473a541b", x"b18bf867e56d97e2");
            when 21568072 => data <= (x"e33fbaabdf671ca3", x"f93faaecaab45f29", x"7dbd0a05cc7d91ca", x"1fa101c788bd41c3", x"04097c35d4646c25", x"7f352aabce201506", x"db927c399b12c86e", x"165ccea7886cfbd0");
            when 17601890 => data <= (x"4f840f5a4b2f1335", x"c8a03682eccedd50", x"185af63431e65c34", x"a57bbe09b0320015", x"621e91c7ed79837f", x"971ee6a138e89a56", x"e7200fa01fd072ab", x"1613d9de4157c26f");
            when 4586771 => data <= (x"bf378e7386260fb0", x"df64cfedc89caef2", x"196b3207d7657ea2", x"d51f1524e77fe45a", x"ddcb1a3390ba125f", x"0463e5f3bb282d52", x"3eae120274b773a9", x"1b601314bf015e7f");
            when 28194910 => data <= (x"7821b6637f49eab9", x"baa9ad425366f022", x"a633189bf3adcf64", x"6f476813a933d309", x"52814481dea4dec0", x"b1c4669a1651e4c8", x"7ed056e4d99be3ff", x"8570d49b196cf7b8");
            when 26849587 => data <= (x"16b421da8fdce70b", x"466122e19dc3f6d0", x"ee727744a47d5065", x"fe1cf702a1b92ae8", x"7e73fdb3ad9f7d89", x"ab707b6835655d04", x"94e53e7697b5a82d", x"b5e1794e77a2ed39");
            when 32733779 => data <= (x"ab23f23479213e5b", x"023e63a634499969", x"b792547e69739476", x"cd06990219efc24c", x"efc7b7247f2caf4c", x"3dee3055c89fcc0a", x"e81aa8754233e1b9", x"d7cd9df37d769131");
            when 18534104 => data <= (x"3e6d8393a853c141", x"aebcb21198ca64d7", x"238a001dcfada334", x"8b2eaedf016d0fb6", x"0fa0609a0afa86d9", x"71f1a523a981d406", x"69f162a6360e412d", x"80c226076bbe987a");
            when 22398228 => data <= (x"50702dab5d23faab", x"9224df253a0bef58", x"364dd53e9132dcd0", x"43499014bb7b250b", x"fb4ce6bfbe797730", x"3fd6125d8be00f04", x"2498639c89a01922", x"a8a1080dd01d908a");
            when 11460318 => data <= (x"b507e7e3f3330bbe", x"32f875013305c08d", x"44f788432b8fb404", x"4ad9649abec8e8d4", x"d3bb05413431f602", x"e070227484791ac5", x"8ab7327bf9a6a8f4", x"ca4398187379a1d6");
            when 25897446 => data <= (x"035a8e5841ed8731", x"a76f1166623e0d68", x"a883d202d194471d", x"648b61a75256cc2c", x"9311290f2b7092fb", x"cb763b8269a5116b", x"2615ee788d5df0a4", x"b4e53744a50d5fb2");
            when 7866205 => data <= (x"f69150d4bc6bc4e6", x"e6c7058c0c23c367", x"c8468158cf5febb5", x"26a0ced5124dc1a2", x"5418e228c73f0078", x"da3628bc5cabda15", x"95adf4c34b1d4e4e", x"40bd4b7aadd8f416");
            when 33425296 => data <= (x"01710d294202890c", x"af50101b44e85b68", x"679dc99e14d05e55", x"8aa84cd55fedcde6", x"b8b99842050a91a7", x"167d2e66ad6c83a2", x"3fb10b47326e4a64", x"9e95ee63115855d7");
            when 17537436 => data <= (x"7c806d54d77d2d81", x"8d1fc14614d57342", x"5b32e230a843f4cf", x"0683277fe2c505c4", x"086b585f2de476c0", x"754ec07c6fe476a2", x"de657dc443a021e1", x"e90da273f2d77b4b");
            when 9523881 => data <= (x"4eaab825188bd98b", x"fbbe995f6cf9522c", x"08e0932ad64d77d2", x"f2811785b51702c0", x"2711c084911ae538", x"3a2efd7fe123af6d", x"7f2b12ff2b5aa074", x"8da7ab03bef857c7");
            when 18653383 => data <= (x"6835f151e53bed4e", x"76d8e9b0888cc115", x"1e20463921949628", x"d3dc23888bcc301c", x"87f19b0b944e0bad", x"f5547859a088cd5c", x"80caba2c9cdaff6b", x"f86c59f98c82341e");
            when 29916710 => data <= (x"b76d233f5286c881", x"0c8b1313a3083ac1", x"e772af8e8adbde55", x"91a3524fbe99be8a", x"3bad2348ed911521", x"b3f60812a8983181", x"505525d30ad23354", x"6f5f298548171cc5");
            when 25886687 => data <= (x"615c88a0c8dd2050", x"dbba938e6d225743", x"066ef15b13de13eb", x"3c8c5df1895a1b6e", x"e21d5f78d66a5e66", x"22c3c5b210dffdfc", x"1e47bd4e7002f41c", x"c112a3a733f7b177");
            when 15077665 => data <= (x"565991e5007bd064", x"773483f7667e6600", x"e5dcd35ce46d0468", x"76aeaa5bba266882", x"9b0239cdca823902", x"76154c6a338f41b6", x"deef439c03cd6ea7", x"982661d637a6772c");
            when 20582731 => data <= (x"ef0921b63eefdb0b", x"f5f19a10418fe967", x"1d0aa424a241e047", x"155eede909e57191", x"4d4a964e423a2e14", x"f2119f26a111a9c1", x"db0f97bc6af17fc8", x"5982408f581f6a69");
            when 26009411 => data <= (x"1f1416476dbfd573", x"f09ea64bbe31d0d5", x"364f1865b73b274d", x"2eaa6f26442b45d3", x"c309299f56a0737b", x"5b3ae06df4bb7ee8", x"7dc86401fc66b743", x"1890ddbf7013f6ca");
            when 24777171 => data <= (x"0159e90591787a3e", x"4d8a09abfd311b9d", x"e7b3200cc6a701b3", x"9c6d6b40ffe731e1", x"c3e5c46551fe8403", x"2d93a7a21b488c67", x"efabc1c68fe1a489", x"005e472b109107d9");
            when 27185251 => data <= (x"d254dcfa28d1720f", x"1c477e18c78e3e7f", x"73127c0bb6aeb11e", x"6ac444f53d763f55", x"6121d20a7f21de58", x"a8ab97bbcc2b067b", x"91ff17777bedd344", x"36b34be684a6e387");
            when 31510653 => data <= (x"34823cc5dd9afa59", x"9a05e9478fb937c4", x"0456b903705c442d", x"c218c6c6c7e0ecec", x"a7ac95238533f547", x"e13e551b61d2c704", x"9b4c2d4a8bedb903", x"9a0a525b84dcbe87");
            when 10817891 => data <= (x"6b2ddba01c3de0f8", x"18c5b5bd00c06ce9", x"3232a5927046a190", x"6d892c851794398e", x"9ad28a0475bae3e2", x"f089e1aef3073cab", x"f65137d54a4c5935", x"5126838d65677a86");
            when 32694447 => data <= (x"4cdcb5fbd772dcf6", x"9edd45c222a700fe", x"1e9a120b220973fd", x"460f5bd59ed89024", x"23b4b377b10b4b54", x"3f6519cb22b04092", x"4ed3ce3357cd0ebb", x"090641d318d32ba2");
            when 33157416 => data <= (x"074d07d760e51934", x"9a0f308604be9291", x"4cd28d2da750491f", x"d5863537187b3400", x"a2878963b116d4df", x"beb465e9552a648a", x"6ad141f63e2a0bb2", x"833088ffce1f3fa1");
            when 3083925 => data <= (x"a2a5eb3e7abf5581", x"f4a2337845706b0c", x"7b60103b417050c1", x"2999959fdeed159b", x"2bf4072a82357b8d", x"c286605ae5353fcf", x"93f879023cdcc824", x"14977d61e483e9c3");
            when 7288143 => data <= (x"f84f3b91d6d70e03", x"43f049120e0cce14", x"b08e63cd7e0389b7", x"a7045d6cbc19d13b", x"04c5fe9aaf5f5f34", x"180ad80c98ba1218", x"c3dd9c7f02bca510", x"f3e21aaaf6f1f4b1");
            when 28233267 => data <= (x"202858734495d981", x"2bf428fcea5233e3", x"09c31db2e2041af0", x"f5bb69c17364cd8c", x"cf82b8d3fba32ca7", x"ff2fae49edc9e67a", x"bcc8851cbfc5f0bf", x"5f07017fe00d2301");
            when 25307196 => data <= (x"bbcffe11284bfa3d", x"e73119d1abdeebf1", x"0fae4941ba800917", x"ab0d9f0ebdb0b8b1", x"cd5b5b247de66dd1", x"79e5ad3eecd94978", x"4d4dc514581d903b", x"c604a68c243aa610");
            when 12826993 => data <= (x"8bf12e5f231493ab", x"926366ece49ca8fa", x"6b95ada2bb5e0970", x"39d7d8caf9cee37f", x"48f64d0377b14756", x"e49b2c72acde5ebf", x"a742d0be0c9df438", x"ea151d107b349c18");
            when 20944115 => data <= (x"4eb3910b4ec720ff", x"0ced47cfe859c2a6", x"0a45be43d25596e7", x"1a6836caabd49813", x"531e66cb767fccb1", x"5dac41c2d4b99689", x"71d83660610fd51a", x"b4fe22f3b165932e");
            when 30960061 => data <= (x"c055587e961b1851", x"876dfc06ee7e70b2", x"8e94607723e72ed5", x"119c68c26d656a84", x"99e44560730ed12f", x"c8b2a6eb763a3ab5", x"d14c4f6e7edaadf0", x"0db6264cacaca6e7");
            when 3297178 => data <= (x"76696e8d3fba0e22", x"73261a8d57a5b0f9", x"2dc4873de9cc9446", x"e940fa12eed6a890", x"73dd90ab738bc1a8", x"d46cf9fee6f17c8a", x"d9b60b4efd495603", x"6a6a1659a447d221");
            when 16438995 => data <= (x"df6f70ddd376940b", x"84e2cfe473cda130", x"18ca1c3a6f303081", x"33c814795bea507a", x"25a58a2759c7c492", x"f6efb7eb669f74db", x"c28a287b2535a82c", x"78b3fb438fdc43f0");
            when 11383365 => data <= (x"b8eec9354d9344c0", x"f80bf84cc519729a", x"7df365a6d183378a", x"dae7136e12ebed9a", x"9491a62c9a41d0f4", x"efe1bef2e29a1c44", x"769f6d4b5fbf6b46", x"325a043c7a674f9e");
            when 4328481 => data <= (x"2293d7448ca4d46f", x"e62f246ff1fc2220", x"af88a032b006f4b9", x"afbf5e760766470b", x"183527f2020a52f3", x"fb2e91b8dbd1bae5", x"ca0aa41c05cc5230", x"2d14c1f835c0dd3d");
            when 8657000 => data <= (x"aec0ff10e9e66ecb", x"2f24bf7ae363f7fe", x"a8d2e63cba6ad175", x"656ae3b9f00e3ac3", x"2cd14511c1fd4d66", x"914823418134dadc", x"f404125db181c140", x"473b91e538304977");
            when 18724113 => data <= (x"51c46137ab341912", x"4d3468b346c224b3", x"f18ab2afcff47589", x"9fcc289f3bf99156", x"610709509f80df63", x"e69e4ec5761738d8", x"d248f01d16f93c34", x"b4b2d51eb5c112de");
            when 9502785 => data <= (x"dc215c47b27aa80d", x"60caf80cd73a4f72", x"0032f2ce8af49d71", x"80dacb5a672ab145", x"6324ec56122dce35", x"4c2bd83a1c48f603", x"110060a4bf4752a9", x"619b7e4f5579c75c");
            when 1277430 => data <= (x"2c1be20aad887d27", x"2f950f84cab2cdd1", x"c2b12a5d4c31251d", x"f8e16d14afd8df0f", x"fab6bf5432337ad6", x"e17476346f87046e", x"dabd55d1cac26c0f", x"b666575605a1f4da");
            when 27565102 => data <= (x"d08ed48996aec55f", x"1b42f22229d56ff7", x"4fc5f7790442a1d4", x"2135e3e3a4cb1db7", x"8da7a09e4490c386", x"aa3fe0dc425a618e", x"f8b3cc5992c343e7", x"91a7725132e9ecca");
            when 26588427 => data <= (x"154d952827a0974f", x"2a17834f31a80123", x"eb2fbd48755f75cc", x"fbd85f37584cd36f", x"d15fbef64e34bc3c", x"4d537ffe4b19b0bc", x"359a183e1c56d266", x"f3e91c7b91e4a7cd");
            when 33346163 => data <= (x"e7ce3317be908075", x"cb7f240f480fbcb2", x"2cfc5a77681e6339", x"a7b7df5fecfe781a", x"afbc466421ca20c2", x"ecfb565c0ea9d2ed", x"fa60be3f023ee06d", x"3d23d0e180589c7e");
            when 19519403 => data <= (x"f7b5d84c2b44a482", x"ab43cd3e0ae8053e", x"67aa291dccd24638", x"c1ae66d41a236241", x"e9292fef35d1dd08", x"2eb23a8a09410f58", x"cd68eabf02502fc3", x"fbe764617662a846");
            when 15658209 => data <= (x"5b0edeec58126e2c", x"c32f2805f167d59a", x"abb63a46f4639548", x"f4fe22a7146d014f", x"38bfb5947d1cea15", x"0d6bee6a2b3850f5", x"bab82fc7cccde769", x"de1e9856fa981f9f");
            when 31292117 => data <= (x"802d5257b3f4177e", x"fce2ded0cb777e30", x"10f4ddc7140f74db", x"a033670abb0e0b26", x"9828fe0117a6deb1", x"428044a106326a5c", x"3642a8663b65a97e", x"e49ed3c3a03faa92");
            when 12208779 => data <= (x"8e6d55d9c3e9c48e", x"34d7e02e7d781bed", x"c814085b21477142", x"68cc3f13816a19ac", x"a18dab3499a87122", x"8e46e44aa10cf1d0", x"f0ae9de622bf47b3", x"9f8dfb8e227be252");
            when 22472729 => data <= (x"c29d25ff30dbccaa", x"06fcf8e9ba7e99a8", x"c2581a05256fbe0d", x"68f5e8c192748a80", x"e78f270fcc31fb33", x"d9b75a92c83d4e28", x"863bb20c8c1d9343", x"2dec58207d7b68f7");
            when 11157527 => data <= (x"8bb2832a0543c322", x"096c9e044a732825", x"efad5eae96ecbb46", x"db4afc857665f376", x"8eb234635a794d46", x"fc28f0a2fd5ec1a9", x"3360d9aefbda91d1", x"906146f12d6e525e");
            when 4597460 => data <= (x"f951138bd3a72741", x"543fde582b7629ee", x"7ccc7659b98299b0", x"928d35cecb2e25ab", x"e765770788abf18e", x"f88750d8c14ea078", x"8014335a4d936646", x"5c82ed9aeba5c599");
            when 8517997 => data <= (x"62ab69e7d57fc020", x"e09740b05e57627c", x"005fb3d027550dbd", x"187faad487795ecf", x"779630859b6c02a0", x"7db859daaa6cce74", x"106465ddbf96e626", x"709c1621f39cfbbf");
            when 14615488 => data <= (x"f92e9eac4d40ee17", x"f668c80b79f7d2bf", x"3c4de44d2c5a19c4", x"412ef2246f9e8281", x"a0a9fcf17b654a74", x"83f9a31f985d95c6", x"cb6f5363500c1139", x"c97e621e4b42c2e9");
            when 12296824 => data <= (x"fefef2ab9c30e1ad", x"320e280e143b2512", x"137b2f78e93ae1d9", x"294f9cf4b3e49e36", x"e835327bce6324aa", x"e44db12a6c9ea528", x"5b72ce495d07968f", x"b9fa6d5e953b00ee");
            when 4908639 => data <= (x"c1207d4db0e213c8", x"e66c4dd40c382613", x"20d3c8b8dba1032e", x"d3f23411b0d6126b", x"e2eec950fe734d45", x"90bd0e87530cfb2c", x"90a3bee9bef9e716", x"255a897f7fe844ac");
            when 14903581 => data <= (x"8692494b5223e1c2", x"b51a2c34571da7d1", x"d152563a0f4c0e5e", x"6bbc291610b7346e", x"f810dadae3a5c099", x"1eb5d8e093ec8be7", x"12f73ab970c05942", x"6ff2fae6ec7a4f31");
            when 29850141 => data <= (x"7973d62211129072", x"8011fba079812da8", x"e10df86e922ba1bb", x"4c7a4bf73d432ba2", x"7ee132560156a6d1", x"cd4d622d8fef7afc", x"b1f745aa4b8b7d5d", x"bcc7af8ac6d0758e");
            when 2027298 => data <= (x"2a465aceea9630e6", x"f3366991367ae727", x"473d173953da31ea", x"50a3b1660e6e2a7e", x"4f25e1f7b97f6582", x"176b1adfa1593391", x"c4b0d4b32537a5fb", x"53e853a432ffe6da");
            when 19460932 => data <= (x"52fd037beabc438a", x"29275a50a9e54b4a", x"632557f7aad22600", x"45a9138bd19fc637", x"1f1431bd20a388cd", x"81ddf3dd3af4c5c3", x"dafab55664be710b", x"9e9fb574ce97f1c7");
            when 24960855 => data <= (x"f7b24a43512b1d0f", x"f1f718d8d2ed2c04", x"579bcf4907b13f19", x"30b8c734c82919d2", x"482982b8993e8e96", x"3cbc043453e0a782", x"d683d674c4137eb7", x"cb8db41768f0e0e2");
            when 3852017 => data <= (x"7f69e9fa2cc02d56", x"e2fd35dea8989922", x"202edc1477b3e2d8", x"f851d783e5e64030", x"edae7b2fdcb09530", x"69dd620b517b8743", x"ee155e1681c01427", x"b7fe3601e1f8ba42");
            when 6874458 => data <= (x"a95df3a4fd6b10d0", x"bc32226042e25d72", x"7284c0d867b1c877", x"1c02121a6df9508a", x"459a9bae87087b20", x"7890d03d90c1cffc", x"68d14945a3477204", x"06021030abacb084");
            when 22665199 => data <= (x"755ab9042d957f75", x"9406b52f7dcb8c00", x"f5ef519f893fe175", x"6f873c6aa661701d", x"6dad7d6a571e42fa", x"9b81fe1136b7f43f", x"83ceda15c9279f00", x"892718830b7dd81f");
            when 13069496 => data <= (x"dcbd3c429e0d923a", x"8a7f1e340c156766", x"eb29679410b6a389", x"60c5779df9017def", x"cf26daf09e073a53", x"a340a4f331a10f2a", x"2c20b48ba6eb5297", x"61aed1765efa3f7e");
            when 17200729 => data <= (x"80519dbf23b25951", x"2c74afb923645d2d", x"dc4ee153a4002e20", x"47b41c65303169ca", x"5af9efeb73a78b0d", x"815f9d80512a75f0", x"9376b09fb535cf64", x"1349e84dc75fea86");
            when 11228017 => data <= (x"8b7f7738dfb9b0de", x"5f2839bd532cf323", x"421457e27ec47423", x"b56bb1de27089fcd", x"9277e043f361c7a3", x"17c01772427451dc", x"b8deea5c317cb1b6", x"ad2e3412d8ea7245");
            when 26365665 => data <= (x"2b4d59c71663235d", x"5929d64b7c773c28", x"587fab898bb39cb2", x"d760200ef6926b55", x"3a2fd2b4e460ec22", x"697e40d584f50c73", x"feefb912f3da90ac", x"011e9cc48b498e79");
            when 12667544 => data <= (x"386b4b378aa0faac", x"0569408d766bf401", x"18b72270999c0a3f", x"6b90afa700d45168", x"cfdf4cbcbc87b23f", x"5a9af0b677ee97da", x"4bafc95a1b5c3125", x"daa98e5699b2500a");
            when 5473415 => data <= (x"5ac374a602008ac2", x"0b3187a0d16c15dd", x"6ca6c9cfd2e74fa7", x"f7a011b48e27c70b", x"65ca47012be46086", x"ccc6492e73d79761", x"6f7c770a9f5552e8", x"b4af780723d1422d");
            when 29350532 => data <= (x"f123e65915764927", x"e61957b087b97ea2", x"62b6ac86c1312e78", x"a3ad55762d3bd6cb", x"3e150a6d3105d457", x"f5962c4f23e8063f", x"fc058f78ebf51f1e", x"fd77220ae445dbb2");
            when 6504464 => data <= (x"af7f3d8f70d0718c", x"d5ebc4029c5ab3a6", x"99f1ca56223bc0d1", x"e735f935bd732396", x"91573bd8078a0a71", x"21301658297c1d0a", x"3ccb37edad4df6d2", x"6805bff8df50bb2e");
            when 22712315 => data <= (x"84f474bbf911bea5", x"e33f1fbeeb72cbce", x"70f7f233cb2cdebc", x"2b66e5e065cdd9aa", x"38ffab7d52ac8ce5", x"dd9c33468c4ed9ae", x"8f6bcb6a0d13d6cd", x"642edc20c47a3425");
            when 22921254 => data <= (x"42798c40b31823e7", x"acd458e63dc5cd36", x"247a4b65bbb0623e", x"751bb108f0393565", x"c0174df4af29d912", x"8f8e6e1e3a91ce8b", x"97adb5c16482d993", x"566fb988c1f000bb");
            when 20716644 => data <= (x"9e49694dd3fe5ef3", x"a02bb7a744af283a", x"dc24ecc74d1fb77b", x"6fe25b16bebdc135", x"14a5c2d88814cdd3", x"41cb2dda8018a93c", x"7de323c86a01a63e", x"69ce101ef0b295ca");
            when 6041035 => data <= (x"b559b9060b0c8250", x"a0004427dcb382a4", x"9d208a733fc22334", x"1691e25dead9fb3b", x"568246e127aabbe7", x"5563f569bb076520", x"681328f7ddb6c240", x"8fc7731e030ae337");
            when 16954023 => data <= (x"dcef5f1ee4d63dee", x"bf093901643efe19", x"ecd5406fb1565797", x"21c1443eec6c3aae", x"c7eea13143a1b9c1", x"03906d8938a0589d", x"fb40917265d309a5", x"a4f2e9754bbaf400");
            when 28792578 => data <= (x"32cc09bf0eb42b8d", x"163663e422be2ab3", x"d1d03adb4d1890c8", x"b037ae8c789dc9cf", x"ea252051d87fba93", x"4e7f4a906aebf8a4", x"dd910850a6bc20ed", x"dea45dfaeee790ba");
            when 19663947 => data <= (x"a639ca00c9c8d4bb", x"07c1bf76bb0079d9", x"1ec9ced772f9d4be", x"e1f463281bc18c40", x"1bc6e09ff7557088", x"2bac17d7bbdf2880", x"591d7cd156255497", x"a35451166334745d");
            when 19455341 => data <= (x"5fadb38fcad83758", x"d7c38d6a6063c10c", x"7f84b91075c47f89", x"69c670a597f58429", x"cfeb9518efe95cc1", x"1c104ad915fcf899", x"96a92f1edf476af5", x"8dc9cfc419521fbe");
            when 2108751 => data <= (x"b255f999403d082b", x"2dab86ff9f9d1c0c", x"f53ac10e4499b34f", x"97ad7a1991120b0f", x"022694283a8a58ff", x"ceeea926e59bc523", x"9951de3be56abfa2", x"c437c0f8fdab3b92");
            when 5534133 => data <= (x"bdccc98974f4309d", x"2608cf596dc298bd", x"6323a92eb15ce3e2", x"73fb62cb90df9a39", x"3ab249fa73158b5c", x"eb0d187e4eb953df", x"2ad812365a6bb09c", x"312f21f96668ee78");
            when 10283719 => data <= (x"fd43b076f08e51d4", x"19755a6a1c63d8f2", x"6d203259fccbfafa", x"e9ed05050370f941", x"fd95bb4077e10930", x"cd321aa973864eba", x"3064177725839d7f", x"15e32c2927c4c1fa");
            when 33246267 => data <= (x"bfffce38c99a85ba", x"37a53e96d325f2ea", x"b45342bfd0537633", x"ee921b0076d2561e", x"c9b74c976011098f", x"9e842387900c4a19", x"6c49a1463ad8e875", x"0dbb3beb136d552f");
            when 23154258 => data <= (x"2e04c576ad4682e1", x"71fad22750cb9697", x"b4cce345a0a68207", x"3af64336b2994c86", x"a2aabe2a14cef39e", x"821ae3dc26b8c042", x"4873895be01602a8", x"502b22b1ca75b88c");
            when 31950520 => data <= (x"6d6e0f7bae12a9cc", x"7ffc0ebb4106a069", x"228566006d1b1626", x"1e33e135d4ba812e", x"5f92a9c2b57d337e", x"015d61fead9e59de", x"8e04a218d68ed5aa", x"11f78b8f27247aeb");
            when 19098401 => data <= (x"8919b30d964f0f38", x"0ea9328f37fc7c3a", x"9c877473e55e7183", x"a2edc3ffba68e6b2", x"933ae5e91af60b68", x"8fd18e90b7774b73", x"df04bfae3d61ddce", x"11083547322d192b");
            when 32310686 => data <= (x"579fcd14ff52ee7b", x"a8f80b6184e60ab6", x"06ca13f69b9e8c81", x"86237bcec8b23cd3", x"2ed75a0b550b44ad", x"c46d09bbc7b8f78c", x"8a17a9f4b510df8b", x"161b56c5992b0c7b");
            when 26774721 => data <= (x"71e496194f62429c", x"81a74504a2074857", x"f1526ebcdac633c2", x"9d114b67f0e84ab6", x"a022db7078e674ce", x"7e43e07e6fcf70ba", x"7f6469cf7b518bf6", x"c13a1fe655fe2a9b");
            when 25312928 => data <= (x"6d9b56f0ff96a2bb", x"588b6288f34fd3b2", x"05346592a3ea0b59", x"c2a64c00b1ee706d", x"a2e6c6fe2013a0e8", x"749a5f1b4bef756f", x"2448bb77bde29283", x"87a11739971a9956");
            when 10274914 => data <= (x"f8aa35a4d3018518", x"2c097f7582470cd6", x"d8651c5d70631815", x"c1b10e8498a2d90b", x"7ec5dc55ba1cfb8a", x"9492b2e5b4f34aba", x"d589c9e73db675d7", x"f029fb628d2f87dd");
            when 26779862 => data <= (x"694bef4b063f9f8c", x"b6721f117b655b95", x"5b930c05cbc95e8b", x"a633d9b5114e26af", x"f60fd0b31cd282d8", x"694e26b565c9c9a7", x"9c7f8f9908a66ad5", x"32f6761d78be2e26");
            when 26682883 => data <= (x"73011c28a9f2117d", x"3f186bdaeadbe64d", x"cb791a2f1323f6a8", x"5d1137747cd3245d", x"134fb6a3617579e2", x"eb86a389b3d6c600", x"96162b5a52c9d6d3", x"70e26e2a715642ba");
            when 21132164 => data <= (x"049330341b86286d", x"bf0a3cf53d7b836b", x"8fec15ddc852bb84", x"b36cde854b8a9d8a", x"f79fef19e63ab0ad", x"36b1406f578d7d1a", x"7341a4268db0ca62", x"54340af0a53522cd");
            when 8922805 => data <= (x"c89cd70f374b0ac7", x"930e6b4662ff8c35", x"bfca3f1f43beb083", x"ddfb30d95dacd156", x"954b51d1eed4195c", x"b3d4cf9825827b71", x"a2ded7a46bdb4af4", x"95d779d9f9b0f4af");
            when 7048550 => data <= (x"82ee8b8a72035864", x"adfbb934dfa192cc", x"c7d446abf7b8279a", x"959e5f72b567e86d", x"c88474877c8cd466", x"7a939c09c7d6a7a9", x"2ebb56bb241db3e1", x"4522fc635fc3f6d0");
            when 10825265 => data <= (x"aca15da14e4b23c3", x"32a8292cd2821992", x"a5557203b9995067", x"a9827ae0faba9889", x"87c2aa77448ddca9", x"9f61dc0b1e28c1a2", x"a3f286f2c0b60c71", x"eb92e865b2ca65bc");
            when 14678471 => data <= (x"2993d3f9354d91ad", x"24771a9928952a6e", x"9457fc0b8ff2bc10", x"cf194b706285f172", x"88b9a65212e4e2e3", x"362333116b027447", x"73d521dfbcbfcc2a", x"ce908d00cae5d5de");
            when 4591596 => data <= (x"d31fc8209ac1302b", x"c451d39a71bbca50", x"8e15b73753252013", x"f9e78a4276e2ccd8", x"7afc2df6c9190aaa", x"f4f50d32dada3806", x"b861fb61b8b3a95c", x"ac4153918a5a04d1");
            when 6682576 => data <= (x"f648f25246fdf700", x"28a0e213c9dd0f93", x"3ec6b67435bfa5be", x"541f1d8f153fa082", x"8de3f54dccf9ad61", x"897195fe752e074a", x"7984c8b60887fe78", x"9ad84d87b7f184d8");
            when 3500889 => data <= (x"2efd9c734578906a", x"0075bbe227b86811", x"dc0f49e720e8592a", x"878443c67b30927d", x"9d6eb2839ce40367", x"c8c1a19d1aee82e2", x"aeda35fa46758752", x"c233348b424e5de4");
            when 328688 => data <= (x"ef77fa4b60449eb8", x"42e7d0be2a8c41e9", x"806e18caee574201", x"7e39f0826fd14674", x"6476a240a95acc50", x"18cc6617a00f0a55", x"4d80fa78e681a1ca", x"fc7e0a89e1feaaf5");
            when 5837153 => data <= (x"ad09bb1cc28e277e", x"b5788da77755094c", x"36cc088550902f15", x"890425dfa423b8a2", x"03c88644c930970c", x"d742cde2505bd826", x"79c774c9b92df803", x"1063beba27f9fe9a");
            when 31135772 => data <= (x"01dffb8ef9c09d3e", x"132a068794888e20", x"0bb91fcbb4bda282", x"dc4e0a2209af6b2c", x"6561aa52b210d50b", x"94b669d685f544fe", x"7ed132cbab044ff4", x"d6a457212634200e");
            when 29536560 => data <= (x"bfb2c85f8c4d396e", x"a282f8e60cf0c344", x"d56246e80b8a9214", x"9402d5a7fc67ef92", x"86263a9092ec981a", x"faf2cf7f56eb1918", x"5a567b5d7213409b", x"fd908a11d8f38f6b");
            when 13087466 => data <= (x"363eeea019aec7bc", x"a128af04f02c92d5", x"31f298d00842e725", x"01a00f8b0274ca8c", x"80b3c97bcdf1a804", x"3a10b70eeece204b", x"21818f49ac1f7a95", x"e209f931ecf5be21");
            when 24909478 => data <= (x"07c2c8b398cc19be", x"d06420acfb1f2880", x"aa45489af177ab5c", x"bcdfd6ad8e516d44", x"d47c726a37659e28", x"1e383e418dcae73d", x"eaf9060b7bbe45be", x"e73f592b97013ef7");
            when 1720322 => data <= (x"a895d2462d0e5469", x"551bc5f12f3e7ff2", x"9296603cf57cd6da", x"58466ab070492117", x"725071b2482fb741", x"e687b8d333df1dc6", x"d41b9dfb0c0c0d9f", x"60ceb14d033c8f1a");
            when 25449788 => data <= (x"fa4539bd19dae41e", x"32276ca105f228d7", x"387ed6158ba56ad1", x"3a7fe66e10f180fe", x"25c81d7b3b78d247", x"2113805dedf6136c", x"b0369235e5c6755e", x"25914db35cb607c7");
            when 33353774 => data <= (x"bfb76a72989ef9e9", x"a09c352417ccdcb6", x"150672596bc69891", x"ac31b24d3fc61c98", x"7175e6094d34f885", x"8919302d8e3bbdeb", x"34efd10e000ef3ec", x"f9ef5f0587afd732");
            when 24847321 => data <= (x"4770bb1f1a70ca84", x"7917ce2959f3f600", x"9c274d703dcd030d", x"8d9cc2d0be185bba", x"323dcd72a230fc06", x"428b79b2bf9f4053", x"6de24fef0fa24171", x"a4f7547b6f17d6b7");
            when 13497475 => data <= (x"c03b4bf6c160d151", x"27e9d1f278d024c8", x"2322aa0989bed183", x"e419052a141cd3d1", x"638190df25fe2c01", x"d4daaf2dcac63aed", x"ad210ee8fa05c416", x"42c7a08e1b49553f");
            when 1060804 => data <= (x"fa3edbdb43a33f8b", x"63116b2b7e2897b0", x"b43246fca65730cb", x"3e0f2490a86727ff", x"0f75110e3e704c39", x"28f366df4b625312", x"bd8a7c06030a969d", x"d08fe02c180ba782");
            when 8089859 => data <= (x"0c12ab12ee29d79a", x"0d19651c3d5cf1a0", x"ecb01d7e6bb9aac6", x"42340f2ae446c03f", x"4b1c4facffc68ada", x"70ecd5a2a34dae4c", x"278c23a630346b72", x"1ca43dc48da2b457");
            when 28521657 => data <= (x"6d93639e2fc6fbe3", x"6c2e086d57b14ccf", x"064794018131da2b", x"21b2a041c35b972b", x"7820e662aac10efb", x"709f81d2918ab60b", x"5bed50b670e78a6a", x"fbad33d9a162c074");
            when 30880305 => data <= (x"68709ebc5a9ccdbd", x"3e001a5639bb5026", x"4426aa83262e1600", x"8de5a0d8a52262b3", x"dc4332fd7ea5e2e0", x"85fb7f896733e020", x"134ad27b487a512f", x"f4d1a6f279d4bae8");
            when 10780265 => data <= (x"a4fdca1a33085edf", x"52b750d90e7dd09c", x"2abb8a5af0c4b7f7", x"5b312779a2789f6e", x"d28b05e0a89e3070", x"178b19d8a4163b57", x"604898805e8363ec", x"0b33f3c721eb2ca6");
            when 13759947 => data <= (x"fde6139f038a4387", x"2a95a497457866df", x"41c05401bb96d4ba", x"e244c1ad3931104d", x"4de3230b99179af5", x"24f6ea7da225a668", x"0a9772676208f000", x"c3b10683cb6bb7db");
            when 6752431 => data <= (x"a1b013ce4a06219f", x"826b863f31f559c9", x"9c53f84b22b5b53a", x"20dff2e8addac474", x"5e89685b636239c6", x"ebbfda18656d816a", x"d1a45325cfd20454", x"48acecc218e93bcf");
            when 24237940 => data <= (x"10a22027b436c10f", x"4b1699d2aa5ee595", x"20d8ecf09138d69c", x"1c99036571c5f3db", x"770b8f3ddd1db9d6", x"9a28987cc7022883", x"838ce577b1f1a2ca", x"2a96fe6db3141809");
            when 9813608 => data <= (x"029709983f9f13d0", x"bd0983775e6dc5e5", x"bb0d0c33f248b55b", x"d04afeb5e0709326", x"3a8df79a6740b045", x"de168eb839b7341a", x"13ba78870b713b55", x"cd8e8badb2ce71d7");
            when 20831584 => data <= (x"42c0d8992dad95b3", x"a5492cb7b6746138", x"3dca20064037e8aa", x"ecdcdde199b8d6b6", x"77e96c2cfa76d100", x"0aece26a740e657d", x"9ffa01c3ce422069", x"27bd490611bf8fef");
            when 30182809 => data <= (x"54e418c7efc7ff5c", x"6f5e264f370aefb0", x"7773e55f701c395c", x"70f1cb61b4bdde8a", x"66f28accca1c9b74", x"7600278e04665efa", x"2bffe33fc1fcdd8f", x"db252e25e42bdb77");
            when 8050791 => data <= (x"70b8dc1ffad92722", x"aff5039f205ac6db", x"c42e558678548ae4", x"0ef7e1545b0b55d7", x"08933d1078a7f886", x"9443862df2854c39", x"6c37ce08ce5c93c9", x"8b663f88ca03d716");
            when 4325763 => data <= (x"4e71f5058da8ae01", x"93445cc0e3c74c6f", x"b8637b272ac4b5cb", x"0b9f7ba4017effab", x"630444cdd69ff720", x"0c5b082b3e3feb72", x"a7bd9cea065f0f81", x"4929e9dc568db2eb");
            when 29175277 => data <= (x"7efd97d7b603b77e", x"81deba5586723ca1", x"9129c4f86a58d3d0", x"1e2ea6767b47812c", x"ea4ce9f871470ab4", x"2708522add94a662", x"80f3828e3aec511b", x"c91ece0a6acc3d39");
            when 21079991 => data <= (x"aca12db685ce52fe", x"28d8b959a34c264f", x"e2936bbc90c56fae", x"08e046f22f23e121", x"5112ebb033915c1b", x"0883fb6201294417", x"3953032d0c512db7", x"108def7e98e0f5d6");
            when 11676056 => data <= (x"accb7b2cfb4b7868", x"011dd3600c3faf47", x"abf19e9dfea592d4", x"7ebc8c75bb16edac", x"3e7ce7c2cfdfe800", x"b627042c5a92215a", x"6688ef2ae2548cee", x"d0c736fd66a19cce");
            when 22599584 => data <= (x"8d74e34a698f911c", x"d64655fea69edf5d", x"9f582227ea0e1b7d", x"f0150461638ed9aa", x"58608f4c46f7928f", x"586af9f8aa05b184", x"99fec509713d258b", x"29ea94b4a978304e");
            when 20626472 => data <= (x"743ccd8b80de30c7", x"29a5278db09b1031", x"3b04d839376f1ad8", x"a741a9069c143125", x"95d7a872897b687b", x"0ec75ad8266a49b3", x"e00f86fc797a5103", x"90be14d872ea107b");
            when 32040677 => data <= (x"b541e5d70d7e0c90", x"1004c617e12c9438", x"84f6970a519ef0bf", x"702ddbf3ac278d1d", x"9540426b5a0490b2", x"e0fac38ab0fcc6f2", x"a7fbcb936a225d03", x"e38825f9863e1e80");
            when 29473710 => data <= (x"20afaef0111e15e2", x"f159ed90df08ad47", x"092ffac8150b07eb", x"996854ce02811064", x"bfc094acc6c27523", x"c6ffcb509cc23af1", x"01f3bcbf0c992a59", x"498a3be4ad85f3d4");
            when 19798101 => data <= (x"0790b21f6ecc2f9e", x"5b5fd3866ee9b11a", x"c5a713584b55597a", x"faa8d4ab08d06355", x"6e205443002cba1a", x"72b6b1b514180f28", x"51bee078859b8184", x"3a81cc81b9380606");
            when 26158921 => data <= (x"0bbd5f89b6ea9c95", x"9a85377c34e4725a", x"d721fa08a849a9c3", x"5d925d0f4c296f81", x"2493aef6f3d50ae9", x"87e1034f79361ee7", x"8d5d3eb957fd952e", x"e515ef559493ab5e");
            when 21289983 => data <= (x"b00db841081dade7", x"9186cf62d29130e0", x"1374df835f3db09e", x"683bbccaa78e2c6b", x"91ecea90905d4f0b", x"1df7f002c78d22c4", x"d44b13d2c03e4c92", x"a3bd1beb04e5080d");
            when 23827913 => data <= (x"6b3e24bd7f2fc3a0", x"746c782acbb017a3", x"96cee4b2b606e4a9", x"43a0dcc74d617f71", x"27543117377cf7b0", x"8c1ced4cd7e27c6d", x"b1f1f94590eb2950", x"b3b6e66fe474364a");
            when 17282184 => data <= (x"daf2768b7b8781d3", x"7e0ba5587424af29", x"a524132bf1cdc616", x"7e0c1769dd20ffeb", x"53318922c92a2f9d", x"92e2e604ac364532", x"75c4f3e1055865f8", x"a68acf8eac40e2e5");
            when 12408061 => data <= (x"e336eafad948e8c6", x"098dc5029e2999d0", x"f739d85aea940ca2", x"3f591b8b44dce32f", x"e5e88e5e4a5ea34a", x"deccf2d8a7e63f13", x"77ffc17c57e0ce44", x"1eae7306ab7274e4");
            when 29276611 => data <= (x"f430ba78d7422073", x"81dea2e947fa4511", x"95f279e495264200", x"ac221178a31388ea", x"97a90720c0089294", x"81703e0e24c6422a", x"50cd6f38e3dda9b5", x"4d3869e8bbfe5436");
            when 24948753 => data <= (x"39ab1f2cf112c4b3", x"dcaa5d42adf91575", x"56d97ca2048dfc21", x"b5dd90a137de2727", x"f9f7ee50cfe90d98", x"90b2f49dfcbc2ad8", x"2af1c0300c9f4642", x"71993bf7221af472");
            when 30623537 => data <= (x"fc555d6bb1b60ada", x"9946f88be769b49e", x"7029e29ce32e23ac", x"db490a5de51a233f", x"24e5a58ed8420477", x"d76458b210ef91b7", x"150d948e68baa075", x"52f55bd1e831bc00");
            when 32220921 => data <= (x"0c15146c2e33d81f", x"0f4f2b51672bc618", x"f5a24d5e8e7d4a0e", x"852f8456bb7ae4c3", x"ec6bbd2c5958c834", x"4e22fe22d586039a", x"30a3add70a5fe136", x"9de71cce123f10f8");
            when 12369130 => data <= (x"b30ada21bbfe9ca0", x"08b69446209aa21e", x"ecab703082838e90", x"d7c7eabe236677cb", x"b582204a77801024", x"5aa79a16075132f8", x"b3e7dd01e20adbc5", x"09b143d76db1d8eb");
            when 6605619 => data <= (x"0ddef16720ccb598", x"4181e3ea42e23bff", x"4ae92d3b0c725316", x"04226beee4cd0e96", x"f2f8d0107c3a3a6a", x"9977a02c57a364c7", x"559f043d0b858fd0", x"915b6758ae874004");
            when 16287969 => data <= (x"ac632f55c612f36b", x"51e02b1581015290", x"6c781c1407c1e25f", x"b4a731217e6e835a", x"8fd01e529d95a40c", x"7f5b2cc29d6d4023", x"97bdd442463db199", x"74d0df9100b9b478");
            when 3970041 => data <= (x"09a402b0c627ee09", x"3d074ed105d56ca2", x"8a98ec4cca6dcb7d", x"a8e2ba6dcf839e8c", x"d4bd968a016944bc", x"af87359993a77575", x"4c597a9849255b45", x"8d3aadd32c70ed13");
            when 28268182 => data <= (x"1237e728e67d1b9d", x"d2797e8910118c2d", x"d18af3dfcf07cc60", x"a6a8783a20e5cd3c", x"6cb115e6f7f491c4", x"5db40ad04b199d75", x"1e7bf78d4942aa68", x"c686da644f7a06e9");
            when 11275385 => data <= (x"7d2d7fe478d4e646", x"921b000f937dfbe1", x"13b3ed8e8e3e6304", x"18b75a55a0014c3a", x"840e8de5c6190685", x"4013412dfc49cf2d", x"ba2d8f55ead697bf", x"a986f5590380dc86");
            when 4563296 => data <= (x"a78122d4f7264aae", x"96053101a5a7a60c", x"97768ce3f6b1a032", x"0dcfe4d8ad5e4839", x"206590c23dd1ad13", x"6d188ebfa6a2bbea", x"45f08556784f60fb", x"62472981e5b71c90");
            when 27140916 => data <= (x"cc8f8a042b80ee6b", x"d07159320ed2abf9", x"f7e6965583c83130", x"0458dc9cc08ebf72", x"ae72920a12ecd7f4", x"e74c65bbbb2c65ee", x"f4340b157d1a7a15", x"ded3d2646d12f3fe");
            when 20691376 => data <= (x"5c3ff7213dcd7b8f", x"bd56268e30d18a88", x"c6dd45d2691f98e0", x"51e30eedf415da68", x"9438ad72a353ba06", x"6653dd3a63d6a619", x"2dd3173f67ab3c62", x"82046ccb7c68413c");
            when 19758244 => data <= (x"4516e48f4001f025", x"6a8bacf681bfdec2", x"ae502d488fe49409", x"2a36e2fd9793eeda", x"d93acd3ea52222e6", x"21a76fb8f62fc81d", x"99b9328694c5e07a", x"91ba88525faae9bc");
            when 22207166 => data <= (x"6cf12f3c506242cd", x"5c74e619d9ba8ec1", x"2a0a263ed17a6fb3", x"f167228b16e30a69", x"f72d411710aa9e2f", x"6e52c8716330d9b3", x"409a75f9ac431df9", x"0fe0e0e190f3fdee");
            when 2956502 => data <= (x"890316e6f06a89c2", x"3ae3bacc293274dc", x"f62955d983a4dd19", x"73a7492fd8078867", x"2df84e2c810f4ed1", x"4071e930f1c8f291", x"56a59c3f3e0a6309", x"ad86340147d9ee4d");
            when 13668453 => data <= (x"7cc1f5adfdd46c9c", x"67975063449ce8ba", x"f7c8d1117265043e", x"fdb803b5f426b3a9", x"3f2dca5c22a65e48", x"4fd0f669837d94ee", x"3148f600b1cf6c18", x"6bbbc5f722f85b6f");
            when 27737809 => data <= (x"1edf06b2df6566a9", x"d74e0d846f8cf6ea", x"ffbd3a0a9d41fb90", x"28b5c1e2c5343aec", x"23b8d075fd4075e5", x"8451164636a82af2", x"d4b0d4ac4baf52ff", x"2ee8561e0452fdd1");
            when 11142824 => data <= (x"72ed8b9668e07d02", x"1378f0bb19ea12db", x"b79f44476a62facf", x"42ca8783f2ebc31c", x"30c8dfa0bef03bf6", x"b54234c7805ded69", x"4c15740faa7d0b18", x"a841dd6c1adc127a");
            when 21168767 => data <= (x"d3c45ea72594b226", x"657283dab7223945", x"8f39bb4aaf0e31e2", x"9649135c00e7e104", x"463017408387a461", x"52872a8c232fe0a8", x"b677b707301e1444", x"1fb308db287bc930");
            when 28114580 => data <= (x"8841ebfe3782a955", x"73e2a5bc334cd26e", x"ba5a6f7825582aff", x"4e6c3fc4085a360e", x"bc686d337fa88721", x"dc64468ebaba5df4", x"9c64fbba5c69c8c4", x"307771e0c0f4cd13");
            when 297382 => data <= (x"297dc5a29526ae83", x"ef997b6ffc623cc0", x"7f9f8d1cd1d4364c", x"bc60e97e0c94b162", x"89422306df51a815", x"f5bfb775fba24e79", x"f7bd025b5c6c352d", x"90dcf876d3f8147f");
            when 13603496 => data <= (x"d466e3fcea31626c", x"5a40921bbbd62911", x"6c7a7370b20cbd4c", x"5db3a626cd83b592", x"2e3df34ce5f8fd4b", x"5b12f5b3b419c644", x"03389beb0cae4e26", x"f3e9abfedc21a377");
            when 17929015 => data <= (x"5162d1e31876a1a0", x"dfed99fe36afcb80", x"1242053f34aedeff", x"600b9e138f8ebb9d", x"d512e134d8c81062", x"dc64a016fad10b86", x"902647c2a1b2b746", x"bd2c85ba92d3415e");
            when 24133818 => data <= (x"210c08ff1a64d55c", x"cf628915ac5f8af1", x"a286d77407816e71", x"13bd909f05ffd7aa", x"f80d7467dabd4d28", x"fa89448a9a4190c1", x"55e357a2f546b21f", x"aa124253b621a526");
            when 29141181 => data <= (x"6f1919908ee31c71", x"69a5aa8261cb3f4d", x"00a742440fb6435b", x"ed39e8e73bd5bed1", x"ca30c0657b0c8f63", x"f7d2b118db2adf13", x"cce6468dd63dfd4f", x"7296905a610a4483");
            when 4203934 => data <= (x"b12317aa34c25389", x"87df0e1f2f01806a", x"121fe5ce60b2dcd4", x"46cc329e4dea110f", x"7445d30417d46452", x"96c9583a75b7579e", x"a46a4d06eeb1ae52", x"6e69ded2d723fec0");
            when 16739833 => data <= (x"66b605de7ee1773e", x"e93abec965f0b820", x"976e0f231621f2b0", x"2e9550bc044697c7", x"484edd8628a53263", x"7fef081e4abfc368", x"4b877e5a1e91c9f9", x"8e2e95d2a3dd58aa");
            when 28084737 => data <= (x"23655f7320ab358b", x"5d48e24ea90142cb", x"4b9ab5ff5489ad0d", x"5254af1d24a22b37", x"6bf7f2b5b3c7442e", x"4c29f87dcdd35393", x"13270c7cf90e7c4e", x"db27fa165a83eecf");
            when 1240137 => data <= (x"aaed79478a1b9e29", x"63c81242df45ba92", x"a29d45298ada5e31", x"d2498574e1fc22ad", x"82c32f1b3c6aca41", x"8304d799f5929364", x"9b4ee5d203d3b5fb", x"f59aa2e02e205e2d");
            when 5165073 => data <= (x"059b535c3023341b", x"f8a4d22b5792a89b", x"00fb22055bf6ae52", x"35fb48dc10d3db14", x"cd7cee32b66d2f6c", x"9b5cbd04df760d93", x"e380fe4f51e79208", x"210d9e6d7d93955d");
            when 17120387 => data <= (x"1ba125378feef6bd", x"baaea155b78f77be", x"6bf26dc95d4b89b8", x"1dec1209562ff542", x"4f43a98f20f58f7b", x"4b8f376b2006270f", x"94036e8484a0a861", x"5efdb55a659d0c37");
            when 28712565 => data <= (x"661bc4f8c249a3ae", x"178e31b6e6dae1e6", x"023f5991d3c214ea", x"ddb4c4f7128d2fe8", x"e5203511a5832941", x"cfa0fe1a26b8c720", x"c5f64555822e18e5", x"e3d908e480afa032");
            when 3713103 => data <= (x"f251a330bf9e4d9f", x"b56e1aa06bc78251", x"b6c696ba82670742", x"554e9d5c037a9996", x"b3a495d6e8cef4db", x"d020894d213a2ec5", x"a75f128cad7aac07", x"68467727b46eba69");
            when 16673004 => data <= (x"0ff1de00277e1769", x"bd7662c1c4bfe7f7", x"5e1c4062f0712273", x"a259fd812a5f3038", x"68768b68bb63d3e3", x"9a4a9689a29e95c1", x"ef1dacce2660c7a2", x"ac46ae19e615baac");
            when 25059055 => data <= (x"7b7c17c52a889e2a", x"3b11bf0a81734264", x"96ffd13308beb279", x"73dda737ca66adc5", x"b651e9b60978e9ce", x"6eac089e766227ed", x"832daba1c699f7da", x"47eec58cd41518e5");
            when 24722983 => data <= (x"76b55ddeb5a936c4", x"cda8e32375b7d017", x"9a35f5b278a6b1af", x"e843e10356cc1786", x"a558ebf26c9b4a29", x"5b0811d770a84c5e", x"9d40c24b6fe7a4e3", x"bacd254fd32b66f8");
            when 18924519 => data <= (x"761611b303ece734", x"32f7b964662a0415", x"64a0270ea7030d99", x"5c32e1e89722618c", x"56a38c6c3154771a", x"dae6441aeca237f8", x"a57ff0f8343eb0bd", x"9dc6fcb2cf78035c");
            when 33766630 => data <= (x"962c622c55687801", x"382a06cd3c27b345", x"134bde1aca78e19b", x"edaa9c4954b8e120", x"581ff1e44892b0a9", x"f78300e0a67493dd", x"476f73b653af2fdb", x"5abf5c15dfa7a078");
            when 8381887 => data <= (x"c0d4086cb157dfa5", x"7200f6bfd1f96325", x"0044af530f7227e5", x"41df3f406c1a500f", x"2b6d14bcba3c9c34", x"947a1ebee3a37d0c", x"69054a3b3853534b", x"1e22d4d184b34d3d");
            when 5721477 => data <= (x"5d51c2746f6aa0ec", x"6c68b48ae215366d", x"64f7bd67c8871974", x"df5cd2d1f7e7ddc1", x"4f434e1eb154b0e9", x"380401cf4482f5c8", x"7d29c95114c58659", x"fd76d808899fc79c");
            when 18678087 => data <= (x"8186b4d233a81f0f", x"7b837080720bedaf", x"8989fd0832c16840", x"67932eb20fe5500e", x"0228d955aaa9ddb7", x"c40573780094fc08", x"63fa4dbf3fd9286d", x"4186ea75572f1326");
            when 25779616 => data <= (x"b295516456a32036", x"97964d19f252a180", x"c353acde0d878125", x"d792b1179ddbda90", x"b41d8162a5e942d8", x"903a0970203946c5", x"bf9fb2a2931a1a77", x"e97bc7b25f068be1");
            when 13974985 => data <= (x"29912cfd6c18462f", x"0964dd13d7e97d52", x"9217d9fedbd475ef", x"60b1f6f633077d01", x"00fd09c8ea56aa22", x"f0732136162e26d7", x"1e652cc5cd4d5d19", x"679947521425a0e0");
            when 14798958 => data <= (x"859c131d78c137db", x"a3c9ef38d5b1b45b", x"840b5ae668d9b427", x"6bf53b3bbc523a91", x"6e7656a33e7f8491", x"13996fc325a88252", x"11da089c6a5c78d1", x"28c4f52e6372f974");
            when 12415666 => data <= (x"d8092cd4af16cb50", x"1485a05a4317a8c4", x"42c340736b52200f", x"83be2b3e9868baf5", x"7a968b266099d9ea", x"782b50b812016b37", x"d1f2ccee4a561c6d", x"e2b78320782bd751");
            when 33562258 => data <= (x"efbe66acdb78dbd9", x"42ae0f8dcbfdedbb", x"58053db05e889789", x"bc0849c5964c8918", x"8116cf4ca644c0d5", x"5a9f7c03786bab22", x"2369c983fd4f6d0c", x"e096430ee88e9d92");
            when 20519770 => data <= (x"0f3e7b02623cdf2b", x"19365cb0f35b7e4c", x"45adabb994d8a26d", x"004bbda92a948015", x"2b61bfcbe8c02978", x"9af9234701e9b5de", x"44e0636c585ae638", x"192439d1e6a180f5");
            when 11917666 => data <= (x"6a19c6e1e632b5ef", x"786d84ad61ea6095", x"bd4d79fbd9c43fc4", x"653b090551daaaab", x"ea1d4e1b3aecca1d", x"546c09ad11c3647d", x"b6084255b46c372c", x"03843db28c1100e2");
            when 3440569 => data <= (x"68c36a3b67aa36d4", x"b3698f0b1780510d", x"441a700b9339bb1d", x"d5ef4cd990ec534d", x"c89e2ad400f6aeb7", x"3c2441831629007d", x"132dc773dc3dc1f3", x"07823b695f38e4c1");
            when 32962438 => data <= (x"07ef5b9b2b4feb2e", x"42344f63a4de2024", x"9dfb0fdd69daf3c6", x"ad7085d9932d8aec", x"7e5efa882af160a0", x"b5d368a0a855eac9", x"6ae166f7f6bcfdb2", x"7ac06d10ece65c5e");
            when 23914225 => data <= (x"ff5d440aa1b83774", x"a896808fb656f034", x"4a6781f52821b670", x"76a2886452bbe8e5", x"b9741f9aa442f076", x"3915a20a82a5a942", x"51c89fac3e7d6002", x"ebfee3752c0aa808");
            when 32524318 => data <= (x"86b07123c4065f1e", x"002099c0d155c135", x"18f1e535067c32cc", x"1513fcbd13493d03", x"eb36f0737f6844b3", x"64759db91b12b04e", x"89543e0d2a3b4e4c", x"a05a428deb86832b");
            when 4859099 => data <= (x"473fe2fe443d0286", x"105e58b5906d7f4f", x"e2af76930bacf22d", x"ab211d2178c62096", x"31c8db9a9853ffe7", x"722b23af9f71a35d", x"921f5a1c0cf6d6cd", x"ddbb02d4dc7a59e7");
            when 25675445 => data <= (x"195a782a407033a7", x"fce4b9c74b1cc846", x"cc8584fbbc4e4e30", x"a566b835f1d20b27", x"5db3f087b104ed8f", x"b73a6f72d30dd64c", x"c6bc0e77e7589927", x"bd063b28dd48fbb7");
            when 33247937 => data <= (x"90e6514592feee29", x"be893800d92cea4c", x"20fecbef722ddaaa", x"a9ccc34641c25002", x"f549869f219292e3", x"4083aeb25f1916cf", x"2c816f101e6dd78b", x"594a14c679acff91");
            when 10016582 => data <= (x"189e257bf9c34a4f", x"21e74e88509f8bd0", x"8c875fdcdcbe669a", x"55c9e7a8fd2469f8", x"1bd5f6131f450dbb", x"1d4f62bbf73ccd88", x"ee2d2d4b8de5b29a", x"2fbcfc71ddaac44a");
            when 14055595 => data <= (x"3ef6b9534f8006e8", x"858aa363a59aaa1b", x"3490c7d946c12484", x"4e941d8afe68191a", x"d0397e6cdd7169d9", x"1a2be21c7dfc4b2c", x"f460fa96f568fa7b", x"f3b6b7bdf8efa25a");
            when 2020156 => data <= (x"846881ddc080642c", x"91d0ccb59e647cf0", x"2ecc1d6dad0b7e52", x"f826b631c9c12cf2", x"e6453677f4287a87", x"2fb7ceae441d674a", x"a35f26b2d96d4f25", x"e175a8e114f1a0eb");
            when 30030505 => data <= (x"e77c8005fd922c89", x"4d1e7c3c6ecf590e", x"2bff68c69b19f045", x"6d2ddde150ca2be5", x"afd070f02173ff87", x"328ee21058e08c81", x"b1698223ffd6706e", x"90afb90c1a17efde");
            when 8617169 => data <= (x"26c7b819a1f1f1be", x"469b39798676faee", x"97aa83db03f746b6", x"fa7423188451a782", x"85b2b830dc79984d", x"f16784a252375a21", x"d18e2f7d2606f685", x"82e9026a0df86b94");
            when 31377517 => data <= (x"96e3fe483ba65deb", x"0c418fff32061fcc", x"0f5c68633ad689f7", x"fb58cd9281810d1f", x"2a73423753658ef4", x"60eaa0be9c923899", x"3c238454910c4114", x"2d01291806143400");
            when 27946321 => data <= (x"cca87319c24cfc2b", x"7a62944deb8a74cf", x"607c89558009e276", x"8fd0f13118ebc157", x"5343341ac94070dd", x"63e17721be55573b", x"4ad599ff3c28664a", x"671e058963eee71d");
            when 407792 => data <= (x"5a52e4e5114cd05f", x"9a8d95a5f351aa67", x"5c311e49be8bc0b3", x"b07991e545e605f6", x"8cd64e1ede9170c4", x"a78c7eb44eb3fd3c", x"a0720d1702e9bb7a", x"548100a1b04ede85");
            when 26579151 => data <= (x"c28023e743387896", x"28a0dfb9bedc0f0e", x"5c35a973047c4f66", x"8f850c814ba6df9c", x"b360f2b4673390b0", x"2dd493d91cf6525d", x"48c3077fd52be9d5", x"bc3055c41f7a44eb");
            when 32475890 => data <= (x"4c20b9c882b967b3", x"bcd4e2b25a6cb19c", x"a408b6e69a732d4f", x"84a5092f169222bc", x"f565c1bdebe0df9d", x"6d85dd9fd5d4041f", x"74753aa31c45d1e4", x"f8eb278f88094dcf");
            when 2296847 => data <= (x"6ae9b14f9c2b014a", x"79e45e98ef457e9f", x"76ee9117a99ed8ee", x"d77669a583161690", x"1396605ac991fa90", x"8f44c29250cf7df2", x"c68263d881e4b0be", x"c43f09148ca10c11");
            when 20556989 => data <= (x"ec962a5b012e55a0", x"766d62a9ef764183", x"6e512749b9873d88", x"4394e3f70828f884", x"826b820ba6565b93", x"dbba53e861080c7d", x"ec754aadbde9ff8c", x"61225199e88ffcc6");
            when 13748254 => data <= (x"d94bac44adbe90aa", x"d8f464c3fa2b6458", x"789aab0702b8c499", x"e558b14ab6ae83c2", x"b4fbc0cea78912d0", x"4a02856bcf9002a7", x"4066359aac0d1464", x"fc323bda23dceca6");
            when 24263142 => data <= (x"f3bb04c53c35409c", x"8603231b2c9101fa", x"eea0d50d345d8dc7", x"701e72e1e4430947", x"d9057ed5b1d1b6ba", x"db815f65d0512a7d", x"a820e2a52a64fc91", x"68757e6d9a56c54e");
            when 27657692 => data <= (x"874292af6e6ba4ad", x"07edd1db7e01a089", x"f3a76d4ea2e1b267", x"079c22f375722c6a", x"5f55a089a24d504c", x"091d5168c193704d", x"b909968a09d046eb", x"c87211be2bfb020e");
            when 29611312 => data <= (x"00e91e211e599c92", x"0074798ddb2a7cd3", x"89fc01ec0968a9e9", x"1cc1cc55086c5881", x"fb447fd53a034cce", x"242c97c2d254b3bd", x"93ef94fcf664625a", x"d8755a136c401342");
            when 20935452 => data <= (x"68fe20939f53b1e5", x"ad1b6e7a826ba89c", x"32069d1126f08f68", x"5a3c37c046091582", x"69aba2bbe460d4fd", x"26f289b98423e963", x"f4af7b6769ca2ca7", x"97645f0140dc830e");
            when 27675905 => data <= (x"f270ebd198804007", x"1fa1cb46a7098b7b", x"d0db85aa1005332e", x"e5b681739ec08fe0", x"e4d247cd16dff172", x"f48fd165e4bb1fed", x"37d9717b3cd9f744", x"73abf21870f54ced");
            when 10683825 => data <= (x"a3eb13ec00fc333a", x"75dad2fc0061ad92", x"b538ca629226a9c8", x"d0f8c5a78d10b3cb", x"811a028b19c0f6b8", x"aabe3b1185b89cbf", x"316e5c164452af78", x"019af27886052cd4");
            when 15777353 => data <= (x"1508309f4ae92f0f", x"6893e5e9b89b46ce", x"315fa203acee7f54", x"bb0aae8663eeebe6", x"0a5201d8bfa43f8b", x"08af10c5c37033bd", x"a43b7065ebdf5d25", x"dd1cfbda4f0db4ac");
            when 27512872 => data <= (x"ff580d257647ce22", x"a58f35fb79695083", x"85c501d830146a33", x"09c9b13b1bba2506", x"743ec7cd74903d47", x"158b390ac53012bf", x"911ee00c9dd1a8cd", x"17fd9ce5edf1931d"); 
            when others => data <= (others => (others => '0'));
        end case;

    end process;

end behavioral;