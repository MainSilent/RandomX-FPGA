library ieee;
use ieee.std_logic_1164.all;


package aes_sbox is

    function lutEnc0 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector;

    function lutEnc1 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector;

    function lutEnc2 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector;

    function lutEnc3 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector;

    function lutDec0 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector;

    function lutDec1 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector;

    function lutDec2 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector;

    function lutDec3 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector;

end package;


package body aes_sbox is
    
    ------------------------------ ENC ------------------------------

    function lutEnc0 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector is variable output : std_logic_vector(31 downto 0);
    begin
		case input is
            when x"00" => output := x"a56363c6";
            when x"01" => output := x"847c7cf8";
            when x"02" => output := x"997777ee";
            when x"03" => output := x"8d7b7bf6";
            when x"04" => output := x"0df2f2ff";
            when x"05" => output := x"bd6b6bd6";
            when x"06" => output := x"b16f6fde";
            when x"07" => output := x"54c5c591";
            when x"08" => output := x"50303060";
            when x"09" => output := x"03010102";
            when x"0a" => output := x"a96767ce";
            when x"0b" => output := x"7d2b2b56";
            when x"0c" => output := x"19fefee7";
            when x"0d" => output := x"62d7d7b5";
            when x"0e" => output := x"e6abab4d";
            when x"0f" => output := x"9a7676ec";
            when x"10" => output := x"45caca8f";
            when x"11" => output := x"9d82821f";
            when x"12" => output := x"40c9c989";
            when x"13" => output := x"877d7dfa";
            when x"14" => output := x"15fafaef";
            when x"15" => output := x"eb5959b2";
            when x"16" => output := x"c947478e";
            when x"17" => output := x"0bf0f0fb";
            when x"18" => output := x"ecadad41";
            when x"19" => output := x"67d4d4b3";
            when x"1a" => output := x"fda2a25f";
            when x"1b" => output := x"eaafaf45";
            when x"1c" => output := x"bf9c9c23";
            when x"1d" => output := x"f7a4a453";
            when x"1e" => output := x"967272e4";
            when x"1f" => output := x"5bc0c09b";
            when x"20" => output := x"c2b7b775";
            when x"21" => output := x"1cfdfde1";
            when x"22" => output := x"ae93933d";
            when x"23" => output := x"6a26264c";
            when x"24" => output := x"5a36366c";
            when x"25" => output := x"413f3f7e";
            when x"26" => output := x"02f7f7f5";
            when x"27" => output := x"4fcccc83";
            when x"28" => output := x"5c343468";
            when x"29" => output := x"f4a5a551";
            when x"2a" => output := x"34e5e5d1";
            when x"2b" => output := x"08f1f1f9";
            when x"2c" => output := x"937171e2";
            when x"2d" => output := x"73d8d8ab";
            when x"2e" => output := x"53313162";
            when x"2f" => output := x"3f15152a";
            when x"30" => output := x"0c040408";
            when x"31" => output := x"52c7c795";
            when x"32" => output := x"65232346";
            when x"33" => output := x"5ec3c39d";
            when x"34" => output := x"28181830";
            when x"35" => output := x"a1969637";
            when x"36" => output := x"0f05050a";
            when x"37" => output := x"b59a9a2f";
            when x"38" => output := x"0907070e";
            when x"39" => output := x"36121224";
            when x"3a" => output := x"9b80801b";
            when x"3b" => output := x"3de2e2df";
            when x"3c" => output := x"26ebebcd";
            when x"3d" => output := x"6927274e";
            when x"3e" => output := x"cdb2b27f";
            when x"3f" => output := x"9f7575ea";
            when x"40" => output := x"1b090912";
            when x"41" => output := x"9e83831d";
            when x"42" => output := x"742c2c58";
            when x"43" => output := x"2e1a1a34";
            when x"44" => output := x"2d1b1b36";
            when x"45" => output := x"b26e6edc";
            when x"46" => output := x"ee5a5ab4";
            when x"47" => output := x"fba0a05b";
            when x"48" => output := x"f65252a4";
            when x"49" => output := x"4d3b3b76";
            when x"4a" => output := x"61d6d6b7";
            when x"4b" => output := x"ceb3b37d";
            when x"4c" => output := x"7b292952";
            when x"4d" => output := x"3ee3e3dd";
            when x"4e" => output := x"712f2f5e";
            when x"4f" => output := x"97848413";
            when x"50" => output := x"f55353a6";
            when x"51" => output := x"68d1d1b9";
            when x"52" => output := x"00000000";
            when x"53" => output := x"2cededc1";
            when x"54" => output := x"60202040";
            when x"55" => output := x"1ffcfce3";
            when x"56" => output := x"c8b1b179";
            when x"57" => output := x"ed5b5bb6";
            when x"58" => output := x"be6a6ad4";
            when x"59" => output := x"46cbcb8d";
            when x"5a" => output := x"d9bebe67";
            when x"5b" => output := x"4b393972";
            when x"5c" => output := x"de4a4a94";
            when x"5d" => output := x"d44c4c98";
            when x"5e" => output := x"e85858b0";
            when x"5f" => output := x"4acfcf85";
            when x"60" => output := x"6bd0d0bb";
            when x"61" => output := x"2aefefc5";
            when x"62" => output := x"e5aaaa4f";
            when x"63" => output := x"16fbfbed";
            when x"64" => output := x"c5434386";
            when x"65" => output := x"d74d4d9a";
            when x"66" => output := x"55333366";
            when x"67" => output := x"94858511";
            when x"68" => output := x"cf45458a";
            when x"69" => output := x"10f9f9e9";
            when x"6a" => output := x"06020204";
            when x"6b" => output := x"817f7ffe";
            when x"6c" => output := x"f05050a0";
            when x"6d" => output := x"443c3c78";
            when x"6e" => output := x"ba9f9f25";
            when x"6f" => output := x"e3a8a84b";
            when x"70" => output := x"f35151a2";
            when x"71" => output := x"fea3a35d";
            when x"72" => output := x"c0404080";
            when x"73" => output := x"8a8f8f05";
            when x"74" => output := x"ad92923f";
            when x"75" => output := x"bc9d9d21";
            when x"76" => output := x"48383870";
            when x"77" => output := x"04f5f5f1";
            when x"78" => output := x"dfbcbc63";
            when x"79" => output := x"c1b6b677";
            when x"7a" => output := x"75dadaaf";
            when x"7b" => output := x"63212142";
            when x"7c" => output := x"30101020";
            when x"7d" => output := x"1affffe5";
            when x"7e" => output := x"0ef3f3fd";
            when x"7f" => output := x"6dd2d2bf";
            when x"80" => output := x"4ccdcd81";
            when x"81" => output := x"140c0c18";
            when x"82" => output := x"35131326";
            when x"83" => output := x"2fececc3";
            when x"84" => output := x"e15f5fbe";
            when x"85" => output := x"a2979735";
            when x"86" => output := x"cc444488";
            when x"87" => output := x"3917172e";
            when x"88" => output := x"57c4c493";
            when x"89" => output := x"f2a7a755";
            when x"8a" => output := x"827e7efc";
            when x"8b" => output := x"473d3d7a";
            when x"8c" => output := x"ac6464c8";
            when x"8d" => output := x"e75d5dba";
            when x"8e" => output := x"2b191932";
            when x"8f" => output := x"957373e6";
            when x"90" => output := x"a06060c0";
            when x"91" => output := x"98818119";
            when x"92" => output := x"d14f4f9e";
            when x"93" => output := x"7fdcdca3";
            when x"94" => output := x"66222244";
            when x"95" => output := x"7e2a2a54";
            when x"96" => output := x"ab90903b";
            when x"97" => output := x"8388880b";
            when x"98" => output := x"ca46468c";
            when x"99" => output := x"29eeeec7";
            when x"9a" => output := x"d3b8b86b";
            when x"9b" => output := x"3c141428";
            when x"9c" => output := x"79dedea7";
            when x"9d" => output := x"e25e5ebc";
            when x"9e" => output := x"1d0b0b16";
            when x"9f" => output := x"76dbdbad";
            when x"a0" => output := x"3be0e0db";
            when x"a1" => output := x"56323264";
            when x"a2" => output := x"4e3a3a74";
            when x"a3" => output := x"1e0a0a14";
            when x"a4" => output := x"db494992";
            when x"a5" => output := x"0a06060c";
            when x"a6" => output := x"6c242448";
            when x"a7" => output := x"e45c5cb8";
            when x"a8" => output := x"5dc2c29f";
            when x"a9" => output := x"6ed3d3bd";
            when x"aa" => output := x"efacac43";
            when x"ab" => output := x"a66262c4";
            when x"ac" => output := x"a8919139";
            when x"ad" => output := x"a4959531";
            when x"ae" => output := x"37e4e4d3";
            when x"af" => output := x"8b7979f2";
            when x"b0" => output := x"32e7e7d5";
            when x"b1" => output := x"43c8c88b";
            when x"b2" => output := x"5937376e";
            when x"b3" => output := x"b76d6dda";
            when x"b4" => output := x"8c8d8d01";
            when x"b5" => output := x"64d5d5b1";
            when x"b6" => output := x"d24e4e9c";
            when x"b7" => output := x"e0a9a949";
            when x"b8" => output := x"b46c6cd8";
            when x"b9" => output := x"fa5656ac";
            when x"ba" => output := x"07f4f4f3";
            when x"bb" => output := x"25eaeacf";
            when x"bc" => output := x"af6565ca";
            when x"bd" => output := x"8e7a7af4";
            when x"be" => output := x"e9aeae47";
            when x"bf" => output := x"18080810";
            when x"c0" => output := x"d5baba6f";
            when x"c1" => output := x"887878f0";
            when x"c2" => output := x"6f25254a";
            when x"c3" => output := x"722e2e5c";
            when x"c4" => output := x"241c1c38";
            when x"c5" => output := x"f1a6a657";
            when x"c6" => output := x"c7b4b473";
            when x"c7" => output := x"51c6c697";
            when x"c8" => output := x"23e8e8cb";
            when x"c9" => output := x"7cdddda1";
            when x"ca" => output := x"9c7474e8";
            when x"cb" => output := x"211f1f3e";
            when x"cc" => output := x"dd4b4b96";
            when x"cd" => output := x"dcbdbd61";
            when x"ce" => output := x"868b8b0d";
            when x"cf" => output := x"858a8a0f";
            when x"d0" => output := x"907070e0";
            when x"d1" => output := x"423e3e7c";
            when x"d2" => output := x"c4b5b571";
            when x"d3" => output := x"aa6666cc";
            when x"d4" => output := x"d8484890";
            when x"d5" => output := x"05030306";
            when x"d6" => output := x"01f6f6f7";
            when x"d7" => output := x"120e0e1c";
            when x"d8" => output := x"a36161c2";
            when x"d9" => output := x"5f35356a";
            when x"da" => output := x"f95757ae";
            when x"db" => output := x"d0b9b969";
            when x"dc" => output := x"91868617";
            when x"dd" => output := x"58c1c199";
            when x"de" => output := x"271d1d3a";
            when x"df" => output := x"b99e9e27";
            when x"e0" => output := x"38e1e1d9";
            when x"e1" => output := x"13f8f8eb";
            when x"e2" => output := x"b398982b";
            when x"e3" => output := x"33111122";
            when x"e4" => output := x"bb6969d2";
            when x"e5" => output := x"70d9d9a9";
            when x"e6" => output := x"898e8e07";
            when x"e7" => output := x"a7949433";
            when x"e8" => output := x"b69b9b2d";
            when x"e9" => output := x"221e1e3c";
            when x"ea" => output := x"92878715";
            when x"eb" => output := x"20e9e9c9";
            when x"ec" => output := x"49cece87";
            when x"ed" => output := x"ff5555aa";
            when x"ee" => output := x"78282850";
            when x"ef" => output := x"7adfdfa5";
            when x"f0" => output := x"8f8c8c03";
            when x"f1" => output := x"f8a1a159";
            when x"f2" => output := x"80898909";
            when x"f3" => output := x"170d0d1a";
            when x"f4" => output := x"dabfbf65";
            when x"f5" => output := x"31e6e6d7";
            when x"f6" => output := x"c6424284";
            when x"f7" => output := x"b86868d0";
            when x"f8" => output := x"c3414182";
            when x"f9" => output := x"b0999929";
            when x"fa" => output := x"772d2d5a";
            when x"fb" => output := x"110f0f1e";
            when x"fc" => output := x"cbb0b07b";
            when x"fd" => output := x"fc5454a8";
            when x"fe" => output := x"d6bbbb6d";
            when x"ff" => output := x"3a16162c";
			when others => null;
		end case;

        return output;
    end;

    function lutEnc1 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector is variable output : std_logic_vector(31 downto 0);
    begin
        case input is
            when x"00" => output := x"6363c6a5";
            when x"01" => output := x"7c7cf884";
            when x"02" => output := x"7777ee99";
            when x"03" => output := x"7b7bf68d";
            when x"04" => output := x"f2f2ff0d";
            when x"05" => output := x"6b6bd6bd";
            when x"06" => output := x"6f6fdeb1";
            when x"07" => output := x"c5c59154";
            when x"08" => output := x"30306050";
            when x"09" => output := x"01010203";
            when x"0a" => output := x"6767cea9";
            when x"0b" => output := x"2b2b567d";
            when x"0c" => output := x"fefee719";
            when x"0d" => output := x"d7d7b562";
            when x"0e" => output := x"abab4de6";
            when x"0f" => output := x"7676ec9a";
            when x"10" => output := x"caca8f45";
            when x"11" => output := x"82821f9d";
            when x"12" => output := x"c9c98940";
            when x"13" => output := x"7d7dfa87";
            when x"14" => output := x"fafaef15";
            when x"15" => output := x"5959b2eb";
            when x"16" => output := x"47478ec9";
            when x"17" => output := x"f0f0fb0b";
            when x"18" => output := x"adad41ec";
            when x"19" => output := x"d4d4b367";
            when x"1a" => output := x"a2a25ffd";
            when x"1b" => output := x"afaf45ea";
            when x"1c" => output := x"9c9c23bf";
            when x"1d" => output := x"a4a453f7";
            when x"1e" => output := x"7272e496";
            when x"1f" => output := x"c0c09b5b";
            when x"20" => output := x"b7b775c2";
            when x"21" => output := x"fdfde11c";
            when x"22" => output := x"93933dae";
            when x"23" => output := x"26264c6a";
            when x"24" => output := x"36366c5a";
            when x"25" => output := x"3f3f7e41";
            when x"26" => output := x"f7f7f502";
            when x"27" => output := x"cccc834f";
            when x"28" => output := x"3434685c";
            when x"29" => output := x"a5a551f4";
            when x"2a" => output := x"e5e5d134";
            when x"2b" => output := x"f1f1f908";
            when x"2c" => output := x"7171e293";
            when x"2d" => output := x"d8d8ab73";
            when x"2e" => output := x"31316253";
            when x"2f" => output := x"15152a3f";
            when x"30" => output := x"0404080c";
            when x"31" => output := x"c7c79552";
            when x"32" => output := x"23234665";
            when x"33" => output := x"c3c39d5e";
            when x"34" => output := x"18183028";
            when x"35" => output := x"969637a1";
            when x"36" => output := x"05050a0f";
            when x"37" => output := x"9a9a2fb5";
            when x"38" => output := x"07070e09";
            when x"39" => output := x"12122436";
            when x"3a" => output := x"80801b9b";
            when x"3b" => output := x"e2e2df3d";
            when x"3c" => output := x"ebebcd26";
            when x"3d" => output := x"27274e69";
            when x"3e" => output := x"b2b27fcd";
            when x"3f" => output := x"7575ea9f";
            when x"40" => output := x"0909121b";
            when x"41" => output := x"83831d9e";
            when x"42" => output := x"2c2c5874";
            when x"43" => output := x"1a1a342e";
            when x"44" => output := x"1b1b362d";
            when x"45" => output := x"6e6edcb2";
            when x"46" => output := x"5a5ab4ee";
            when x"47" => output := x"a0a05bfb";
            when x"48" => output := x"5252a4f6";
            when x"49" => output := x"3b3b764d";
            when x"4a" => output := x"d6d6b761";
            when x"4b" => output := x"b3b37dce";
            when x"4c" => output := x"2929527b";
            when x"4d" => output := x"e3e3dd3e";
            when x"4e" => output := x"2f2f5e71";
            when x"4f" => output := x"84841397";
            when x"50" => output := x"5353a6f5";
            when x"51" => output := x"d1d1b968";
            when x"52" => output := x"00000000";
            when x"53" => output := x"ededc12c";
            when x"54" => output := x"20204060";
            when x"55" => output := x"fcfce31f";
            when x"56" => output := x"b1b179c8";
            when x"57" => output := x"5b5bb6ed";
            when x"58" => output := x"6a6ad4be";
            when x"59" => output := x"cbcb8d46";
            when x"5a" => output := x"bebe67d9";
            when x"5b" => output := x"3939724b";
            when x"5c" => output := x"4a4a94de";
            when x"5d" => output := x"4c4c98d4";
            when x"5e" => output := x"5858b0e8";
            when x"5f" => output := x"cfcf854a";
            when x"60" => output := x"d0d0bb6b";
            when x"61" => output := x"efefc52a";
            when x"62" => output := x"aaaa4fe5";
            when x"63" => output := x"fbfbed16";
            when x"64" => output := x"434386c5";
            when x"65" => output := x"4d4d9ad7";
            when x"66" => output := x"33336655";
            when x"67" => output := x"85851194";
            when x"68" => output := x"45458acf";
            when x"69" => output := x"f9f9e910";
            when x"6a" => output := x"02020406";
            when x"6b" => output := x"7f7ffe81";
            when x"6c" => output := x"5050a0f0";
            when x"6d" => output := x"3c3c7844";
            when x"6e" => output := x"9f9f25ba";
            when x"6f" => output := x"a8a84be3";
            when x"70" => output := x"5151a2f3";
            when x"71" => output := x"a3a35dfe";
            when x"72" => output := x"404080c0";
            when x"73" => output := x"8f8f058a";
            when x"74" => output := x"92923fad";
            when x"75" => output := x"9d9d21bc";
            when x"76" => output := x"38387048";
            when x"77" => output := x"f5f5f104";
            when x"78" => output := x"bcbc63df";
            when x"79" => output := x"b6b677c1";
            when x"7a" => output := x"dadaaf75";
            when x"7b" => output := x"21214263";
            when x"7c" => output := x"10102030";
            when x"7d" => output := x"ffffe51a";
            when x"7e" => output := x"f3f3fd0e";
            when x"7f" => output := x"d2d2bf6d";
            when x"80" => output := x"cdcd814c";
            when x"81" => output := x"0c0c1814";
            when x"82" => output := x"13132635";
            when x"83" => output := x"ececc32f";
            when x"84" => output := x"5f5fbee1";
            when x"85" => output := x"979735a2";
            when x"86" => output := x"444488cc";
            when x"87" => output := x"17172e39";
            when x"88" => output := x"c4c49357";
            when x"89" => output := x"a7a755f2";
            when x"8a" => output := x"7e7efc82";
            when x"8b" => output := x"3d3d7a47";
            when x"8c" => output := x"6464c8ac";
            when x"8d" => output := x"5d5dbae7";
            when x"8e" => output := x"1919322b";
            when x"8f" => output := x"7373e695";
            when x"90" => output := x"6060c0a0";
            when x"91" => output := x"81811998";
            when x"92" => output := x"4f4f9ed1";
            when x"93" => output := x"dcdca37f";
            when x"94" => output := x"22224466";
            when x"95" => output := x"2a2a547e";
            when x"96" => output := x"90903bab";
            when x"97" => output := x"88880b83";
            when x"98" => output := x"46468cca";
            when x"99" => output := x"eeeec729";
            when x"9a" => output := x"b8b86bd3";
            when x"9b" => output := x"1414283c";
            when x"9c" => output := x"dedea779";
            when x"9d" => output := x"5e5ebce2";
            when x"9e" => output := x"0b0b161d";
            when x"9f" => output := x"dbdbad76";
            when x"a0" => output := x"e0e0db3b";
            when x"a1" => output := x"32326456";
            when x"a2" => output := x"3a3a744e";
            when x"a3" => output := x"0a0a141e";
            when x"a4" => output := x"494992db";
            when x"a5" => output := x"06060c0a";
            when x"a6" => output := x"2424486c";
            when x"a7" => output := x"5c5cb8e4";
            when x"a8" => output := x"c2c29f5d";
            when x"a9" => output := x"d3d3bd6e";
            when x"aa" => output := x"acac43ef";
            when x"ab" => output := x"6262c4a6";
            when x"ac" => output := x"919139a8";
            when x"ad" => output := x"959531a4";
            when x"ae" => output := x"e4e4d337";
            when x"af" => output := x"7979f28b";
            when x"b0" => output := x"e7e7d532";
            when x"b1" => output := x"c8c88b43";
            when x"b2" => output := x"37376e59";
            when x"b3" => output := x"6d6ddab7";
            when x"b4" => output := x"8d8d018c";
            when x"b5" => output := x"d5d5b164";
            when x"b6" => output := x"4e4e9cd2";
            when x"b7" => output := x"a9a949e0";
            when x"b8" => output := x"6c6cd8b4";
            when x"b9" => output := x"5656acfa";
            when x"ba" => output := x"f4f4f307";
            when x"bb" => output := x"eaeacf25";
            when x"bc" => output := x"6565caaf";
            when x"bd" => output := x"7a7af48e";
            when x"be" => output := x"aeae47e9";
            when x"bf" => output := x"08081018";
            when x"c0" => output := x"baba6fd5";
            when x"c1" => output := x"7878f088";
            when x"c2" => output := x"25254a6f";
            when x"c3" => output := x"2e2e5c72";
            when x"c4" => output := x"1c1c3824";
            when x"c5" => output := x"a6a657f1";
            when x"c6" => output := x"b4b473c7";
            when x"c7" => output := x"c6c69751";
            when x"c8" => output := x"e8e8cb23";
            when x"c9" => output := x"dddda17c";
            when x"ca" => output := x"7474e89c";
            when x"cb" => output := x"1f1f3e21";
            when x"cc" => output := x"4b4b96dd";
            when x"cd" => output := x"bdbd61dc";
            when x"ce" => output := x"8b8b0d86";
            when x"cf" => output := x"8a8a0f85";
            when x"d0" => output := x"7070e090";
            when x"d1" => output := x"3e3e7c42";
            when x"d2" => output := x"b5b571c4";
            when x"d3" => output := x"6666ccaa";
            when x"d4" => output := x"484890d8";
            when x"d5" => output := x"03030605";
            when x"d6" => output := x"f6f6f701";
            when x"d7" => output := x"0e0e1c12";
            when x"d8" => output := x"6161c2a3";
            when x"d9" => output := x"35356a5f";
            when x"da" => output := x"5757aef9";
            when x"db" => output := x"b9b969d0";
            when x"dc" => output := x"86861791";
            when x"dd" => output := x"c1c19958";
            when x"de" => output := x"1d1d3a27";
            when x"df" => output := x"9e9e27b9";
            when x"e0" => output := x"e1e1d938";
            when x"e1" => output := x"f8f8eb13";
            when x"e2" => output := x"98982bb3";
            when x"e3" => output := x"11112233";
            when x"e4" => output := x"6969d2bb";
            when x"e5" => output := x"d9d9a970";
            when x"e6" => output := x"8e8e0789";
            when x"e7" => output := x"949433a7";
            when x"e8" => output := x"9b9b2db6";
            when x"e9" => output := x"1e1e3c22";
            when x"ea" => output := x"87871592";
            when x"eb" => output := x"e9e9c920";
            when x"ec" => output := x"cece8749";
            when x"ed" => output := x"5555aaff";
            when x"ee" => output := x"28285078";
            when x"ef" => output := x"dfdfa57a";
            when x"f0" => output := x"8c8c038f";
            when x"f1" => output := x"a1a159f8";
            when x"f2" => output := x"89890980";
            when x"f3" => output := x"0d0d1a17";
            when x"f4" => output := x"bfbf65da";
            when x"f5" => output := x"e6e6d731";
            when x"f6" => output := x"424284c6";
            when x"f7" => output := x"6868d0b8";
            when x"f8" => output := x"414182c3";
            when x"f9" => output := x"999929b0";
            when x"fa" => output := x"2d2d5a77";
            when x"fb" => output := x"0f0f1e11";
            when x"fc" => output := x"b0b07bcb";
            when x"fd" => output := x"5454a8fc";
            when x"fe" => output := x"bbbb6dd6";
            when x"ff" => output := x"16162c3a";
            when others => null;
        end case;

        return output;
    end;

    function lutEnc2 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector is variable output : std_logic_vector(31 downto 0);
    begin
        case input is
            when x"00" => output := x"63c6a563";
            when x"01" => output := x"7cf8847c";
            when x"02" => output := x"77ee9977";
            when x"03" => output := x"7bf68d7b";
            when x"04" => output := x"f2ff0df2";
            when x"05" => output := x"6bd6bd6b";
            when x"06" => output := x"6fdeb16f";
            when x"07" => output := x"c59154c5";
            when x"08" => output := x"30605030";
            when x"09" => output := x"01020301";
            when x"0a" => output := x"67cea967";
            when x"0b" => output := x"2b567d2b";
            when x"0c" => output := x"fee719fe";
            when x"0d" => output := x"d7b562d7";
            when x"0e" => output := x"ab4de6ab";
            when x"0f" => output := x"76ec9a76";
            when x"10" => output := x"ca8f45ca";
            when x"11" => output := x"821f9d82";
            when x"12" => output := x"c98940c9";
            when x"13" => output := x"7dfa877d";
            when x"14" => output := x"faef15fa";
            when x"15" => output := x"59b2eb59";
            when x"16" => output := x"478ec947";
            when x"17" => output := x"f0fb0bf0";
            when x"18" => output := x"ad41ecad";
            when x"19" => output := x"d4b367d4";
            when x"1a" => output := x"a25ffda2";
            when x"1b" => output := x"af45eaaf";
            when x"1c" => output := x"9c23bf9c";
            when x"1d" => output := x"a453f7a4";
            when x"1e" => output := x"72e49672";
            when x"1f" => output := x"c09b5bc0";
            when x"20" => output := x"b775c2b7";
            when x"21" => output := x"fde11cfd";
            when x"22" => output := x"933dae93";
            when x"23" => output := x"264c6a26";
            when x"24" => output := x"366c5a36";
            when x"25" => output := x"3f7e413f";
            when x"26" => output := x"f7f502f7";
            when x"27" => output := x"cc834fcc";
            when x"28" => output := x"34685c34";
            when x"29" => output := x"a551f4a5";
            when x"2a" => output := x"e5d134e5";
            when x"2b" => output := x"f1f908f1";
            when x"2c" => output := x"71e29371";
            when x"2d" => output := x"d8ab73d8";
            when x"2e" => output := x"31625331";
            when x"2f" => output := x"152a3f15";
            when x"30" => output := x"04080c04";
            when x"31" => output := x"c79552c7";
            when x"32" => output := x"23466523";
            when x"33" => output := x"c39d5ec3";
            when x"34" => output := x"18302818";
            when x"35" => output := x"9637a196";
            when x"36" => output := x"050a0f05";
            when x"37" => output := x"9a2fb59a";
            when x"38" => output := x"070e0907";
            when x"39" => output := x"12243612";
            when x"3a" => output := x"801b9b80";
            when x"3b" => output := x"e2df3de2";
            when x"3c" => output := x"ebcd26eb";
            when x"3d" => output := x"274e6927";
            when x"3e" => output := x"b27fcdb2";
            when x"3f" => output := x"75ea9f75";
            when x"40" => output := x"09121b09";
            when x"41" => output := x"831d9e83";
            when x"42" => output := x"2c58742c";
            when x"43" => output := x"1a342e1a";
            when x"44" => output := x"1b362d1b";
            when x"45" => output := x"6edcb26e";
            when x"46" => output := x"5ab4ee5a";
            when x"47" => output := x"a05bfba0";
            when x"48" => output := x"52a4f652";
            when x"49" => output := x"3b764d3b";
            when x"4a" => output := x"d6b761d6";
            when x"4b" => output := x"b37dceb3";
            when x"4c" => output := x"29527b29";
            when x"4d" => output := x"e3dd3ee3";
            when x"4e" => output := x"2f5e712f";
            when x"4f" => output := x"84139784";
            when x"50" => output := x"53a6f553";
            when x"51" => output := x"d1b968d1";
            when x"52" => output := x"00000000";
            when x"53" => output := x"edc12ced";
            when x"54" => output := x"20406020";
            when x"55" => output := x"fce31ffc";
            when x"56" => output := x"b179c8b1";
            when x"57" => output := x"5bb6ed5b";
            when x"58" => output := x"6ad4be6a";
            when x"59" => output := x"cb8d46cb";
            when x"5a" => output := x"be67d9be";
            when x"5b" => output := x"39724b39";
            when x"5c" => output := x"4a94de4a";
            when x"5d" => output := x"4c98d44c";
            when x"5e" => output := x"58b0e858";
            when x"5f" => output := x"cf854acf";
            when x"60" => output := x"d0bb6bd0";
            when x"61" => output := x"efc52aef";
            when x"62" => output := x"aa4fe5aa";
            when x"63" => output := x"fbed16fb";
            when x"64" => output := x"4386c543";
            when x"65" => output := x"4d9ad74d";
            when x"66" => output := x"33665533";
            when x"67" => output := x"85119485";
            when x"68" => output := x"458acf45";
            when x"69" => output := x"f9e910f9";
            when x"6a" => output := x"02040602";
            when x"6b" => output := x"7ffe817f";
            when x"6c" => output := x"50a0f050";
            when x"6d" => output := x"3c78443c";
            when x"6e" => output := x"9f25ba9f";
            when x"6f" => output := x"a84be3a8";
            when x"70" => output := x"51a2f351";
            when x"71" => output := x"a35dfea3";
            when x"72" => output := x"4080c040";
            when x"73" => output := x"8f058a8f";
            when x"74" => output := x"923fad92";
            when x"75" => output := x"9d21bc9d";
            when x"76" => output := x"38704838";
            when x"77" => output := x"f5f104f5";
            when x"78" => output := x"bc63dfbc";
            when x"79" => output := x"b677c1b6";
            when x"7a" => output := x"daaf75da";
            when x"7b" => output := x"21426321";
            when x"7c" => output := x"10203010";
            when x"7d" => output := x"ffe51aff";
            when x"7e" => output := x"f3fd0ef3";
            when x"7f" => output := x"d2bf6dd2";
            when x"80" => output := x"cd814ccd";
            when x"81" => output := x"0c18140c";
            when x"82" => output := x"13263513";
            when x"83" => output := x"ecc32fec";
            when x"84" => output := x"5fbee15f";
            when x"85" => output := x"9735a297";
            when x"86" => output := x"4488cc44";
            when x"87" => output := x"172e3917";
            when x"88" => output := x"c49357c4";
            when x"89" => output := x"a755f2a7";
            when x"8a" => output := x"7efc827e";
            when x"8b" => output := x"3d7a473d";
            when x"8c" => output := x"64c8ac64";
            when x"8d" => output := x"5dbae75d";
            when x"8e" => output := x"19322b19";
            when x"8f" => output := x"73e69573";
            when x"90" => output := x"60c0a060";
            when x"91" => output := x"81199881";
            when x"92" => output := x"4f9ed14f";
            when x"93" => output := x"dca37fdc";
            when x"94" => output := x"22446622";
            when x"95" => output := x"2a547e2a";
            when x"96" => output := x"903bab90";
            when x"97" => output := x"880b8388";
            when x"98" => output := x"468cca46";
            when x"99" => output := x"eec729ee";
            when x"9a" => output := x"b86bd3b8";
            when x"9b" => output := x"14283c14";
            when x"9c" => output := x"dea779de";
            when x"9d" => output := x"5ebce25e";
            when x"9e" => output := x"0b161d0b";
            when x"9f" => output := x"dbad76db";
            when x"a0" => output := x"e0db3be0";
            when x"a1" => output := x"32645632";
            when x"a2" => output := x"3a744e3a";
            when x"a3" => output := x"0a141e0a";
            when x"a4" => output := x"4992db49";
            when x"a5" => output := x"060c0a06";
            when x"a6" => output := x"24486c24";
            when x"a7" => output := x"5cb8e45c";
            when x"a8" => output := x"c29f5dc2";
            when x"a9" => output := x"d3bd6ed3";
            when x"aa" => output := x"ac43efac";
            when x"ab" => output := x"62c4a662";
            when x"ac" => output := x"9139a891";
            when x"ad" => output := x"9531a495";
            when x"ae" => output := x"e4d337e4";
            when x"af" => output := x"79f28b79";
            when x"b0" => output := x"e7d532e7";
            when x"b1" => output := x"c88b43c8";
            when x"b2" => output := x"376e5937";
            when x"b3" => output := x"6ddab76d";
            when x"b4" => output := x"8d018c8d";
            when x"b5" => output := x"d5b164d5";
            when x"b6" => output := x"4e9cd24e";
            when x"b7" => output := x"a949e0a9";
            when x"b8" => output := x"6cd8b46c";
            when x"b9" => output := x"56acfa56";
            when x"ba" => output := x"f4f307f4";
            when x"bb" => output := x"eacf25ea";
            when x"bc" => output := x"65caaf65";
            when x"bd" => output := x"7af48e7a";
            when x"be" => output := x"ae47e9ae";
            when x"bf" => output := x"08101808";
            when x"c0" => output := x"ba6fd5ba";
            when x"c1" => output := x"78f08878";
            when x"c2" => output := x"254a6f25";
            when x"c3" => output := x"2e5c722e";
            when x"c4" => output := x"1c38241c";
            when x"c5" => output := x"a657f1a6";
            when x"c6" => output := x"b473c7b4";
            when x"c7" => output := x"c69751c6";
            when x"c8" => output := x"e8cb23e8";
            when x"c9" => output := x"dda17cdd";
            when x"ca" => output := x"74e89c74";
            when x"cb" => output := x"1f3e211f";
            when x"cc" => output := x"4b96dd4b";
            when x"cd" => output := x"bd61dcbd";
            when x"ce" => output := x"8b0d868b";
            when x"cf" => output := x"8a0f858a";
            when x"d0" => output := x"70e09070";
            when x"d1" => output := x"3e7c423e";
            when x"d2" => output := x"b571c4b5";
            when x"d3" => output := x"66ccaa66";
            when x"d4" => output := x"4890d848";
            when x"d5" => output := x"03060503";
            when x"d6" => output := x"f6f701f6";
            when x"d7" => output := x"0e1c120e";
            when x"d8" => output := x"61c2a361";
            when x"d9" => output := x"356a5f35";
            when x"da" => output := x"57aef957";
            when x"db" => output := x"b969d0b9";
            when x"dc" => output := x"86179186";
            when x"dd" => output := x"c19958c1";
            when x"de" => output := x"1d3a271d";
            when x"df" => output := x"9e27b99e";
            when x"e0" => output := x"e1d938e1";
            when x"e1" => output := x"f8eb13f8";
            when x"e2" => output := x"982bb398";
            when x"e3" => output := x"11223311";
            when x"e4" => output := x"69d2bb69";
            when x"e5" => output := x"d9a970d9";
            when x"e6" => output := x"8e07898e";
            when x"e7" => output := x"9433a794";
            when x"e8" => output := x"9b2db69b";
            when x"e9" => output := x"1e3c221e";
            when x"ea" => output := x"87159287";
            when x"eb" => output := x"e9c920e9";
            when x"ec" => output := x"ce8749ce";
            when x"ed" => output := x"55aaff55";
            when x"ee" => output := x"28507828";
            when x"ef" => output := x"dfa57adf";
            when x"f0" => output := x"8c038f8c";
            when x"f1" => output := x"a159f8a1";
            when x"f2" => output := x"89098089";
            when x"f3" => output := x"0d1a170d";
            when x"f4" => output := x"bf65dabf";
            when x"f5" => output := x"e6d731e6";
            when x"f6" => output := x"4284c642";
            when x"f7" => output := x"68d0b868";
            when x"f8" => output := x"4182c341";
            when x"f9" => output := x"9929b099";
            when x"fa" => output := x"2d5a772d";
            when x"fb" => output := x"0f1e110f";
            when x"fc" => output := x"b07bcbb0";
            when x"fd" => output := x"54a8fc54";
            when x"fe" => output := x"bb6dd6bb";
            when x"ff" => output := x"162c3a16";
            when others => null;
        end case;

        return output;
    end;

    function lutEnc3 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector is variable output : std_logic_vector(31 downto 0);
    begin
        case input is
            when x"00" => output := x"c6a56363";
            when x"01" => output := x"f8847c7c";
            when x"02" => output := x"ee997777";
            when x"03" => output := x"f68d7b7b";
            when x"04" => output := x"ff0df2f2";
            when x"05" => output := x"d6bd6b6b";
            when x"06" => output := x"deb16f6f";
            when x"07" => output := x"9154c5c5";
            when x"08" => output := x"60503030";
            when x"09" => output := x"02030101";
            when x"0a" => output := x"cea96767";
            when x"0b" => output := x"567d2b2b";
            when x"0c" => output := x"e719fefe";
            when x"0d" => output := x"b562d7d7";
            when x"0e" => output := x"4de6abab";
            when x"0f" => output := x"ec9a7676";
            when x"10" => output := x"8f45caca";
            when x"11" => output := x"1f9d8282";
            when x"12" => output := x"8940c9c9";
            when x"13" => output := x"fa877d7d";
            when x"14" => output := x"ef15fafa";
            when x"15" => output := x"b2eb5959";
            when x"16" => output := x"8ec94747";
            when x"17" => output := x"fb0bf0f0";
            when x"18" => output := x"41ecadad";
            when x"19" => output := x"b367d4d4";
            when x"1a" => output := x"5ffda2a2";
            when x"1b" => output := x"45eaafaf";
            when x"1c" => output := x"23bf9c9c";
            when x"1d" => output := x"53f7a4a4";
            when x"1e" => output := x"e4967272";
            when x"1f" => output := x"9b5bc0c0";
            when x"20" => output := x"75c2b7b7";
            when x"21" => output := x"e11cfdfd";
            when x"22" => output := x"3dae9393";
            when x"23" => output := x"4c6a2626";
            when x"24" => output := x"6c5a3636";
            when x"25" => output := x"7e413f3f";
            when x"26" => output := x"f502f7f7";
            when x"27" => output := x"834fcccc";
            when x"28" => output := x"685c3434";
            when x"29" => output := x"51f4a5a5";
            when x"2a" => output := x"d134e5e5";
            when x"2b" => output := x"f908f1f1";
            when x"2c" => output := x"e2937171";
            when x"2d" => output := x"ab73d8d8";
            when x"2e" => output := x"62533131";
            when x"2f" => output := x"2a3f1515";
            when x"30" => output := x"080c0404";
            when x"31" => output := x"9552c7c7";
            when x"32" => output := x"46652323";
            when x"33" => output := x"9d5ec3c3";
            when x"34" => output := x"30281818";
            when x"35" => output := x"37a19696";
            when x"36" => output := x"0a0f0505";
            when x"37" => output := x"2fb59a9a";
            when x"38" => output := x"0e090707";
            when x"39" => output := x"24361212";
            when x"3a" => output := x"1b9b8080";
            when x"3b" => output := x"df3de2e2";
            when x"3c" => output := x"cd26ebeb";
            when x"3d" => output := x"4e692727";
            when x"3e" => output := x"7fcdb2b2";
            when x"3f" => output := x"ea9f7575";
            when x"40" => output := x"121b0909";
            when x"41" => output := x"1d9e8383";
            when x"42" => output := x"58742c2c";
            when x"43" => output := x"342e1a1a";
            when x"44" => output := x"362d1b1b";
            when x"45" => output := x"dcb26e6e";
            when x"46" => output := x"b4ee5a5a";
            when x"47" => output := x"5bfba0a0";
            when x"48" => output := x"a4f65252";
            when x"49" => output := x"764d3b3b";
            when x"4a" => output := x"b761d6d6";
            when x"4b" => output := x"7dceb3b3";
            when x"4c" => output := x"527b2929";
            when x"4d" => output := x"dd3ee3e3";
            when x"4e" => output := x"5e712f2f";
            when x"4f" => output := x"13978484";
            when x"50" => output := x"a6f55353";
            when x"51" => output := x"b968d1d1";
            when x"52" => output := x"00000000";
            when x"53" => output := x"c12ceded";
            when x"54" => output := x"40602020";
            when x"55" => output := x"e31ffcfc";
            when x"56" => output := x"79c8b1b1";
            when x"57" => output := x"b6ed5b5b";
            when x"58" => output := x"d4be6a6a";
            when x"59" => output := x"8d46cbcb";
            when x"5a" => output := x"67d9bebe";
            when x"5b" => output := x"724b3939";
            when x"5c" => output := x"94de4a4a";
            when x"5d" => output := x"98d44c4c";
            when x"5e" => output := x"b0e85858";
            when x"5f" => output := x"854acfcf";
            when x"60" => output := x"bb6bd0d0";
            when x"61" => output := x"c52aefef";
            when x"62" => output := x"4fe5aaaa";
            when x"63" => output := x"ed16fbfb";
            when x"64" => output := x"86c54343";
            when x"65" => output := x"9ad74d4d";
            when x"66" => output := x"66553333";
            when x"67" => output := x"11948585";
            when x"68" => output := x"8acf4545";
            when x"69" => output := x"e910f9f9";
            when x"6a" => output := x"04060202";
            when x"6b" => output := x"fe817f7f";
            when x"6c" => output := x"a0f05050";
            when x"6d" => output := x"78443c3c";
            when x"6e" => output := x"25ba9f9f";
            when x"6f" => output := x"4be3a8a8";
            when x"70" => output := x"a2f35151";
            when x"71" => output := x"5dfea3a3";
            when x"72" => output := x"80c04040";
            when x"73" => output := x"058a8f8f";
            when x"74" => output := x"3fad9292";
            when x"75" => output := x"21bc9d9d";
            when x"76" => output := x"70483838";
            when x"77" => output := x"f104f5f5";
            when x"78" => output := x"63dfbcbc";
            when x"79" => output := x"77c1b6b6";
            when x"7a" => output := x"af75dada";
            when x"7b" => output := x"42632121";
            when x"7c" => output := x"20301010";
            when x"7d" => output := x"e51affff";
            when x"7e" => output := x"fd0ef3f3";
            when x"7f" => output := x"bf6dd2d2";
            when x"80" => output := x"814ccdcd";
            when x"81" => output := x"18140c0c";
            when x"82" => output := x"26351313";
            when x"83" => output := x"c32fecec";
            when x"84" => output := x"bee15f5f";
            when x"85" => output := x"35a29797";
            when x"86" => output := x"88cc4444";
            when x"87" => output := x"2e391717";
            when x"88" => output := x"9357c4c4";
            when x"89" => output := x"55f2a7a7";
            when x"8a" => output := x"fc827e7e";
            when x"8b" => output := x"7a473d3d";
            when x"8c" => output := x"c8ac6464";
            when x"8d" => output := x"bae75d5d";
            when x"8e" => output := x"322b1919";
            when x"8f" => output := x"e6957373";
            when x"90" => output := x"c0a06060";
            when x"91" => output := x"19988181";
            when x"92" => output := x"9ed14f4f";
            when x"93" => output := x"a37fdcdc";
            when x"94" => output := x"44662222";
            when x"95" => output := x"547e2a2a";
            when x"96" => output := x"3bab9090";
            when x"97" => output := x"0b838888";
            when x"98" => output := x"8cca4646";
            when x"99" => output := x"c729eeee";
            when x"9a" => output := x"6bd3b8b8";
            when x"9b" => output := x"283c1414";
            when x"9c" => output := x"a779dede";
            when x"9d" => output := x"bce25e5e";
            when x"9e" => output := x"161d0b0b";
            when x"9f" => output := x"ad76dbdb";
            when x"a0" => output := x"db3be0e0";
            when x"a1" => output := x"64563232";
            when x"a2" => output := x"744e3a3a";
            when x"a3" => output := x"141e0a0a";
            when x"a4" => output := x"92db4949";
            when x"a5" => output := x"0c0a0606";
            when x"a6" => output := x"486c2424";
            when x"a7" => output := x"b8e45c5c";
            when x"a8" => output := x"9f5dc2c2";
            when x"a9" => output := x"bd6ed3d3";
            when x"aa" => output := x"43efacac";
            when x"ab" => output := x"c4a66262";
            when x"ac" => output := x"39a89191";
            when x"ad" => output := x"31a49595";
            when x"ae" => output := x"d337e4e4";
            when x"af" => output := x"f28b7979";
            when x"b0" => output := x"d532e7e7";
            when x"b1" => output := x"8b43c8c8";
            when x"b2" => output := x"6e593737";
            when x"b3" => output := x"dab76d6d";
            when x"b4" => output := x"018c8d8d";
            when x"b5" => output := x"b164d5d5";
            when x"b6" => output := x"9cd24e4e";
            when x"b7" => output := x"49e0a9a9";
            when x"b8" => output := x"d8b46c6c";
            when x"b9" => output := x"acfa5656";
            when x"ba" => output := x"f307f4f4";
            when x"bb" => output := x"cf25eaea";
            when x"bc" => output := x"caaf6565";
            when x"bd" => output := x"f48e7a7a";
            when x"be" => output := x"47e9aeae";
            when x"bf" => output := x"10180808";
            when x"c0" => output := x"6fd5baba";
            when x"c1" => output := x"f0887878";
            when x"c2" => output := x"4a6f2525";
            when x"c3" => output := x"5c722e2e";
            when x"c4" => output := x"38241c1c";
            when x"c5" => output := x"57f1a6a6";
            when x"c6" => output := x"73c7b4b4";
            when x"c7" => output := x"9751c6c6";
            when x"c8" => output := x"cb23e8e8";
            when x"c9" => output := x"a17cdddd";
            when x"ca" => output := x"e89c7474";
            when x"cb" => output := x"3e211f1f";
            when x"cc" => output := x"96dd4b4b";
            when x"cd" => output := x"61dcbdbd";
            when x"ce" => output := x"0d868b8b";
            when x"cf" => output := x"0f858a8a";
            when x"d0" => output := x"e0907070";
            when x"d1" => output := x"7c423e3e";
            when x"d2" => output := x"71c4b5b5";
            when x"d3" => output := x"ccaa6666";
            when x"d4" => output := x"90d84848";
            when x"d5" => output := x"06050303";
            when x"d6" => output := x"f701f6f6";
            when x"d7" => output := x"1c120e0e";
            when x"d8" => output := x"c2a36161";
            when x"d9" => output := x"6a5f3535";
            when x"da" => output := x"aef95757";
            when x"db" => output := x"69d0b9b9";
            when x"dc" => output := x"17918686";
            when x"dd" => output := x"9958c1c1";
            when x"de" => output := x"3a271d1d";
            when x"df" => output := x"27b99e9e";
            when x"e0" => output := x"d938e1e1";
            when x"e1" => output := x"eb13f8f8";
            when x"e2" => output := x"2bb39898";
            when x"e3" => output := x"22331111";
            when x"e4" => output := x"d2bb6969";
            when x"e5" => output := x"a970d9d9";
            when x"e6" => output := x"07898e8e";
            when x"e7" => output := x"33a79494";
            when x"e8" => output := x"2db69b9b";
            when x"e9" => output := x"3c221e1e";
            when x"ea" => output := x"15928787";
            when x"eb" => output := x"c920e9e9";
            when x"ec" => output := x"8749cece";
            when x"ed" => output := x"aaff5555";
            when x"ee" => output := x"50782828";
            when x"ef" => output := x"a57adfdf";
            when x"f0" => output := x"038f8c8c";
            when x"f1" => output := x"59f8a1a1";
            when x"f2" => output := x"09808989";
            when x"f3" => output := x"1a170d0d";
            when x"f4" => output := x"65dabfbf";
            when x"f5" => output := x"d731e6e6";
            when x"f6" => output := x"84c64242";
            when x"f7" => output := x"d0b86868";
            when x"f8" => output := x"82c34141";
            when x"f9" => output := x"29b09999";
            when x"fa" => output := x"5a772d2d";
            when x"fb" => output := x"1e110f0f";
            when x"fc" => output := x"7bcbb0b0";
            when x"fd" => output := x"a8fc5454";
            when x"fe" => output := x"6dd6bbbb";
            when x"ff" => output := x"2c3a1616";
            when others => null;
        end case;

        return output;
    end;

    ------------------------------ DEC ------------------------------

    function lutDec0 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector is variable output : std_logic_vector(31 downto 0);
    begin
        case input is
            when x"00" => output := x"50a7f451";
            when x"01" => output := x"5365417e";
            when x"02" => output := x"c3a4171a";
            when x"03" => output := x"965e273a";
            when x"04" => output := x"cb6bab3b";
            when x"05" => output := x"f1459d1f";
            when x"06" => output := x"ab58faac";
            when x"07" => output := x"9303e34b";
            when x"08" => output := x"55fa3020";
            when x"09" => output := x"f66d76ad";
            when x"0a" => output := x"9176cc88";
            when x"0b" => output := x"254c02f5";
            when x"0c" => output := x"fcd7e54f";
            when x"0d" => output := x"d7cb2ac5";
            when x"0e" => output := x"80443526";
            when x"0f" => output := x"8fa362b5";
            when x"10" => output := x"495ab1de";
            when x"11" => output := x"671bba25";
            when x"12" => output := x"980eea45";
            when x"13" => output := x"e1c0fe5d";
            when x"14" => output := x"02752fc3";
            when x"15" => output := x"12f04c81";
            when x"16" => output := x"a397468d";
            when x"17" => output := x"c6f9d36b";
            when x"18" => output := x"e75f8f03";
            when x"19" => output := x"959c9215";
            when x"1a" => output := x"eb7a6dbf";
            when x"1b" => output := x"da595295";
            when x"1c" => output := x"2d83bed4";
            when x"1d" => output := x"d3217458";
            when x"1e" => output := x"2969e049";
            when x"1f" => output := x"44c8c98e";
            when x"20" => output := x"6a89c275";
            when x"21" => output := x"78798ef4";
            when x"22" => output := x"6b3e5899";
            when x"23" => output := x"dd71b927";
            when x"24" => output := x"b64fe1be";
            when x"25" => output := x"17ad88f0";
            when x"26" => output := x"66ac20c9";
            when x"27" => output := x"b43ace7d";
            when x"28" => output := x"184adf63";
            when x"29" => output := x"82311ae5";
            when x"2a" => output := x"60335197";
            when x"2b" => output := x"457f5362";
            when x"2c" => output := x"e07764b1";
            when x"2d" => output := x"84ae6bbb";
            when x"2e" => output := x"1ca081fe";
            when x"2f" => output := x"942b08f9";
            when x"30" => output := x"58684870";
            when x"31" => output := x"19fd458f";
            when x"32" => output := x"876cde94";
            when x"33" => output := x"b7f87b52";
            when x"34" => output := x"23d373ab";
            when x"35" => output := x"e2024b72";
            when x"36" => output := x"578f1fe3";
            when x"37" => output := x"2aab5566";
            when x"38" => output := x"0728ebb2";
            when x"39" => output := x"03c2b52f";
            when x"3a" => output := x"9a7bc586";
            when x"3b" => output := x"a50837d3";
            when x"3c" => output := x"f2872830";
            when x"3d" => output := x"b2a5bf23";
            when x"3e" => output := x"ba6a0302";
            when x"3f" => output := x"5c8216ed";
            when x"40" => output := x"2b1ccf8a";
            when x"41" => output := x"92b479a7";
            when x"42" => output := x"f0f207f3";
            when x"43" => output := x"a1e2694e";
            when x"44" => output := x"cdf4da65";
            when x"45" => output := x"d5be0506";
            when x"46" => output := x"1f6234d1";
            when x"47" => output := x"8afea6c4";
            when x"48" => output := x"9d532e34";
            when x"49" => output := x"a055f3a2";
            when x"4a" => output := x"32e18a05";
            when x"4b" => output := x"75ebf6a4";
            when x"4c" => output := x"39ec830b";
            when x"4d" => output := x"aaef6040";
            when x"4e" => output := x"069f715e";
            when x"4f" => output := x"51106ebd";
            when x"50" => output := x"f98a213e";
            when x"51" => output := x"3d06dd96";
            when x"52" => output := x"ae053edd";
            when x"53" => output := x"46bde64d";
            when x"54" => output := x"b58d5491";
            when x"55" => output := x"055dc471";
            when x"56" => output := x"6fd40604";
            when x"57" => output := x"ff155060";
            when x"58" => output := x"24fb9819";
            when x"59" => output := x"97e9bdd6";
            when x"5a" => output := x"cc434089";
            when x"5b" => output := x"779ed967";
            when x"5c" => output := x"bd42e8b0";
            when x"5d" => output := x"888b8907";
            when x"5e" => output := x"385b19e7";
            when x"5f" => output := x"dbeec879";
            when x"60" => output := x"470a7ca1";
            when x"61" => output := x"e90f427c";
            when x"62" => output := x"c91e84f8";
            when x"63" => output := x"00000000";
            when x"64" => output := x"83868009";
            when x"65" => output := x"48ed2b32";
            when x"66" => output := x"ac70111e";
            when x"67" => output := x"4e725a6c";
            when x"68" => output := x"fbff0efd";
            when x"69" => output := x"5638850f";
            when x"6a" => output := x"1ed5ae3d";
            when x"6b" => output := x"27392d36";
            when x"6c" => output := x"64d90f0a";
            when x"6d" => output := x"21a65c68";
            when x"6e" => output := x"d1545b9b";
            when x"6f" => output := x"3a2e3624";
            when x"70" => output := x"b1670a0c";
            when x"71" => output := x"0fe75793";
            when x"72" => output := x"d296eeb4";
            when x"73" => output := x"9e919b1b";
            when x"74" => output := x"4fc5c080";
            when x"75" => output := x"a220dc61";
            when x"76" => output := x"694b775a";
            when x"77" => output := x"161a121c";
            when x"78" => output := x"0aba93e2";
            when x"79" => output := x"e52aa0c0";
            when x"7a" => output := x"43e0223c";
            when x"7b" => output := x"1d171b12";
            when x"7c" => output := x"0b0d090e";
            when x"7d" => output := x"adc78bf2";
            when x"7e" => output := x"b9a8b62d";
            when x"7f" => output := x"c8a91e14";
            when x"80" => output := x"8519f157";
            when x"81" => output := x"4c0775af";
            when x"82" => output := x"bbdd99ee";
            when x"83" => output := x"fd607fa3";
            when x"84" => output := x"9f2601f7";
            when x"85" => output := x"bcf5725c";
            when x"86" => output := x"c53b6644";
            when x"87" => output := x"347efb5b";
            when x"88" => output := x"7629438b";
            when x"89" => output := x"dcc623cb";
            when x"8a" => output := x"68fcedb6";
            when x"8b" => output := x"63f1e4b8";
            when x"8c" => output := x"cadc31d7";
            when x"8d" => output := x"10856342";
            when x"8e" => output := x"40229713";
            when x"8f" => output := x"2011c684";
            when x"90" => output := x"7d244a85";
            when x"91" => output := x"f83dbbd2";
            when x"92" => output := x"1132f9ae";
            when x"93" => output := x"6da129c7";
            when x"94" => output := x"4b2f9e1d";
            when x"95" => output := x"f330b2dc";
            when x"96" => output := x"ec52860d";
            when x"97" => output := x"d0e3c177";
            when x"98" => output := x"6c16b32b";
            when x"99" => output := x"99b970a9";
            when x"9a" => output := x"fa489411";
            when x"9b" => output := x"2264e947";
            when x"9c" => output := x"c48cfca8";
            when x"9d" => output := x"1a3ff0a0";
            when x"9e" => output := x"d82c7d56";
            when x"9f" => output := x"ef903322";
            when x"a0" => output := x"c74e4987";
            when x"a1" => output := x"c1d138d9";
            when x"a2" => output := x"fea2ca8c";
            when x"a3" => output := x"360bd498";
            when x"a4" => output := x"cf81f5a6";
            when x"a5" => output := x"28de7aa5";
            when x"a6" => output := x"268eb7da";
            when x"a7" => output := x"a4bfad3f";
            when x"a8" => output := x"e49d3a2c";
            when x"a9" => output := x"0d927850";
            when x"aa" => output := x"9bcc5f6a";
            when x"ab" => output := x"62467e54";
            when x"ac" => output := x"c2138df6";
            when x"ad" => output := x"e8b8d890";
            when x"ae" => output := x"5ef7392e";
            when x"af" => output := x"f5afc382";
            when x"b0" => output := x"be805d9f";
            when x"b1" => output := x"7c93d069";
            when x"b2" => output := x"a92dd56f";
            when x"b3" => output := x"b31225cf";
            when x"b4" => output := x"3b99acc8";
            when x"b5" => output := x"a77d1810";
            when x"b6" => output := x"6e639ce8";
            when x"b7" => output := x"7bbb3bdb";
            when x"b8" => output := x"097826cd";
            when x"b9" => output := x"f418596e";
            when x"ba" => output := x"01b79aec";
            when x"bb" => output := x"a89a4f83";
            when x"bc" => output := x"656e95e6";
            when x"bd" => output := x"7ee6ffaa";
            when x"be" => output := x"08cfbc21";
            when x"bf" => output := x"e6e815ef";
            when x"c0" => output := x"d99be7ba";
            when x"c1" => output := x"ce366f4a";
            when x"c2" => output := x"d4099fea";
            when x"c3" => output := x"d67cb029";
            when x"c4" => output := x"afb2a431";
            when x"c5" => output := x"31233f2a";
            when x"c6" => output := x"3094a5c6";
            when x"c7" => output := x"c066a235";
            when x"c8" => output := x"37bc4e74";
            when x"c9" => output := x"a6ca82fc";
            when x"ca" => output := x"b0d090e0";
            when x"cb" => output := x"15d8a733";
            when x"cc" => output := x"4a9804f1";
            when x"cd" => output := x"f7daec41";
            when x"ce" => output := x"0e50cd7f";
            when x"cf" => output := x"2ff69117";
            when x"d0" => output := x"8dd64d76";
            when x"d1" => output := x"4db0ef43";
            when x"d2" => output := x"544daacc";
            when x"d3" => output := x"df0496e4";
            when x"d4" => output := x"e3b5d19e";
            when x"d5" => output := x"1b886a4c";
            when x"d6" => output := x"b81f2cc1";
            when x"d7" => output := x"7f516546";
            when x"d8" => output := x"04ea5e9d";
            when x"d9" => output := x"5d358c01";
            when x"da" => output := x"737487fa";
            when x"db" => output := x"2e410bfb";
            when x"dc" => output := x"5a1d67b3";
            when x"dd" => output := x"52d2db92";
            when x"de" => output := x"335610e9";
            when x"df" => output := x"1347d66d";
            when x"e0" => output := x"8c61d79a";
            when x"e1" => output := x"7a0ca137";
            when x"e2" => output := x"8e14f859";
            when x"e3" => output := x"893c13eb";
            when x"e4" => output := x"ee27a9ce";
            when x"e5" => output := x"35c961b7";
            when x"e6" => output := x"ede51ce1";
            when x"e7" => output := x"3cb1477a";
            when x"e8" => output := x"59dfd29c";
            when x"e9" => output := x"3f73f255";
            when x"ea" => output := x"79ce1418";
            when x"eb" => output := x"bf37c773";
            when x"ec" => output := x"eacdf753";
            when x"ed" => output := x"5baafd5f";
            when x"ee" => output := x"146f3ddf";
            when x"ef" => output := x"86db4478";
            when x"f0" => output := x"81f3afca";
            when x"f1" => output := x"3ec468b9";
            when x"f2" => output := x"2c342438";
            when x"f3" => output := x"5f40a3c2";
            when x"f4" => output := x"72c31d16";
            when x"f5" => output := x"0c25e2bc";
            when x"f6" => output := x"8b493c28";
            when x"f7" => output := x"41950dff";
            when x"f8" => output := x"7101a839";
            when x"f9" => output := x"deb30c08";
            when x"fa" => output := x"9ce4b4d8";
            when x"fb" => output := x"90c15664";
            when x"fc" => output := x"6184cb7b";
            when x"fd" => output := x"70b632d5";
            when x"fe" => output := x"745c6c48";
            when x"ff" => output := x"4257b8d0";
            when others => null;
        end case;

        return output;
    end;

    function lutDec1 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector is variable output : std_logic_vector(31 downto 0);
    begin
        case input is
            when x"00" => output := x"a7f45150";
            when x"01" => output := x"65417e53";
            when x"02" => output := x"a4171ac3";
            when x"03" => output := x"5e273a96";
            when x"04" => output := x"6bab3bcb";
            when x"05" => output := x"459d1ff1";
            when x"06" => output := x"58faacab";
            when x"07" => output := x"03e34b93";
            when x"08" => output := x"fa302055";
            when x"09" => output := x"6d76adf6";
            when x"0a" => output := x"76cc8891";
            when x"0b" => output := x"4c02f525";
            when x"0c" => output := x"d7e54ffc";
            when x"0d" => output := x"cb2ac5d7";
            when x"0e" => output := x"44352680";
            when x"0f" => output := x"a362b58f";
            when x"10" => output := x"5ab1de49";
            when x"11" => output := x"1bba2567";
            when x"12" => output := x"0eea4598";
            when x"13" => output := x"c0fe5de1";
            when x"14" => output := x"752fc302";
            when x"15" => output := x"f04c8112";
            when x"16" => output := x"97468da3";
            when x"17" => output := x"f9d36bc6";
            when x"18" => output := x"5f8f03e7";
            when x"19" => output := x"9c921595";
            when x"1a" => output := x"7a6dbfeb";
            when x"1b" => output := x"595295da";
            when x"1c" => output := x"83bed42d";
            when x"1d" => output := x"217458d3";
            when x"1e" => output := x"69e04929";
            when x"1f" => output := x"c8c98e44";
            when x"20" => output := x"89c2756a";
            when x"21" => output := x"798ef478";
            when x"22" => output := x"3e58996b";
            when x"23" => output := x"71b927dd";
            when x"24" => output := x"4fe1beb6";
            when x"25" => output := x"ad88f017";
            when x"26" => output := x"ac20c966";
            when x"27" => output := x"3ace7db4";
            when x"28" => output := x"4adf6318";
            when x"29" => output := x"311ae582";
            when x"2a" => output := x"33519760";
            when x"2b" => output := x"7f536245";
            when x"2c" => output := x"7764b1e0";
            when x"2d" => output := x"ae6bbb84";
            when x"2e" => output := x"a081fe1c";
            when x"2f" => output := x"2b08f994";
            when x"30" => output := x"68487058";
            when x"31" => output := x"fd458f19";
            when x"32" => output := x"6cde9487";
            when x"33" => output := x"f87b52b7";
            when x"34" => output := x"d373ab23";
            when x"35" => output := x"024b72e2";
            when x"36" => output := x"8f1fe357";
            when x"37" => output := x"ab55662a";
            when x"38" => output := x"28ebb207";
            when x"39" => output := x"c2b52f03";
            when x"3a" => output := x"7bc5869a";
            when x"3b" => output := x"0837d3a5";
            when x"3c" => output := x"872830f2";
            when x"3d" => output := x"a5bf23b2";
            when x"3e" => output := x"6a0302ba";
            when x"3f" => output := x"8216ed5c";
            when x"40" => output := x"1ccf8a2b";
            when x"41" => output := x"b479a792";
            when x"42" => output := x"f207f3f0";
            when x"43" => output := x"e2694ea1";
            when x"44" => output := x"f4da65cd";
            when x"45" => output := x"be0506d5";
            when x"46" => output := x"6234d11f";
            when x"47" => output := x"fea6c48a";
            when x"48" => output := x"532e349d";
            when x"49" => output := x"55f3a2a0";
            when x"4a" => output := x"e18a0532";
            when x"4b" => output := x"ebf6a475";
            when x"4c" => output := x"ec830b39";
            when x"4d" => output := x"ef6040aa";
            when x"4e" => output := x"9f715e06";
            when x"4f" => output := x"106ebd51";
            when x"50" => output := x"8a213ef9";
            when x"51" => output := x"06dd963d";
            when x"52" => output := x"053eddae";
            when x"53" => output := x"bde64d46";
            when x"54" => output := x"8d5491b5";
            when x"55" => output := x"5dc47105";
            when x"56" => output := x"d406046f";
            when x"57" => output := x"155060ff";
            when x"58" => output := x"fb981924";
            when x"59" => output := x"e9bdd697";
            when x"5a" => output := x"434089cc";
            when x"5b" => output := x"9ed96777";
            when x"5c" => output := x"42e8b0bd";
            when x"5d" => output := x"8b890788";
            when x"5e" => output := x"5b19e738";
            when x"5f" => output := x"eec879db";
            when x"60" => output := x"0a7ca147";
            when x"61" => output := x"0f427ce9";
            when x"62" => output := x"1e84f8c9";
            when x"63" => output := x"00000000";
            when x"64" => output := x"86800983";
            when x"65" => output := x"ed2b3248";
            when x"66" => output := x"70111eac";
            when x"67" => output := x"725a6c4e";
            when x"68" => output := x"ff0efdfb";
            when x"69" => output := x"38850f56";
            when x"6a" => output := x"d5ae3d1e";
            when x"6b" => output := x"392d3627";
            when x"6c" => output := x"d90f0a64";
            when x"6d" => output := x"a65c6821";
            when x"6e" => output := x"545b9bd1";
            when x"6f" => output := x"2e36243a";
            when x"70" => output := x"670a0cb1";
            when x"71" => output := x"e757930f";
            when x"72" => output := x"96eeb4d2";
            when x"73" => output := x"919b1b9e";
            when x"74" => output := x"c5c0804f";
            when x"75" => output := x"20dc61a2";
            when x"76" => output := x"4b775a69";
            when x"77" => output := x"1a121c16";
            when x"78" => output := x"ba93e20a";
            when x"79" => output := x"2aa0c0e5";
            when x"7a" => output := x"e0223c43";
            when x"7b" => output := x"171b121d";
            when x"7c" => output := x"0d090e0b";
            when x"7d" => output := x"c78bf2ad";
            when x"7e" => output := x"a8b62db9";
            when x"7f" => output := x"a91e14c8";
            when x"80" => output := x"19f15785";
            when x"81" => output := x"0775af4c";
            when x"82" => output := x"dd99eebb";
            when x"83" => output := x"607fa3fd";
            when x"84" => output := x"2601f79f";
            when x"85" => output := x"f5725cbc";
            when x"86" => output := x"3b6644c5";
            when x"87" => output := x"7efb5b34";
            when x"88" => output := x"29438b76";
            when x"89" => output := x"c623cbdc";
            when x"8a" => output := x"fcedb668";
            when x"8b" => output := x"f1e4b863";
            when x"8c" => output := x"dc31d7ca";
            when x"8d" => output := x"85634210";
            when x"8e" => output := x"22971340";
            when x"8f" => output := x"11c68420";
            when x"90" => output := x"244a857d";
            when x"91" => output := x"3dbbd2f8";
            when x"92" => output := x"32f9ae11";
            when x"93" => output := x"a129c76d";
            when x"94" => output := x"2f9e1d4b";
            when x"95" => output := x"30b2dcf3";
            when x"96" => output := x"52860dec";
            when x"97" => output := x"e3c177d0";
            when x"98" => output := x"16b32b6c";
            when x"99" => output := x"b970a999";
            when x"9a" => output := x"489411fa";
            when x"9b" => output := x"64e94722";
            when x"9c" => output := x"8cfca8c4";
            when x"9d" => output := x"3ff0a01a";
            when x"9e" => output := x"2c7d56d8";
            when x"9f" => output := x"903322ef";
            when x"a0" => output := x"4e4987c7";
            when x"a1" => output := x"d138d9c1";
            when x"a2" => output := x"a2ca8cfe";
            when x"a3" => output := x"0bd49836";
            when x"a4" => output := x"81f5a6cf";
            when x"a5" => output := x"de7aa528";
            when x"a6" => output := x"8eb7da26";
            when x"a7" => output := x"bfad3fa4";
            when x"a8" => output := x"9d3a2ce4";
            when x"a9" => output := x"9278500d";
            when x"aa" => output := x"cc5f6a9b";
            when x"ab" => output := x"467e5462";
            when x"ac" => output := x"138df6c2";
            when x"ad" => output := x"b8d890e8";
            when x"ae" => output := x"f7392e5e";
            when x"af" => output := x"afc382f5";
            when x"b0" => output := x"805d9fbe";
            when x"b1" => output := x"93d0697c";
            when x"b2" => output := x"2dd56fa9";
            when x"b3" => output := x"1225cfb3";
            when x"b4" => output := x"99acc83b";
            when x"b5" => output := x"7d1810a7";
            when x"b6" => output := x"639ce86e";
            when x"b7" => output := x"bb3bdb7b";
            when x"b8" => output := x"7826cd09";
            when x"b9" => output := x"18596ef4";
            when x"ba" => output := x"b79aec01";
            when x"bb" => output := x"9a4f83a8";
            when x"bc" => output := x"6e95e665";
            when x"bd" => output := x"e6ffaa7e";
            when x"be" => output := x"cfbc2108";
            when x"bf" => output := x"e815efe6";
            when x"c0" => output := x"9be7bad9";
            when x"c1" => output := x"366f4ace";
            when x"c2" => output := x"099fead4";
            when x"c3" => output := x"7cb029d6";
            when x"c4" => output := x"b2a431af";
            when x"c5" => output := x"233f2a31";
            when x"c6" => output := x"94a5c630";
            when x"c7" => output := x"66a235c0";
            when x"c8" => output := x"bc4e7437";
            when x"c9" => output := x"ca82fca6";
            when x"ca" => output := x"d090e0b0";
            when x"cb" => output := x"d8a73315";
            when x"cc" => output := x"9804f14a";
            when x"cd" => output := x"daec41f7";
            when x"ce" => output := x"50cd7f0e";
            when x"cf" => output := x"f691172f";
            when x"d0" => output := x"d64d768d";
            when x"d1" => output := x"b0ef434d";
            when x"d2" => output := x"4daacc54";
            when x"d3" => output := x"0496e4df";
            when x"d4" => output := x"b5d19ee3";
            when x"d5" => output := x"886a4c1b";
            when x"d6" => output := x"1f2cc1b8";
            when x"d7" => output := x"5165467f";
            when x"d8" => output := x"ea5e9d04";
            when x"d9" => output := x"358c015d";
            when x"da" => output := x"7487fa73";
            when x"db" => output := x"410bfb2e";
            when x"dc" => output := x"1d67b35a";
            when x"dd" => output := x"d2db9252";
            when x"de" => output := x"5610e933";
            when x"df" => output := x"47d66d13";
            when x"e0" => output := x"61d79a8c";
            when x"e1" => output := x"0ca1377a";
            when x"e2" => output := x"14f8598e";
            when x"e3" => output := x"3c13eb89";
            when x"e4" => output := x"27a9ceee";
            when x"e5" => output := x"c961b735";
            when x"e6" => output := x"e51ce1ed";
            when x"e7" => output := x"b1477a3c";
            when x"e8" => output := x"dfd29c59";
            when x"e9" => output := x"73f2553f";
            when x"ea" => output := x"ce141879";
            when x"eb" => output := x"37c773bf";
            when x"ec" => output := x"cdf753ea";
            when x"ed" => output := x"aafd5f5b";
            when x"ee" => output := x"6f3ddf14";
            when x"ef" => output := x"db447886";
            when x"f0" => output := x"f3afca81";
            when x"f1" => output := x"c468b93e";
            when x"f2" => output := x"3424382c";
            when x"f3" => output := x"40a3c25f";
            when x"f4" => output := x"c31d1672";
            when x"f5" => output := x"25e2bc0c";
            when x"f6" => output := x"493c288b";
            when x"f7" => output := x"950dff41";
            when x"f8" => output := x"01a83971";
            when x"f9" => output := x"b30c08de";
            when x"fa" => output := x"e4b4d89c";
            when x"fb" => output := x"c1566490";
            when x"fc" => output := x"84cb7b61";
            when x"fd" => output := x"b632d570";
            when x"fe" => output := x"5c6c4874";
            when x"ff" => output := x"57b8d042";
            when others => null;
        end case;

        return output;
    end;

    function lutDec2 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector is variable output : std_logic_vector(31 downto 0);
    begin
        case input is
            when x"00" => output := x"f45150a7";
            when x"01" => output := x"417e5365";
            when x"02" => output := x"171ac3a4";
            when x"03" => output := x"273a965e";
            when x"04" => output := x"ab3bcb6b";
            when x"05" => output := x"9d1ff145";
            when x"06" => output := x"faacab58";
            when x"07" => output := x"e34b9303";
            when x"08" => output := x"302055fa";
            when x"09" => output := x"76adf66d";
            when x"0a" => output := x"cc889176";
            when x"0b" => output := x"02f5254c";
            when x"0c" => output := x"e54ffcd7";
            when x"0d" => output := x"2ac5d7cb";
            when x"0e" => output := x"35268044";
            when x"0f" => output := x"62b58fa3";
            when x"10" => output := x"b1de495a";
            when x"11" => output := x"ba25671b";
            when x"12" => output := x"ea45980e";
            when x"13" => output := x"fe5de1c0";
            when x"14" => output := x"2fc30275";
            when x"15" => output := x"4c8112f0";
            when x"16" => output := x"468da397";
            when x"17" => output := x"d36bc6f9";
            when x"18" => output := x"8f03e75f";
            when x"19" => output := x"9215959c";
            when x"1a" => output := x"6dbfeb7a";
            when x"1b" => output := x"5295da59";
            when x"1c" => output := x"bed42d83";
            when x"1d" => output := x"7458d321";
            when x"1e" => output := x"e0492969";
            when x"1f" => output := x"c98e44c8";
            when x"20" => output := x"c2756a89";
            when x"21" => output := x"8ef47879";
            when x"22" => output := x"58996b3e";
            when x"23" => output := x"b927dd71";
            when x"24" => output := x"e1beb64f";
            when x"25" => output := x"88f017ad";
            when x"26" => output := x"20c966ac";
            when x"27" => output := x"ce7db43a";
            when x"28" => output := x"df63184a";
            when x"29" => output := x"1ae58231";
            when x"2a" => output := x"51976033";
            when x"2b" => output := x"5362457f";
            when x"2c" => output := x"64b1e077";
            when x"2d" => output := x"6bbb84ae";
            when x"2e" => output := x"81fe1ca0";
            when x"2f" => output := x"08f9942b";
            when x"30" => output := x"48705868";
            when x"31" => output := x"458f19fd";
            when x"32" => output := x"de94876c";
            when x"33" => output := x"7b52b7f8";
            when x"34" => output := x"73ab23d3";
            when x"35" => output := x"4b72e202";
            when x"36" => output := x"1fe3578f";
            when x"37" => output := x"55662aab";
            when x"38" => output := x"ebb20728";
            when x"39" => output := x"b52f03c2";
            when x"3a" => output := x"c5869a7b";
            when x"3b" => output := x"37d3a508";
            when x"3c" => output := x"2830f287";
            when x"3d" => output := x"bf23b2a5";
            when x"3e" => output := x"0302ba6a";
            when x"3f" => output := x"16ed5c82";
            when x"40" => output := x"cf8a2b1c";
            when x"41" => output := x"79a792b4";
            when x"42" => output := x"07f3f0f2";
            when x"43" => output := x"694ea1e2";
            when x"44" => output := x"da65cdf4";
            when x"45" => output := x"0506d5be";
            when x"46" => output := x"34d11f62";
            when x"47" => output := x"a6c48afe";
            when x"48" => output := x"2e349d53";
            when x"49" => output := x"f3a2a055";
            when x"4a" => output := x"8a0532e1";
            when x"4b" => output := x"f6a475eb";
            when x"4c" => output := x"830b39ec";
            when x"4d" => output := x"6040aaef";
            when x"4e" => output := x"715e069f";
            when x"4f" => output := x"6ebd5110";
            when x"50" => output := x"213ef98a";
            when x"51" => output := x"dd963d06";
            when x"52" => output := x"3eddae05";
            when x"53" => output := x"e64d46bd";
            when x"54" => output := x"5491b58d";
            when x"55" => output := x"c471055d";
            when x"56" => output := x"06046fd4";
            when x"57" => output := x"5060ff15";
            when x"58" => output := x"981924fb";
            when x"59" => output := x"bdd697e9";
            when x"5a" => output := x"4089cc43";
            when x"5b" => output := x"d967779e";
            when x"5c" => output := x"e8b0bd42";
            when x"5d" => output := x"8907888b";
            when x"5e" => output := x"19e7385b";
            when x"5f" => output := x"c879dbee";
            when x"60" => output := x"7ca1470a";
            when x"61" => output := x"427ce90f";
            when x"62" => output := x"84f8c91e";
            when x"63" => output := x"00000000";
            when x"64" => output := x"80098386";
            when x"65" => output := x"2b3248ed";
            when x"66" => output := x"111eac70";
            when x"67" => output := x"5a6c4e72";
            when x"68" => output := x"0efdfbff";
            when x"69" => output := x"850f5638";
            when x"6a" => output := x"ae3d1ed5";
            when x"6b" => output := x"2d362739";
            when x"6c" => output := x"0f0a64d9";
            when x"6d" => output := x"5c6821a6";
            when x"6e" => output := x"5b9bd154";
            when x"6f" => output := x"36243a2e";
            when x"70" => output := x"0a0cb167";
            when x"71" => output := x"57930fe7";
            when x"72" => output := x"eeb4d296";
            when x"73" => output := x"9b1b9e91";
            when x"74" => output := x"c0804fc5";
            when x"75" => output := x"dc61a220";
            when x"76" => output := x"775a694b";
            when x"77" => output := x"121c161a";
            when x"78" => output := x"93e20aba";
            when x"79" => output := x"a0c0e52a";
            when x"7a" => output := x"223c43e0";
            when x"7b" => output := x"1b121d17";
            when x"7c" => output := x"090e0b0d";
            when x"7d" => output := x"8bf2adc7";
            when x"7e" => output := x"b62db9a8";
            when x"7f" => output := x"1e14c8a9";
            when x"80" => output := x"f1578519";
            when x"81" => output := x"75af4c07";
            when x"82" => output := x"99eebbdd";
            when x"83" => output := x"7fa3fd60";
            when x"84" => output := x"01f79f26";
            when x"85" => output := x"725cbcf5";
            when x"86" => output := x"6644c53b";
            when x"87" => output := x"fb5b347e";
            when x"88" => output := x"438b7629";
            when x"89" => output := x"23cbdcc6";
            when x"8a" => output := x"edb668fc";
            when x"8b" => output := x"e4b863f1";
            when x"8c" => output := x"31d7cadc";
            when x"8d" => output := x"63421085";
            when x"8e" => output := x"97134022";
            when x"8f" => output := x"c6842011";
            when x"90" => output := x"4a857d24";
            when x"91" => output := x"bbd2f83d";
            when x"92" => output := x"f9ae1132";
            when x"93" => output := x"29c76da1";
            when x"94" => output := x"9e1d4b2f";
            when x"95" => output := x"b2dcf330";
            when x"96" => output := x"860dec52";
            when x"97" => output := x"c177d0e3";
            when x"98" => output := x"b32b6c16";
            when x"99" => output := x"70a999b9";
            when x"9a" => output := x"9411fa48";
            when x"9b" => output := x"e9472264";
            when x"9c" => output := x"fca8c48c";
            when x"9d" => output := x"f0a01a3f";
            when x"9e" => output := x"7d56d82c";
            when x"9f" => output := x"3322ef90";
            when x"a0" => output := x"4987c74e";
            when x"a1" => output := x"38d9c1d1";
            when x"a2" => output := x"ca8cfea2";
            when x"a3" => output := x"d498360b";
            when x"a4" => output := x"f5a6cf81";
            when x"a5" => output := x"7aa528de";
            when x"a6" => output := x"b7da268e";
            when x"a7" => output := x"ad3fa4bf";
            when x"a8" => output := x"3a2ce49d";
            when x"a9" => output := x"78500d92";
            when x"aa" => output := x"5f6a9bcc";
            when x"ab" => output := x"7e546246";
            when x"ac" => output := x"8df6c213";
            when x"ad" => output := x"d890e8b8";
            when x"ae" => output := x"392e5ef7";
            when x"af" => output := x"c382f5af";
            when x"b0" => output := x"5d9fbe80";
            when x"b1" => output := x"d0697c93";
            when x"b2" => output := x"d56fa92d";
            when x"b3" => output := x"25cfb312";
            when x"b4" => output := x"acc83b99";
            when x"b5" => output := x"1810a77d";
            when x"b6" => output := x"9ce86e63";
            when x"b7" => output := x"3bdb7bbb";
            when x"b8" => output := x"26cd0978";
            when x"b9" => output := x"596ef418";
            when x"ba" => output := x"9aec01b7";
            when x"bb" => output := x"4f83a89a";
            when x"bc" => output := x"95e6656e";
            when x"bd" => output := x"ffaa7ee6";
            when x"be" => output := x"bc2108cf";
            when x"bf" => output := x"15efe6e8";
            when x"c0" => output := x"e7bad99b";
            when x"c1" => output := x"6f4ace36";
            when x"c2" => output := x"9fead409";
            when x"c3" => output := x"b029d67c";
            when x"c4" => output := x"a431afb2";
            when x"c5" => output := x"3f2a3123";
            when x"c6" => output := x"a5c63094";
            when x"c7" => output := x"a235c066";
            when x"c8" => output := x"4e7437bc";
            when x"c9" => output := x"82fca6ca";
            when x"ca" => output := x"90e0b0d0";
            when x"cb" => output := x"a73315d8";
            when x"cc" => output := x"04f14a98";
            when x"cd" => output := x"ec41f7da";
            when x"ce" => output := x"cd7f0e50";
            when x"cf" => output := x"91172ff6";
            when x"d0" => output := x"4d768dd6";
            when x"d1" => output := x"ef434db0";
            when x"d2" => output := x"aacc544d";
            when x"d3" => output := x"96e4df04";
            when x"d4" => output := x"d19ee3b5";
            when x"d5" => output := x"6a4c1b88";
            when x"d6" => output := x"2cc1b81f";
            when x"d7" => output := x"65467f51";
            when x"d8" => output := x"5e9d04ea";
            when x"d9" => output := x"8c015d35";
            when x"da" => output := x"87fa7374";
            when x"db" => output := x"0bfb2e41";
            when x"dc" => output := x"67b35a1d";
            when x"dd" => output := x"db9252d2";
            when x"de" => output := x"10e93356";
            when x"df" => output := x"d66d1347";
            when x"e0" => output := x"d79a8c61";
            when x"e1" => output := x"a1377a0c";
            when x"e2" => output := x"f8598e14";
            when x"e3" => output := x"13eb893c";
            when x"e4" => output := x"a9ceee27";
            when x"e5" => output := x"61b735c9";
            when x"e6" => output := x"1ce1ede5";
            when x"e7" => output := x"477a3cb1";
            when x"e8" => output := x"d29c59df";
            when x"e9" => output := x"f2553f73";
            when x"ea" => output := x"141879ce";
            when x"eb" => output := x"c773bf37";
            when x"ec" => output := x"f753eacd";
            when x"ed" => output := x"fd5f5baa";
            when x"ee" => output := x"3ddf146f";
            when x"ef" => output := x"447886db";
            when x"f0" => output := x"afca81f3";
            when x"f1" => output := x"68b93ec4";
            when x"f2" => output := x"24382c34";
            when x"f3" => output := x"a3c25f40";
            when x"f4" => output := x"1d1672c3";
            when x"f5" => output := x"e2bc0c25";
            when x"f6" => output := x"3c288b49";
            when x"f7" => output := x"0dff4195";
            when x"f8" => output := x"a8397101";
            when x"f9" => output := x"0c08deb3";
            when x"fa" => output := x"b4d89ce4";
            when x"fb" => output := x"566490c1";
            when x"fc" => output := x"cb7b6184";
            when x"fd" => output := x"32d570b6";
            when x"fe" => output := x"6c48745c";
            when x"ff" => output := x"b8d04257";
            when others => null;
        end case;

        return output;
    end;

    function lutDec3 (input : in std_logic_vector(7 downto 0))
        return std_logic_vector is variable output : std_logic_vector(31 downto 0);
    begin
        case input is
            when x"00" => output := x"5150a7f4";
            when x"01" => output := x"7e536541";
            when x"02" => output := x"1ac3a417";
            when x"03" => output := x"3a965e27";
            when x"04" => output := x"3bcb6bab";
            when x"05" => output := x"1ff1459d";
            when x"06" => output := x"acab58fa";
            when x"07" => output := x"4b9303e3";
            when x"08" => output := x"2055fa30";
            when x"09" => output := x"adf66d76";
            when x"0a" => output := x"889176cc";
            when x"0b" => output := x"f5254c02";
            when x"0c" => output := x"4ffcd7e5";
            when x"0d" => output := x"c5d7cb2a";
            when x"0e" => output := x"26804435";
            when x"0f" => output := x"b58fa362";
            when x"10" => output := x"de495ab1";
            when x"11" => output := x"25671bba";
            when x"12" => output := x"45980eea";
            when x"13" => output := x"5de1c0fe";
            when x"14" => output := x"c302752f";
            when x"15" => output := x"8112f04c";
            when x"16" => output := x"8da39746";
            when x"17" => output := x"6bc6f9d3";
            when x"18" => output := x"03e75f8f";
            when x"19" => output := x"15959c92";
            when x"1a" => output := x"bfeb7a6d";
            when x"1b" => output := x"95da5952";
            when x"1c" => output := x"d42d83be";
            when x"1d" => output := x"58d32174";
            when x"1e" => output := x"492969e0";
            when x"1f" => output := x"8e44c8c9";
            when x"20" => output := x"756a89c2";
            when x"21" => output := x"f478798e";
            when x"22" => output := x"996b3e58";
            when x"23" => output := x"27dd71b9";
            when x"24" => output := x"beb64fe1";
            when x"25" => output := x"f017ad88";
            when x"26" => output := x"c966ac20";
            when x"27" => output := x"7db43ace";
            when x"28" => output := x"63184adf";
            when x"29" => output := x"e582311a";
            when x"2a" => output := x"97603351";
            when x"2b" => output := x"62457f53";
            when x"2c" => output := x"b1e07764";
            when x"2d" => output := x"bb84ae6b";
            when x"2e" => output := x"fe1ca081";
            when x"2f" => output := x"f9942b08";
            when x"30" => output := x"70586848";
            when x"31" => output := x"8f19fd45";
            when x"32" => output := x"94876cde";
            when x"33" => output := x"52b7f87b";
            when x"34" => output := x"ab23d373";
            when x"35" => output := x"72e2024b";
            when x"36" => output := x"e3578f1f";
            when x"37" => output := x"662aab55";
            when x"38" => output := x"b20728eb";
            when x"39" => output := x"2f03c2b5";
            when x"3a" => output := x"869a7bc5";
            when x"3b" => output := x"d3a50837";
            when x"3c" => output := x"30f28728";
            when x"3d" => output := x"23b2a5bf";
            when x"3e" => output := x"02ba6a03";
            when x"3f" => output := x"ed5c8216";
            when x"40" => output := x"8a2b1ccf";
            when x"41" => output := x"a792b479";
            when x"42" => output := x"f3f0f207";
            when x"43" => output := x"4ea1e269";
            when x"44" => output := x"65cdf4da";
            when x"45" => output := x"06d5be05";
            when x"46" => output := x"d11f6234";
            when x"47" => output := x"c48afea6";
            when x"48" => output := x"349d532e";
            when x"49" => output := x"a2a055f3";
            when x"4a" => output := x"0532e18a";
            when x"4b" => output := x"a475ebf6";
            when x"4c" => output := x"0b39ec83";
            when x"4d" => output := x"40aaef60";
            when x"4e" => output := x"5e069f71";
            when x"4f" => output := x"bd51106e";
            when x"50" => output := x"3ef98a21";
            when x"51" => output := x"963d06dd";
            when x"52" => output := x"ddae053e";
            when x"53" => output := x"4d46bde6";
            when x"54" => output := x"91b58d54";
            when x"55" => output := x"71055dc4";
            when x"56" => output := x"046fd406";
            when x"57" => output := x"60ff1550";
            when x"58" => output := x"1924fb98";
            when x"59" => output := x"d697e9bd";
            when x"5a" => output := x"89cc4340";
            when x"5b" => output := x"67779ed9";
            when x"5c" => output := x"b0bd42e8";
            when x"5d" => output := x"07888b89";
            when x"5e" => output := x"e7385b19";
            when x"5f" => output := x"79dbeec8";
            when x"60" => output := x"a1470a7c";
            when x"61" => output := x"7ce90f42";
            when x"62" => output := x"f8c91e84";
            when x"63" => output := x"00000000";
            when x"64" => output := x"09838680";
            when x"65" => output := x"3248ed2b";
            when x"66" => output := x"1eac7011";
            when x"67" => output := x"6c4e725a";
            when x"68" => output := x"fdfbff0e";
            when x"69" => output := x"0f563885";
            when x"6a" => output := x"3d1ed5ae";
            when x"6b" => output := x"3627392d";
            when x"6c" => output := x"0a64d90f";
            when x"6d" => output := x"6821a65c";
            when x"6e" => output := x"9bd1545b";
            when x"6f" => output := x"243a2e36";
            when x"70" => output := x"0cb1670a";
            when x"71" => output := x"930fe757";
            when x"72" => output := x"b4d296ee";
            when x"73" => output := x"1b9e919b";
            when x"74" => output := x"804fc5c0";
            when x"75" => output := x"61a220dc";
            when x"76" => output := x"5a694b77";
            when x"77" => output := x"1c161a12";
            when x"78" => output := x"e20aba93";
            when x"79" => output := x"c0e52aa0";
            when x"7a" => output := x"3c43e022";
            when x"7b" => output := x"121d171b";
            when x"7c" => output := x"0e0b0d09";
            when x"7d" => output := x"f2adc78b";
            when x"7e" => output := x"2db9a8b6";
            when x"7f" => output := x"14c8a91e";
            when x"80" => output := x"578519f1";
            when x"81" => output := x"af4c0775";
            when x"82" => output := x"eebbdd99";
            when x"83" => output := x"a3fd607f";
            when x"84" => output := x"f79f2601";
            when x"85" => output := x"5cbcf572";
            when x"86" => output := x"44c53b66";
            when x"87" => output := x"5b347efb";
            when x"88" => output := x"8b762943";
            when x"89" => output := x"cbdcc623";
            when x"8a" => output := x"b668fced";
            when x"8b" => output := x"b863f1e4";
            when x"8c" => output := x"d7cadc31";
            when x"8d" => output := x"42108563";
            when x"8e" => output := x"13402297";
            when x"8f" => output := x"842011c6";
            when x"90" => output := x"857d244a";
            when x"91" => output := x"d2f83dbb";
            when x"92" => output := x"ae1132f9";
            when x"93" => output := x"c76da129";
            when x"94" => output := x"1d4b2f9e";
            when x"95" => output := x"dcf330b2";
            when x"96" => output := x"0dec5286";
            when x"97" => output := x"77d0e3c1";
            when x"98" => output := x"2b6c16b3";
            when x"99" => output := x"a999b970";
            when x"9a" => output := x"11fa4894";
            when x"9b" => output := x"472264e9";
            when x"9c" => output := x"a8c48cfc";
            when x"9d" => output := x"a01a3ff0";
            when x"9e" => output := x"56d82c7d";
            when x"9f" => output := x"22ef9033";
            when x"a0" => output := x"87c74e49";
            when x"a1" => output := x"d9c1d138";
            when x"a2" => output := x"8cfea2ca";
            when x"a3" => output := x"98360bd4";
            when x"a4" => output := x"a6cf81f5";
            when x"a5" => output := x"a528de7a";
            when x"a6" => output := x"da268eb7";
            when x"a7" => output := x"3fa4bfad";
            when x"a8" => output := x"2ce49d3a";
            when x"a9" => output := x"500d9278";
            when x"aa" => output := x"6a9bcc5f";
            when x"ab" => output := x"5462467e";
            when x"ac" => output := x"f6c2138d";
            when x"ad" => output := x"90e8b8d8";
            when x"ae" => output := x"2e5ef739";
            when x"af" => output := x"82f5afc3";
            when x"b0" => output := x"9fbe805d";
            when x"b1" => output := x"697c93d0";
            when x"b2" => output := x"6fa92dd5";
            when x"b3" => output := x"cfb31225";
            when x"b4" => output := x"c83b99ac";
            when x"b5" => output := x"10a77d18";
            when x"b6" => output := x"e86e639c";
            when x"b7" => output := x"db7bbb3b";
            when x"b8" => output := x"cd097826";
            when x"b9" => output := x"6ef41859";
            when x"ba" => output := x"ec01b79a";
            when x"bb" => output := x"83a89a4f";
            when x"bc" => output := x"e6656e95";
            when x"bd" => output := x"aa7ee6ff";
            when x"be" => output := x"2108cfbc";
            when x"bf" => output := x"efe6e815";
            when x"c0" => output := x"bad99be7";
            when x"c1" => output := x"4ace366f";
            when x"c2" => output := x"ead4099f";
            when x"c3" => output := x"29d67cb0";
            when x"c4" => output := x"31afb2a4";
            when x"c5" => output := x"2a31233f";
            when x"c6" => output := x"c63094a5";
            when x"c7" => output := x"35c066a2";
            when x"c8" => output := x"7437bc4e";
            when x"c9" => output := x"fca6ca82";
            when x"ca" => output := x"e0b0d090";
            when x"cb" => output := x"3315d8a7";
            when x"cc" => output := x"f14a9804";
            when x"cd" => output := x"41f7daec";
            when x"ce" => output := x"7f0e50cd";
            when x"cf" => output := x"172ff691";
            when x"d0" => output := x"768dd64d";
            when x"d1" => output := x"434db0ef";
            when x"d2" => output := x"cc544daa";
            when x"d3" => output := x"e4df0496";
            when x"d4" => output := x"9ee3b5d1";
            when x"d5" => output := x"4c1b886a";
            when x"d6" => output := x"c1b81f2c";
            when x"d7" => output := x"467f5165";
            when x"d8" => output := x"9d04ea5e";
            when x"d9" => output := x"015d358c";
            when x"da" => output := x"fa737487";
            when x"db" => output := x"fb2e410b";
            when x"dc" => output := x"b35a1d67";
            when x"dd" => output := x"9252d2db";
            when x"de" => output := x"e9335610";
            when x"df" => output := x"6d1347d6";
            when x"e0" => output := x"9a8c61d7";
            when x"e1" => output := x"377a0ca1";
            when x"e2" => output := x"598e14f8";
            when x"e3" => output := x"eb893c13";
            when x"e4" => output := x"ceee27a9";
            when x"e5" => output := x"b735c961";
            when x"e6" => output := x"e1ede51c";
            when x"e7" => output := x"7a3cb147";
            when x"e8" => output := x"9c59dfd2";
            when x"e9" => output := x"553f73f2";
            when x"ea" => output := x"1879ce14";
            when x"eb" => output := x"73bf37c7";
            when x"ec" => output := x"53eacdf7";
            when x"ed" => output := x"5f5baafd";
            when x"ee" => output := x"df146f3d";
            when x"ef" => output := x"7886db44";
            when x"f0" => output := x"ca81f3af";
            when x"f1" => output := x"b93ec468";
            when x"f2" => output := x"382c3424";
            when x"f3" => output := x"c25f40a3";
            when x"f4" => output := x"1672c31d";
            when x"f5" => output := x"bc0c25e2";
            when x"f6" => output := x"288b493c";
            when x"f7" => output := x"ff41950d";
            when x"f8" => output := x"397101a8";
            when x"f9" => output := x"08deb30c";
            when x"fa" => output := x"d89ce4b4";
            when x"fb" => output := x"6490c156";
            when x"fc" => output := x"7b6184cb";
            when x"fd" => output := x"d570b632";
            when x"fe" => output := x"48745c6c";
            when x"ff" => output := x"d04257b8";
            when others => null;
        end case;

        return output;
    end;

end aes_sbox;